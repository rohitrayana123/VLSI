magic
tech c035u
timestamp 1394714437
<< error_s >>
rect 27146 30021 27154 30031
rect 27156 30001 27164 30021
rect 27366 30009 27374 30023
rect 27466 30009 27470 30023
rect 27650 30021 27654 30031
rect 27746 30021 27754 30031
rect 27156 29983 27158 30001
rect 27372 29983 27374 30009
rect 27468 29983 27470 30009
rect 27564 29983 27566 30021
rect 27660 30001 27664 30021
rect 27756 30001 27764 30021
rect 27966 30009 27974 30023
rect 28066 30009 28070 30023
rect 28250 30021 28254 30031
rect 28346 30021 28354 30031
rect 27660 29983 27662 30001
rect 27756 29983 27758 30001
rect 27972 29983 27974 30009
rect 28068 29983 28070 30009
rect 28164 29983 28166 30021
rect 28260 30001 28264 30021
rect 28356 30001 28364 30021
rect 28566 30009 28574 30023
rect 28666 30009 28670 30023
rect 28850 30021 28854 30031
rect 28946 30021 28954 30031
rect 28260 29983 28262 30001
rect 28356 29983 28358 30001
rect 28572 29984 28574 30009
rect 28537 29983 28595 29984
rect 28668 29983 28670 30009
rect 28764 29983 28766 30021
rect 28860 30001 28864 30021
rect 28956 30001 28964 30021
rect 29166 30009 29174 30023
rect 29266 30009 29270 30023
rect 29450 30021 29454 30031
rect 29546 30021 29554 30031
rect 28860 29983 28862 30001
rect 28956 29984 28958 30001
rect 28921 29983 28979 29984
rect 29172 29983 29174 30009
rect 29268 29983 29270 30009
rect 29364 29983 29366 30021
rect 29460 30001 29464 30021
rect 29556 30001 29564 30021
rect 29766 30009 29774 30023
rect 29866 30009 29870 30023
rect 30050 30021 30054 30031
rect 30146 30021 30154 30031
rect 29460 29983 29462 30001
rect 29556 29983 29558 30001
rect 29772 29983 29774 30009
rect 29868 29983 29870 30009
rect 29964 29983 29966 30021
rect 30060 30001 30064 30021
rect 30156 30001 30164 30021
rect 30366 30009 30374 30023
rect 30060 29983 30062 30001
rect 30156 29983 30158 30001
rect 30372 29983 30374 30009
rect 30466 30008 30470 30023
rect 30566 30021 30567 30024
rect 30650 30021 30654 30031
rect 30746 30021 30754 30031
rect 30543 30000 30546 30007
rect 30556 30000 30557 30007
rect 30564 30000 30567 30021
rect 30660 30001 30664 30021
rect 30756 30001 30764 30021
rect 30966 30009 30974 30023
rect 31066 30009 31070 30023
rect 31250 30021 31254 30031
rect 31346 30021 31354 30031
rect 30409 29983 30443 29984
rect 30660 29983 30662 30001
rect 30756 29983 30758 30001
rect 30972 29983 30974 30009
rect 31068 29983 31070 30009
rect 31164 29983 31166 30021
rect 31260 30001 31264 30021
rect 31356 30001 31364 30021
rect 31566 30009 31574 30023
rect 31666 30009 31670 30023
rect 31850 30021 31854 30031
rect 31946 30021 31954 30031
rect 31260 29983 31262 30001
rect 31356 29983 31358 30001
rect 31572 29984 31574 30009
rect 31668 29984 31670 30009
rect 31764 29984 31766 30021
rect 31860 30001 31864 30021
rect 31956 30001 31964 30021
rect 32166 30008 32175 30024
rect 31860 29984 31862 30001
rect 31956 29984 31958 30001
rect 32174 30000 32175 30008
rect 31465 29983 31499 29984
rect 27087 29979 30443 29983
rect 30456 29979 30522 29983
rect 30546 29979 31499 29983
rect 31561 29979 31595 29984
rect 31657 29979 31691 29984
rect 31753 29979 31787 29984
rect 31849 29979 31883 29984
rect 31945 29979 31979 29984
rect 27087 29976 27101 29979
rect 27156 29959 27158 29979
rect 27169 29959 27227 29960
rect 27372 29959 27374 29979
rect 27468 29959 27470 29979
rect 27564 29959 27566 29979
rect 27660 29959 27662 29979
rect 27756 29959 27758 29979
rect 27972 29959 27974 29979
rect 28068 29959 28070 29979
rect 28164 29959 28166 29979
rect 28260 29959 28262 29979
rect 28356 29959 28358 29979
rect 28561 29974 28564 29979
rect 28572 29974 28574 29979
rect 28571 29960 28574 29974
rect 28572 29959 28574 29960
rect 28668 29976 28670 29979
rect 28668 29959 28671 29976
rect 28764 29959 28766 29979
rect 28860 29959 28862 29979
rect 28945 29974 28948 29979
rect 28956 29974 28958 29979
rect 28955 29960 28958 29974
rect 29172 29959 29174 29979
rect 29268 29960 29270 29979
rect 29257 29959 29291 29960
rect 29364 29959 29366 29979
rect 29460 29959 29462 29979
rect 29556 29959 29558 29979
rect 29772 29959 29774 29979
rect 29868 29959 29870 29979
rect 29964 29959 29966 29979
rect 30060 29959 30062 29979
rect 30156 29959 30158 29979
rect 30372 29960 30374 29979
rect 30337 29959 30395 29960
rect 30660 29959 30662 29979
rect 30756 29959 30758 29979
rect 30972 29959 30974 29979
rect 31068 29960 31070 29979
rect 31164 29960 31166 29979
rect 31260 29960 31262 29979
rect 31356 29960 31358 29979
rect 31561 29974 31564 29979
rect 31572 29976 31574 29979
rect 31572 29974 31575 29976
rect 31657 29974 31660 29979
rect 31668 29976 31670 29979
rect 31668 29974 31671 29976
rect 31753 29974 31756 29979
rect 31764 29976 31766 29979
rect 31764 29974 31767 29976
rect 31849 29974 31852 29979
rect 31860 29976 31862 29979
rect 31860 29974 31863 29976
rect 31945 29974 31948 29979
rect 31956 29976 31958 29979
rect 31956 29974 31959 29976
rect 31571 29960 31575 29974
rect 31667 29960 31671 29974
rect 31763 29960 31767 29974
rect 31859 29960 31863 29974
rect 31955 29960 31959 29974
rect 31057 29959 31091 29960
rect 27063 29955 28637 29959
rect 27063 29952 27077 29955
rect 27060 29935 27063 29952
rect 27156 29935 27158 29955
rect 27276 29936 27279 29952
rect 27241 29935 27269 29936
rect 27039 29931 27269 29935
rect 27039 29928 27053 29931
rect 27060 29928 27063 29931
rect 27060 29911 27062 29928
rect 27156 29911 27158 29931
rect 27241 29926 27244 29931
rect 27255 29928 27269 29931
rect 27276 29935 27299 29936
rect 27372 29935 27374 29955
rect 27468 29935 27470 29955
rect 27564 29935 27566 29955
rect 27660 29935 27662 29955
rect 27756 29935 27758 29955
rect 27972 29935 27974 29955
rect 28068 29935 28070 29955
rect 28164 29935 28166 29955
rect 28260 29935 28262 29955
rect 28356 29935 28358 29955
rect 28417 29935 28451 29936
rect 27276 29931 28451 29935
rect 28537 29935 28571 29936
rect 28572 29935 28574 29955
rect 28623 29952 28637 29955
rect 28647 29955 29021 29959
rect 28647 29952 28661 29955
rect 28668 29952 28671 29955
rect 28668 29935 28670 29952
rect 28764 29935 28766 29955
rect 28860 29935 28862 29955
rect 29007 29952 29021 29955
rect 29031 29955 30509 29959
rect 30522 29955 31091 29959
rect 31153 29955 31187 29960
rect 31249 29955 31283 29960
rect 31345 29955 31379 29960
rect 29031 29952 29045 29955
rect 29172 29935 29174 29955
rect 29257 29950 29260 29955
rect 29268 29950 29270 29955
rect 29267 29936 29270 29950
rect 29364 29952 29366 29955
rect 29209 29935 29243 29936
rect 29364 29935 29367 29952
rect 29460 29935 29462 29955
rect 29556 29935 29558 29955
rect 29641 29935 29699 29936
rect 29772 29935 29774 29955
rect 29868 29935 29870 29955
rect 29964 29935 29966 29955
rect 30060 29935 30062 29955
rect 30156 29935 30158 29955
rect 30361 29950 30364 29955
rect 30372 29950 30374 29955
rect 30495 29952 30509 29955
rect 30371 29936 30374 29950
rect 30660 29935 30662 29955
rect 30756 29935 30758 29955
rect 30972 29936 30974 29955
rect 31057 29950 31060 29955
rect 31068 29950 31070 29955
rect 31153 29950 31156 29955
rect 31164 29952 31166 29955
rect 31164 29950 31167 29952
rect 31249 29950 31252 29955
rect 31260 29952 31262 29955
rect 31260 29950 31263 29952
rect 31345 29950 31348 29955
rect 31356 29952 31358 29955
rect 31574 29952 31575 29960
rect 31670 29952 31671 29960
rect 31766 29952 31767 29960
rect 31862 29952 31863 29960
rect 31958 29952 31959 29960
rect 32054 29952 32055 29976
rect 31356 29950 31359 29952
rect 31067 29936 31070 29950
rect 31163 29936 31167 29950
rect 31259 29936 31263 29950
rect 31355 29936 31359 29950
rect 28537 29931 29243 29935
rect 29256 29931 29322 29935
rect 29343 29931 30437 29935
rect 27276 29928 27293 29931
rect 27372 29928 27374 29931
rect 27265 29926 27268 29928
rect 27276 29926 27278 29928
rect 27251 29912 27254 29926
rect 27275 29912 27278 29926
rect 27252 29911 27254 29912
rect 27372 29911 27375 29928
rect 27468 29911 27470 29931
rect 27564 29911 27566 29931
rect 27660 29911 27662 29931
rect 27756 29911 27758 29931
rect 27972 29911 27974 29931
rect 28068 29911 28070 29931
rect 28164 29911 28166 29931
rect 28260 29911 28262 29931
rect 28356 29911 28358 29931
rect 27015 29907 27341 29911
rect 27015 29904 27029 29907
rect 27012 29887 27015 29904
rect 27060 29887 27062 29907
rect 27156 29887 27158 29907
rect 27252 29887 27254 29907
rect 27327 29904 27341 29907
rect 27351 29907 28517 29911
rect 27351 29904 27365 29907
rect 27372 29904 27375 29907
rect 27468 29887 27470 29907
rect 27564 29887 27566 29907
rect 27660 29887 27662 29907
rect 27756 29887 27758 29907
rect 27972 29887 27974 29907
rect 28068 29887 28070 29907
rect 28164 29887 28166 29907
rect 28260 29887 28262 29907
rect 28356 29887 28358 29907
rect 28503 29904 28517 29907
rect 28572 29887 28574 29931
rect 28668 29911 28670 29931
rect 28764 29911 28766 29931
rect 28860 29911 28862 29931
rect 29172 29911 29174 29931
rect 29343 29928 29357 29931
rect 29364 29928 29367 29931
rect 29460 29911 29462 29931
rect 29556 29911 29558 29931
rect 29641 29926 29644 29931
rect 29772 29928 29774 29931
rect 29651 29912 29654 29926
rect 29652 29911 29654 29912
rect 29772 29911 29775 29928
rect 29868 29912 29870 29931
rect 29964 29912 29966 29931
rect 30060 29912 30062 29931
rect 30156 29912 30158 29931
rect 30423 29928 30437 29931
rect 30447 29931 30922 29935
rect 30961 29931 30995 29936
rect 30447 29928 30461 29931
rect 29857 29911 29891 29912
rect 28623 29907 29309 29911
rect 29322 29907 29741 29911
rect 28623 29904 28637 29907
rect 28668 29887 28670 29907
rect 28764 29887 28766 29907
rect 28860 29887 28862 29907
rect 29172 29888 29174 29907
rect 29295 29904 29309 29907
rect 28921 29887 28955 29888
rect 29161 29887 29195 29888
rect 26991 29883 29195 29887
rect 29209 29887 29243 29888
rect 29460 29887 29462 29907
rect 29556 29888 29558 29907
rect 29652 29888 29654 29907
rect 29727 29904 29741 29907
rect 29751 29907 29891 29911
rect 29953 29907 29987 29912
rect 30049 29907 30083 29912
rect 30145 29907 30179 29912
rect 30265 29907 30299 29912
rect 30337 29911 30371 29912
rect 30660 29911 30662 29931
rect 30756 29912 30758 29931
rect 30961 29926 30964 29931
rect 30972 29926 30974 29931
rect 31166 29928 31167 29936
rect 31262 29928 31263 29936
rect 31358 29928 31359 29936
rect 30971 29912 30974 29926
rect 30721 29911 30779 29912
rect 30337 29907 30779 29911
rect 30865 29907 30899 29912
rect 29751 29904 29765 29907
rect 29772 29904 29775 29907
rect 29857 29902 29860 29907
rect 29868 29902 29870 29907
rect 29953 29902 29956 29907
rect 29964 29904 29966 29907
rect 29964 29902 29967 29904
rect 30049 29902 30052 29907
rect 30060 29904 30062 29907
rect 30060 29902 30063 29904
rect 30145 29902 30148 29907
rect 30156 29904 30158 29907
rect 30156 29902 30159 29904
rect 29867 29888 29870 29902
rect 29963 29888 29967 29902
rect 30059 29888 30063 29902
rect 30155 29888 30159 29902
rect 30361 29894 30365 29902
rect 30351 29888 30361 29894
rect 30660 29888 30662 29907
rect 30745 29902 30748 29907
rect 30756 29902 30758 29907
rect 31070 29904 31071 29928
rect 30755 29888 30758 29902
rect 29545 29887 29579 29888
rect 29209 29883 29579 29887
rect 29641 29887 29675 29888
rect 29641 29883 29890 29887
rect 26991 29880 27005 29883
rect 27012 29880 27015 29883
rect 26988 29863 26991 29880
rect 27012 29863 27014 29880
rect 27060 29863 27062 29883
rect 27156 29863 27158 29883
rect 27252 29864 27254 29883
rect 27217 29863 27275 29864
rect 27468 29863 27470 29883
rect 27564 29863 27566 29883
rect 27660 29863 27662 29883
rect 27756 29863 27758 29883
rect 27972 29863 27974 29883
rect 28068 29863 28070 29883
rect 28164 29863 28166 29883
rect 28260 29864 28262 29883
rect 28249 29863 28283 29864
rect 26967 29859 28283 29863
rect 26967 29856 26981 29859
rect 26988 29856 26991 29859
rect 26964 29839 26967 29856
rect 26988 29839 26990 29856
rect 27012 29839 27014 29859
rect 27060 29839 27062 29859
rect 27156 29839 27158 29859
rect 27241 29854 27244 29859
rect 27252 29854 27254 29859
rect 27251 29840 27254 29854
rect 27468 29839 27470 29859
rect 27564 29839 27566 29859
rect 27660 29839 27662 29859
rect 27756 29839 27758 29859
rect 27972 29839 27974 29859
rect 28068 29840 28070 29859
rect 28057 29839 28091 29840
rect 26943 29835 27317 29839
rect 26943 29832 26957 29835
rect 26964 29832 26967 29835
rect 26940 29815 26943 29832
rect 26964 29815 26966 29832
rect 26988 29815 26990 29835
rect 27012 29815 27014 29835
rect 27060 29815 27062 29835
rect 27156 29815 27158 29835
rect 27303 29832 27317 29835
rect 27327 29835 28091 29839
rect 27327 29832 27341 29835
rect 27468 29815 27470 29835
rect 27564 29815 27566 29835
rect 27660 29815 27662 29835
rect 27756 29815 27758 29835
rect 27972 29815 27974 29835
rect 28057 29830 28060 29835
rect 28068 29830 28070 29835
rect 28067 29816 28070 29830
rect 28164 29832 28166 29859
rect 28249 29854 28252 29859
rect 28260 29854 28262 29859
rect 28259 29840 28262 29854
rect 28356 29856 28358 29883
rect 28356 29832 28359 29856
rect 26919 29811 28157 29815
rect 26919 29808 26933 29811
rect 26940 29808 26943 29811
rect 26916 29791 26919 29808
rect 26940 29791 26942 29808
rect 26964 29791 26966 29811
rect 26988 29791 26990 29811
rect 27012 29791 27014 29811
rect 27060 29791 27062 29811
rect 27156 29791 27158 29811
rect 27468 29791 27470 29811
rect 27564 29791 27566 29811
rect 27660 29791 27662 29811
rect 27756 29791 27758 29811
rect 27972 29791 27974 29811
rect 28143 29808 28157 29811
rect 28164 29808 28167 29832
rect 28572 29791 28574 29883
rect 28668 29791 28670 29883
rect 28764 29791 28766 29883
rect 28860 29791 28862 29883
rect 29161 29878 29164 29883
rect 29172 29878 29174 29883
rect 29171 29864 29174 29878
rect 29460 29864 29462 29883
rect 29545 29878 29548 29883
rect 29556 29878 29558 29883
rect 29641 29878 29644 29883
rect 29652 29880 29654 29883
rect 29966 29880 29967 29888
rect 30062 29880 30063 29888
rect 30158 29880 30159 29888
rect 30423 29887 30443 29888
rect 30423 29883 30634 29887
rect 30649 29883 30683 29888
rect 30720 29883 30778 29887
rect 30423 29880 30437 29883
rect 29652 29878 29655 29880
rect 30649 29878 30652 29883
rect 30660 29878 30662 29883
rect 30974 29880 30975 29904
rect 29555 29864 29558 29878
rect 29651 29864 29655 29878
rect 30659 29864 30662 29878
rect 29065 29863 29099 29864
rect 28920 29859 28986 29863
rect 29007 29859 29099 29863
rect 29449 29859 29483 29864
rect 29761 29859 29795 29864
rect 30553 29859 30587 29864
rect 29007 29856 29021 29859
rect 29137 29835 29150 29840
rect 29151 29832 29165 29840
rect 29174 29832 29175 29856
rect 29449 29854 29452 29859
rect 29460 29854 29462 29859
rect 30735 29858 30738 29864
rect 30744 29858 30749 29864
rect 30735 29856 30749 29858
rect 30758 29856 30759 29867
rect 29459 29840 29462 29854
rect 29870 29832 29871 29856
rect 30662 29832 30663 29856
rect 29223 29808 29237 29815
rect 29247 29808 29261 29815
rect 29857 29806 29860 29816
rect 29870 29806 29871 29808
rect 29953 29806 29956 29816
rect 29966 29806 29967 29808
rect 30049 29806 30052 29816
rect 30062 29806 30063 29808
rect 30145 29806 30148 29816
rect 30158 29806 30159 29808
rect 29867 29792 29871 29806
rect 29963 29792 29967 29806
rect 30059 29792 30063 29806
rect 30155 29792 30159 29806
rect 26895 29787 29548 29791
rect 26895 29784 26909 29787
rect 26916 29784 26919 29787
rect 26892 29767 26895 29784
rect 26916 29767 26918 29784
rect 26940 29767 26942 29787
rect 26964 29767 26966 29787
rect 26988 29767 26990 29787
rect 27012 29767 27014 29787
rect 27060 29767 27062 29787
rect 27156 29767 27158 29787
rect 27468 29767 27470 29787
rect 27564 29767 27566 29787
rect 27660 29767 27662 29787
rect 27756 29767 27758 29787
rect 27972 29767 27974 29787
rect 28153 29767 28187 29768
rect 26871 29763 28187 29767
rect 26871 29760 26885 29763
rect 26892 29760 26895 29763
rect 26868 29743 26871 29760
rect 26892 29743 26894 29760
rect 26916 29743 26918 29763
rect 26940 29743 26942 29763
rect 26964 29743 26966 29763
rect 26988 29743 26990 29763
rect 27012 29743 27014 29763
rect 27060 29743 27062 29763
rect 27156 29743 27158 29763
rect 27468 29743 27470 29763
rect 27564 29743 27566 29763
rect 27660 29743 27662 29763
rect 27756 29743 27758 29763
rect 27972 29743 27974 29763
rect 26847 29739 28253 29743
rect 26847 29736 26861 29739
rect 26868 29736 26871 29739
rect 26844 29719 26847 29736
rect 26868 29719 26870 29736
rect 26892 29719 26894 29739
rect 26916 29719 26918 29739
rect 26940 29719 26942 29739
rect 26964 29719 26966 29739
rect 26988 29719 26990 29739
rect 27012 29719 27014 29739
rect 27060 29719 27062 29739
rect 27156 29719 27158 29739
rect 27468 29719 27470 29739
rect 27564 29719 27566 29739
rect 27660 29719 27662 29739
rect 27756 29719 27758 29739
rect 27972 29719 27974 29739
rect 28239 29736 28253 29739
rect 28572 29719 28574 29787
rect 28668 29719 28670 29787
rect 28764 29719 28766 29787
rect 28860 29719 28862 29787
rect 29847 29784 29861 29791
rect 29868 29784 29871 29792
rect 29943 29784 29957 29791
rect 29964 29784 29967 29792
rect 30039 29784 30053 29791
rect 30060 29784 30063 29792
rect 30135 29784 30149 29791
rect 30156 29784 30159 29792
rect 30231 29784 30245 29791
rect 30351 29784 30365 29791
rect 29868 29719 29870 29784
rect 29964 29719 29966 29784
rect 30060 29719 30062 29784
rect 30156 29720 30158 29784
rect 30601 29763 30614 29768
rect 30624 29763 30635 29768
rect 30145 29719 30179 29720
rect 26823 29715 30179 29719
rect 26823 29712 26837 29715
rect 26844 29712 26847 29715
rect 26820 29695 26823 29712
rect 26844 29695 26846 29712
rect 26868 29695 26870 29715
rect 26892 29695 26894 29715
rect 26916 29695 26918 29715
rect 26940 29695 26942 29715
rect 26964 29695 26966 29715
rect 26988 29695 26990 29715
rect 27012 29695 27014 29715
rect 27060 29695 27062 29715
rect 27156 29695 27158 29715
rect 27468 29695 27470 29715
rect 27564 29695 27566 29715
rect 27660 29695 27662 29715
rect 27756 29695 27758 29715
rect 27972 29695 27974 29715
rect 28572 29695 28574 29715
rect 28668 29696 28670 29715
rect 28657 29695 28691 29696
rect 26799 29691 28691 29695
rect 26799 29688 26813 29691
rect 26820 29688 26823 29691
rect 26796 29671 26799 29688
rect 26820 29671 26822 29688
rect 26844 29671 26846 29691
rect 26868 29671 26870 29691
rect 26892 29671 26894 29691
rect 26916 29671 26918 29691
rect 26940 29671 26942 29691
rect 26964 29671 26966 29691
rect 26988 29671 26990 29691
rect 27012 29671 27014 29691
rect 27060 29671 27062 29691
rect 27156 29671 27158 29691
rect 27468 29671 27470 29691
rect 27564 29671 27566 29691
rect 27660 29671 27662 29691
rect 27756 29671 27758 29691
rect 27972 29671 27974 29691
rect 28572 29671 28574 29691
rect 28657 29686 28660 29691
rect 28668 29686 28670 29691
rect 28667 29672 28670 29686
rect 28764 29688 28766 29715
rect 26775 29667 28757 29671
rect 26775 29664 26789 29667
rect 26796 29664 26799 29667
rect 26772 29647 26775 29664
rect 26796 29647 26798 29664
rect 26820 29647 26822 29667
rect 26844 29647 26846 29667
rect 26868 29647 26870 29667
rect 26892 29647 26894 29667
rect 26916 29647 26918 29667
rect 26940 29647 26942 29667
rect 26964 29647 26966 29667
rect 26988 29647 26990 29667
rect 27012 29647 27014 29667
rect 27060 29647 27062 29667
rect 27156 29647 27158 29667
rect 27468 29647 27470 29667
rect 27564 29647 27566 29667
rect 27660 29647 27662 29667
rect 27756 29647 27758 29667
rect 27972 29647 27974 29667
rect 28572 29648 28574 29667
rect 28743 29664 28757 29667
rect 28764 29664 28767 29688
rect 28860 29648 28862 29715
rect 29868 29648 29870 29715
rect 29964 29648 29966 29715
rect 30060 29648 30062 29715
rect 30145 29710 30148 29715
rect 30156 29710 30158 29715
rect 30155 29696 30158 29710
rect 30807 29664 30821 29671
rect 30831 29664 30845 29671
rect 28561 29647 28595 29648
rect 26751 29643 28595 29647
rect 28753 29643 28787 29648
rect 28849 29643 28883 29648
rect 29137 29643 29195 29648
rect 29353 29643 29387 29648
rect 29761 29643 29795 29648
rect 29857 29643 29891 29648
rect 29953 29643 29987 29648
rect 30049 29643 30083 29648
rect 30265 29643 30299 29648
rect 30601 29643 30635 29648
rect 30721 29643 30779 29648
rect 26751 29640 26765 29643
rect 26772 29640 26775 29643
rect 26748 29623 26751 29640
rect 26772 29623 26774 29640
rect 26796 29623 26798 29643
rect 26820 29623 26822 29643
rect 26844 29623 26846 29643
rect 26868 29623 26870 29643
rect 26892 29623 26894 29643
rect 26916 29623 26918 29643
rect 26940 29623 26942 29643
rect 26964 29623 26966 29643
rect 26988 29623 26990 29643
rect 27012 29623 27014 29643
rect 27060 29623 27062 29643
rect 27156 29623 27158 29643
rect 27468 29623 27470 29643
rect 27564 29623 27566 29643
rect 27660 29623 27662 29643
rect 27756 29623 27758 29643
rect 27972 29623 27974 29643
rect 28561 29638 28564 29643
rect 28572 29638 28574 29643
rect 28849 29638 28852 29643
rect 28860 29640 28862 29643
rect 28860 29638 28863 29640
rect 29857 29638 29860 29643
rect 29868 29640 29870 29643
rect 29868 29638 29871 29640
rect 29953 29638 29956 29643
rect 29964 29640 29966 29643
rect 29964 29638 29967 29640
rect 30049 29638 30052 29643
rect 30060 29640 30062 29643
rect 30060 29638 30063 29640
rect 28571 29624 28574 29638
rect 28859 29624 28863 29638
rect 29867 29624 29871 29638
rect 29963 29624 29967 29638
rect 30059 29624 30063 29638
rect 26727 29619 28661 29623
rect 26727 29616 26741 29619
rect 26748 29616 26751 29619
rect 26703 29568 26717 29575
rect 26724 29568 26727 29592
rect 26724 29552 26726 29568
rect 26748 29552 26750 29616
rect 26772 29552 26774 29619
rect 26796 29552 26798 29619
rect 26820 29552 26822 29619
rect 26844 29552 26846 29619
rect 26868 29552 26870 29619
rect 26892 29552 26894 29619
rect 26916 29552 26918 29619
rect 26940 29552 26942 29619
rect 26964 29552 26966 29619
rect 26988 29552 26990 29619
rect 27012 29552 27014 29619
rect 27060 29600 27062 29619
rect 27049 29599 27083 29600
rect 27156 29599 27158 29619
rect 27193 29599 27251 29600
rect 27468 29599 27470 29619
rect 27564 29599 27566 29619
rect 27660 29599 27662 29619
rect 27756 29599 27758 29619
rect 27972 29600 27974 29619
rect 28647 29616 28661 29619
rect 28862 29616 28863 29624
rect 29870 29616 29871 29624
rect 29966 29616 29967 29624
rect 30062 29616 30063 29624
rect 27865 29599 27899 29600
rect 27049 29595 27899 29599
rect 27961 29595 27995 29600
rect 28345 29595 28379 29600
rect 28417 29595 28451 29600
rect 28465 29595 28499 29600
rect 27049 29590 27052 29595
rect 27060 29590 27062 29595
rect 27059 29576 27062 29590
rect 27156 29592 27158 29595
rect 27156 29575 27159 29592
rect 27361 29575 27395 29576
rect 27468 29575 27470 29595
rect 27564 29575 27566 29595
rect 27660 29575 27662 29595
rect 27756 29576 27758 29595
rect 27961 29590 27964 29595
rect 27972 29592 27974 29595
rect 27972 29590 27975 29592
rect 27971 29576 27975 29590
rect 28441 29582 28445 29590
rect 28431 29576 28441 29582
rect 27135 29571 27293 29575
rect 27135 29568 27149 29571
rect 27156 29568 27159 29571
rect 27279 29568 27293 29571
rect 27303 29571 27730 29575
rect 27745 29571 27779 29576
rect 27303 29568 27317 29571
rect 27468 29568 27470 29571
rect 26689 29547 27035 29552
rect 27145 29551 27203 29552
rect 27468 29551 27471 29568
rect 27564 29551 27566 29571
rect 27660 29552 27662 29571
rect 27745 29566 27748 29571
rect 27756 29566 27758 29571
rect 27974 29568 27975 29576
rect 27755 29552 27758 29566
rect 27649 29551 27683 29552
rect 27145 29547 27346 29551
rect 27360 29547 27426 29551
rect 27447 29547 27683 29551
rect 26689 29542 26692 29547
rect 26713 29542 26716 29547
rect 26724 29544 26726 29547
rect 26724 29542 26727 29544
rect 26699 29528 26702 29542
rect 26713 29534 26717 29542
rect 26723 29534 26727 29542
rect 26737 29542 26740 29547
rect 26748 29544 26750 29547
rect 26748 29542 26751 29544
rect 26737 29534 26741 29542
rect 26747 29534 26751 29542
rect 26761 29542 26764 29547
rect 26772 29544 26774 29547
rect 26772 29542 26775 29544
rect 26761 29534 26765 29542
rect 26771 29534 26775 29542
rect 26785 29542 26788 29547
rect 26796 29544 26798 29547
rect 26796 29542 26799 29544
rect 26785 29534 26789 29542
rect 26795 29534 26799 29542
rect 26809 29542 26812 29547
rect 26820 29544 26822 29547
rect 26820 29542 26823 29544
rect 26809 29534 26813 29542
rect 26819 29534 26823 29542
rect 26833 29542 26836 29547
rect 26844 29544 26846 29547
rect 26844 29542 26847 29544
rect 26833 29534 26837 29542
rect 26843 29534 26847 29542
rect 26857 29542 26860 29547
rect 26868 29544 26870 29547
rect 26868 29542 26871 29544
rect 26857 29534 26861 29542
rect 26867 29534 26871 29542
rect 26881 29542 26884 29547
rect 26892 29544 26894 29547
rect 26892 29542 26895 29544
rect 26881 29534 26885 29542
rect 26891 29534 26895 29542
rect 26905 29542 26908 29547
rect 26916 29544 26918 29547
rect 26916 29542 26919 29544
rect 26905 29534 26909 29542
rect 26915 29534 26919 29542
rect 26929 29542 26932 29547
rect 26940 29544 26942 29547
rect 26940 29542 26943 29544
rect 26929 29534 26933 29542
rect 26939 29534 26943 29542
rect 26953 29542 26956 29547
rect 26964 29544 26966 29547
rect 26964 29542 26967 29544
rect 26953 29534 26957 29542
rect 26963 29534 26967 29542
rect 26977 29542 26980 29547
rect 26988 29544 26990 29547
rect 26988 29542 26991 29544
rect 26977 29534 26981 29542
rect 26987 29534 26991 29542
rect 27001 29542 27004 29547
rect 27012 29544 27014 29547
rect 27447 29544 27461 29547
rect 27468 29544 27471 29547
rect 27012 29542 27015 29544
rect 27001 29534 27005 29542
rect 27011 29534 27015 29542
rect 27025 29534 27029 29542
rect 26703 29528 26713 29534
rect 26723 29528 26737 29534
rect 26747 29528 26761 29534
rect 26771 29528 26785 29534
rect 26795 29528 26809 29534
rect 26819 29528 26833 29534
rect 26843 29528 26857 29534
rect 26867 29528 26881 29534
rect 26891 29528 26905 29534
rect 26915 29528 26929 29534
rect 26939 29528 26953 29534
rect 26963 29528 26977 29534
rect 26987 29528 27001 29534
rect 27011 29528 27025 29534
rect 27564 29528 27566 29547
rect 27649 29542 27652 29547
rect 27660 29542 27662 29547
rect 27659 29528 27662 29542
rect 26726 29520 26727 29528
rect 26750 29520 26751 29528
rect 26774 29520 26775 29528
rect 26798 29520 26799 29528
rect 26822 29520 26823 29528
rect 26846 29520 26847 29528
rect 26870 29520 26871 29528
rect 26894 29520 26895 29528
rect 26918 29520 26919 29528
rect 26942 29520 26943 29528
rect 26966 29520 26967 29528
rect 26990 29520 26991 29528
rect 27014 29520 27015 29528
rect 27457 29527 27491 29528
rect 27336 29523 27402 29527
rect 27426 29523 27491 29527
rect 27553 29523 27587 29528
rect 27553 29518 27556 29523
rect 27564 29520 27566 29523
rect 27758 29520 27759 29544
rect 27564 29518 27567 29520
rect 27563 29504 27567 29518
rect 27566 29496 27567 29504
rect 25599 28323 26630 28327
rect 25599 28320 25613 28323
rect 24999 28299 26654 28303
rect 24999 28296 25013 28299
rect 24879 28275 26678 28279
rect 24879 28272 24893 28275
rect 24615 28251 26702 28255
rect 24615 28248 24629 28251
rect 24540 28231 24543 28248
rect 24519 28227 26726 28231
rect 24519 28224 24533 28227
rect 24540 28224 24543 28227
rect 23473 28207 23507 28208
rect 24540 28207 24542 28224
rect 24793 28207 24851 28208
rect 23343 28203 23507 28207
rect 24399 28203 26750 28207
rect 23343 28200 23357 28203
rect 24399 28200 24413 28203
rect 23268 28183 23271 28200
rect 24540 28183 24542 28203
rect 24924 28183 24927 28200
rect 22215 28179 23021 28183
rect 22215 28176 22229 28179
rect 23007 28176 23021 28179
rect 23247 28179 23573 28183
rect 23247 28176 23261 28179
rect 23268 28176 23271 28179
rect 23559 28176 23573 28179
rect 24255 28179 24893 28183
rect 24255 28176 24269 28179
rect 23268 28159 23270 28176
rect 24540 28160 24542 28179
rect 24879 28176 24893 28179
rect 24903 28179 26774 28183
rect 24903 28176 24917 28179
rect 24924 28176 24927 28179
rect 24529 28159 24587 28160
rect 24924 28159 24926 28176
rect 22071 28155 26798 28159
rect 22071 28152 22085 28155
rect 23268 28135 23270 28155
rect 24015 28152 24029 28155
rect 24529 28150 24532 28155
rect 24540 28150 24542 28155
rect 24539 28136 24542 28150
rect 24924 28135 24926 28155
rect 25129 28135 25163 28136
rect 21951 28131 24629 28135
rect 21951 28128 21965 28131
rect 23268 28111 23270 28131
rect 24615 28128 24629 28131
rect 24639 28131 26822 28135
rect 24639 28128 24653 28131
rect 24924 28111 24926 28131
rect 21831 28107 26846 28111
rect 21831 28104 21845 28107
rect 21635 28088 21639 28102
rect 21471 28083 21629 28087
rect 21471 28080 21485 28083
rect 21615 28080 21629 28083
rect 21636 28080 21639 28088
rect 23161 28087 23219 28088
rect 23268 28087 23270 28107
rect 24924 28087 24926 28107
rect 25215 28104 25229 28107
rect 21711 28083 26870 28087
rect 21711 28080 21725 28083
rect 23268 28080 23270 28083
rect 21636 28064 21638 28080
rect 21625 28063 21683 28064
rect 23268 28063 23271 28080
rect 24924 28063 24926 28083
rect 21327 28059 23261 28063
rect 21327 28056 21341 28059
rect 21625 28054 21628 28059
rect 21636 28054 21638 28059
rect 23247 28056 23261 28059
rect 23268 28059 26894 28063
rect 23268 28056 23285 28059
rect 21635 28040 21638 28054
rect 5329 28039 5363 28040
rect 21756 28039 21759 28056
rect 23257 28039 23315 28040
rect 24924 28039 24926 28059
rect 4863 28035 5363 28039
rect 21255 28035 21725 28039
rect 4863 28032 4877 28035
rect 21255 28032 21269 28035
rect 21711 28032 21725 28035
rect 21735 28035 26918 28039
rect 21735 28032 21749 28035
rect 21756 28032 21759 28035
rect 21756 28015 21758 28032
rect 23281 28030 23284 28035
rect 23291 28016 23294 28030
rect 23292 28015 23294 28016
rect 24924 28015 24926 28035
rect 4839 28011 5429 28015
rect 4839 28008 4853 28011
rect 5415 28008 5429 28011
rect 6927 28011 11741 28015
rect 6927 28008 6941 28011
rect 11727 28008 11741 28011
rect 21207 28011 23357 28015
rect 21207 28008 21221 28011
rect 4753 27991 4787 27992
rect 4551 27987 4787 27991
rect 4801 27991 4835 27992
rect 21241 27991 21299 27992
rect 21756 27991 21758 28011
rect 23292 27991 23294 28011
rect 23343 28008 23357 28011
rect 23367 28011 26942 28015
rect 23367 28008 23381 28011
rect 24924 27991 24926 28011
rect 4801 27987 12005 27991
rect 4551 27984 4565 27987
rect 11991 27984 12005 27987
rect 20751 27987 26966 27991
rect 20751 27984 20765 27987
rect 21265 27982 21268 27987
rect 21275 27968 21278 27982
rect 21276 27967 21278 27968
rect 21756 27967 21758 27987
rect 23292 27967 23294 27987
rect 24924 27967 24926 27987
rect 4444 27963 4853 27967
rect 4839 27960 4853 27963
rect 4887 27963 13181 27967
rect 4887 27960 4901 27963
rect 13167 27960 13181 27963
rect 13599 27963 15437 27967
rect 13599 27960 13613 27963
rect 15423 27960 15437 27963
rect 20631 27963 21341 27967
rect 20631 27960 20645 27963
rect 4476 27943 4479 27960
rect 21276 27943 21278 27963
rect 21327 27960 21341 27963
rect 21351 27963 26990 27967
rect 27001 27963 27014 27968
rect 27024 27963 27035 27968
rect 21351 27960 21365 27963
rect 21756 27943 21758 27963
rect 23292 27943 23294 27963
rect 24924 27943 24926 27963
rect 27492 27943 27495 27960
rect 29857 27958 29860 27968
rect 29870 27958 29871 27960
rect 29953 27958 29956 27968
rect 29966 27958 29967 27960
rect 30049 27958 30052 27968
rect 30062 27958 30063 27960
rect 28441 27950 28445 27958
rect 28431 27944 28441 27950
rect 29867 27944 29871 27958
rect 29963 27944 29967 27958
rect 30059 27944 30063 27958
rect 4335 27939 4444 27943
rect 4455 27939 16013 27943
rect 4335 27936 4349 27939
rect 4455 27936 4469 27939
rect 4476 27936 4479 27939
rect 15999 27936 16013 27939
rect 20295 27939 27076 27943
rect 20295 27936 20309 27939
rect 4476 27919 4478 27936
rect 19643 27920 19647 27934
rect 19644 27919 19647 27920
rect 21276 27919 21278 27939
rect 21756 27919 21758 27939
rect 23292 27919 23294 27939
rect 24924 27919 24926 27939
rect 27087 27936 27101 27943
rect 27231 27936 27245 27943
rect 27471 27939 27652 27943
rect 27471 27936 27485 27939
rect 27492 27936 27495 27939
rect 27783 27936 27797 27943
rect 27807 27939 27844 27943
rect 27807 27936 27821 27939
rect 28047 27936 28061 27943
rect 28431 27936 28445 27943
rect 28503 27936 28517 27943
rect 28551 27936 28565 27943
rect 28935 27936 28949 27943
rect 29223 27936 29237 27943
rect 29247 27936 29261 27943
rect 29439 27936 29453 27943
rect 29847 27936 29861 27943
rect 29868 27936 29871 27944
rect 29943 27936 29957 27943
rect 29964 27936 29967 27944
rect 30039 27936 30053 27943
rect 30060 27936 30063 27944
rect 30135 27936 30149 27943
rect 30351 27936 30365 27943
rect 30687 27936 30701 27943
rect 30807 27936 30821 27943
rect 30831 27936 30845 27943
rect 27001 27919 27035 27920
rect 3964 27915 16733 27919
rect 4476 27895 4478 27915
rect 16719 27912 16733 27915
rect 17319 27915 18269 27919
rect 17319 27912 17333 27915
rect 18255 27912 18269 27915
rect 18399 27915 18869 27919
rect 18399 27912 18413 27915
rect 18855 27912 18869 27915
rect 19623 27915 19685 27919
rect 19623 27912 19637 27915
rect 19644 27912 19647 27915
rect 19671 27912 19685 27915
rect 19719 27915 27035 27919
rect 27337 27919 27371 27920
rect 27492 27919 27494 27936
rect 29868 27920 29870 27936
rect 29964 27920 29966 27936
rect 30060 27920 30062 27936
rect 27745 27919 27779 27920
rect 27337 27915 27779 27919
rect 27961 27915 27995 27920
rect 28345 27915 28379 27920
rect 29161 27915 29195 27920
rect 29353 27915 29387 27920
rect 29761 27915 29795 27920
rect 29857 27915 29891 27920
rect 29953 27915 29987 27920
rect 30049 27915 30083 27920
rect 30265 27915 30299 27920
rect 30601 27915 30635 27920
rect 30721 27915 30779 27920
rect 30889 27915 30923 27920
rect 19719 27912 19733 27915
rect 19644 27895 19646 27912
rect 21121 27895 21179 27896
rect 21276 27895 21278 27915
rect 21756 27896 21758 27915
rect 21745 27895 21803 27896
rect 23292 27895 23294 27915
rect 24924 27895 24926 27915
rect 27423 27895 27443 27896
rect 27492 27895 27494 27915
rect 29857 27910 29860 27915
rect 29868 27912 29870 27915
rect 29868 27910 29871 27912
rect 29953 27910 29956 27915
rect 29964 27912 29966 27915
rect 29964 27910 29967 27912
rect 30049 27910 30052 27915
rect 30060 27912 30062 27915
rect 30060 27910 30063 27912
rect 29867 27896 29871 27910
rect 29963 27896 29967 27910
rect 30059 27896 30063 27910
rect 364 27891 3964 27895
rect 3975 27891 19037 27895
rect 3975 27888 3989 27891
rect 4476 27871 4478 27891
rect 19023 27888 19037 27891
rect 19479 27891 27101 27895
rect 19479 27888 19493 27891
rect 19644 27871 19646 27891
rect 21276 27871 21278 27891
rect 21745 27886 21748 27891
rect 21756 27886 21758 27891
rect 21755 27872 21758 27886
rect 21876 27871 21879 27888
rect 22129 27871 22187 27872
rect 23292 27871 23294 27891
rect 24924 27871 24926 27891
rect 27087 27888 27101 27891
rect 27423 27891 27845 27895
rect 27423 27888 27437 27891
rect 27492 27888 27494 27891
rect 27831 27888 27845 27891
rect 29870 27888 29871 27896
rect 29966 27888 29967 27896
rect 30062 27888 30063 27896
rect 27492 27871 27495 27888
rect 27516 27871 27519 27888
rect -1137 27867 364 27871
rect 375 27867 21221 27871
rect -1137 27864 -1123 27867
rect 375 27864 389 27867
rect -1175 27847 -1141 27848
rect 4476 27847 4478 27867
rect 18097 27847 18131 27848
rect 19393 27847 19451 27848
rect 19644 27847 19646 27867
rect 21207 27864 21221 27867
rect 21231 27867 21845 27871
rect 21231 27864 21245 27867
rect 21276 27847 21278 27867
rect 21831 27864 21845 27867
rect 21855 27867 27485 27871
rect 21855 27864 21869 27867
rect 21876 27864 21879 27867
rect 21876 27847 21878 27864
rect 23292 27847 23294 27867
rect 24924 27847 24926 27867
rect 27471 27864 27485 27867
rect 27492 27867 28060 27871
rect 28263 27867 28444 27871
rect 27492 27864 27509 27867
rect 27516 27864 27519 27867
rect 28263 27864 28277 27867
rect 27516 27847 27518 27864
rect 28177 27847 28211 27848
rect 28465 27847 28499 27848
rect -1209 27843 22229 27847
rect -1209 27840 -1195 27843
rect 4476 27823 4478 27843
rect 17233 27823 17291 27824
rect 19644 27823 19646 27843
rect 20665 27823 20723 27824
rect 21276 27823 21278 27843
rect 21876 27823 21878 27843
rect 22215 27840 22229 27843
rect 22239 27843 28499 27847
rect 28849 27843 28883 27848
rect 28969 27847 29003 27848
rect 28969 27843 29260 27847
rect 22239 27840 22253 27843
rect 23292 27823 23294 27843
rect 24924 27823 24926 27843
rect 27516 27823 27518 27843
rect 29857 27838 29860 27848
rect 29867 27824 29870 27838
rect 28225 27823 28259 27824
rect -1713 27819 19493 27823
rect -1713 27816 -1699 27819
rect -1089 27816 -1075 27819
rect 4476 27799 4478 27819
rect 18183 27816 18197 27819
rect 19479 27816 19493 27819
rect 19503 27819 28214 27823
rect 28225 27819 28277 27823
rect 28300 27819 28565 27823
rect 19503 27816 19517 27819
rect 19644 27799 19646 27819
rect 21276 27799 21278 27819
rect 21876 27800 21878 27819
rect 21865 27799 21923 27800
rect 23292 27799 23294 27819
rect 24924 27799 24926 27819
rect 27516 27799 27518 27819
rect 28263 27816 28277 27819
rect 28551 27816 28565 27819
rect 28935 27816 28949 27824
rect 29055 27819 29452 27823
rect 29751 27819 29860 27823
rect 29055 27816 29069 27819
rect 29751 27816 29765 27819
rect 29943 27816 29957 27823
rect 29966 27816 29967 27840
rect 29665 27799 29723 27800
rect -2145 27795 17333 27799
rect -2145 27792 -2131 27795
rect -1295 27775 -1237 27776
rect 4476 27775 4478 27795
rect 17319 27792 17333 27795
rect 17343 27795 20765 27799
rect 17343 27792 17357 27795
rect 19644 27775 19646 27795
rect 20751 27792 20765 27795
rect 20775 27795 28300 27799
rect 28311 27795 28948 27799
rect 29007 27795 30052 27799
rect 20775 27792 20789 27795
rect 21276 27775 21278 27795
rect 21865 27790 21868 27795
rect 21876 27790 21878 27795
rect 21875 27776 21878 27790
rect 21996 27775 21999 27792
rect 23292 27775 23294 27795
rect 24924 27775 24926 27795
rect 27516 27775 27518 27795
rect 28311 27792 28325 27795
rect 29007 27792 29021 27795
rect 31153 27790 31156 27800
rect 31166 27790 31167 27792
rect 31249 27790 31252 27800
rect 31262 27790 31263 27792
rect 31345 27790 31348 27800
rect 31358 27790 31359 27792
rect 31657 27790 31660 27800
rect 31670 27790 31671 27792
rect 31753 27790 31756 27800
rect 31766 27790 31767 27792
rect 31849 27790 31852 27800
rect 31862 27790 31863 27792
rect 31163 27776 31167 27790
rect 31259 27776 31263 27790
rect 31355 27776 31359 27790
rect 31667 27776 31671 27790
rect 31763 27776 31767 27790
rect 31859 27776 31863 27790
rect -2457 27771 21965 27775
rect -2457 27768 -2443 27771
rect -3383 27751 -3349 27752
rect -1164 27751 -1161 27768
rect 1801 27751 1835 27752
rect 1897 27751 1931 27752
rect 2377 27751 2411 27752
rect 3409 27751 3443 27752
rect 4476 27751 4478 27771
rect 6457 27751 6491 27752
rect 12913 27751 12947 27752
rect 13585 27751 13619 27752
rect 13777 27751 13811 27752
rect 19644 27751 19646 27771
rect 20473 27751 20507 27752
rect 21276 27751 21278 27771
rect 21951 27768 21965 27771
rect 21975 27771 29765 27775
rect 21975 27768 21989 27771
rect 21996 27768 21999 27771
rect 21996 27751 21998 27768
rect 23292 27751 23294 27771
rect 24924 27751 24926 27771
rect 27516 27751 27518 27771
rect 29751 27768 29765 27771
rect 29775 27771 30148 27775
rect 29775 27768 29789 27771
rect 30351 27768 30365 27775
rect 30687 27768 30701 27775
rect 30807 27768 30821 27775
rect 30831 27768 30845 27775
rect 30975 27768 30989 27775
rect 31119 27768 31133 27775
rect 31143 27768 31157 27775
rect 31164 27768 31167 27776
rect 31239 27768 31253 27775
rect 31260 27768 31263 27776
rect 31335 27768 31349 27775
rect 31356 27768 31359 27776
rect 31431 27768 31445 27775
rect 31647 27768 31661 27775
rect 31668 27768 31671 27776
rect 31743 27768 31757 27775
rect 31764 27768 31767 27776
rect 31839 27768 31853 27775
rect 31860 27768 31863 27776
rect 31935 27768 31949 27775
rect 31958 27768 31959 27792
rect 31164 27751 31166 27768
rect 31260 27751 31262 27768
rect 31356 27751 31358 27768
rect 31668 27751 31670 27768
rect 31764 27751 31766 27768
rect 31860 27752 31862 27768
rect 31849 27751 31883 27752
rect -5073 27747 -1195 27751
rect -5073 27744 -5059 27747
rect -1209 27744 -1195 27747
rect -1185 27747 31883 27751
rect -1185 27744 -1171 27747
rect -1164 27744 -1161 27747
rect -5148 27727 -5145 27744
rect -1164 27727 -1162 27744
rect 1907 27728 1911 27742
rect 1908 27727 1911 27728
rect 4476 27727 4478 27747
rect 18313 27727 18371 27728
rect 19644 27727 19646 27747
rect 21276 27727 21278 27747
rect 21996 27727 21998 27747
rect 23292 27727 23294 27747
rect 24121 27727 24155 27728
rect 24924 27727 24926 27747
rect 27516 27727 27518 27747
rect 30265 27727 30299 27728
rect -5169 27723 30299 27727
rect 30721 27723 30755 27728
rect -5169 27720 -5155 27723
rect -5148 27720 -5145 27723
rect -3297 27720 -3283 27723
rect -5148 27703 -5146 27720
rect -1164 27703 -1162 27723
rect 1887 27720 1901 27723
rect 1908 27720 1911 27723
rect 1983 27720 1997 27723
rect 2463 27720 2477 27723
rect 3495 27720 3509 27723
rect 1908 27703 1910 27720
rect 4476 27703 4478 27723
rect 6543 27720 6557 27723
rect 12999 27720 13013 27723
rect 13671 27720 13685 27723
rect 13863 27720 13877 27723
rect 19644 27703 19646 27723
rect 20559 27720 20573 27723
rect 20209 27703 20267 27704
rect 21276 27703 21278 27723
rect 21996 27704 21998 27723
rect 21985 27703 22043 27704
rect 23292 27703 23294 27723
rect 24313 27703 24371 27704
rect 24924 27703 24926 27723
rect 27409 27703 27467 27704
rect 27516 27703 27518 27723
rect 28921 27703 28979 27704
rect 29665 27703 29699 27704
rect -5732 27699 18413 27703
rect -5808 27685 -5804 27693
rect -5148 27679 -5146 27699
rect -1164 27679 -1162 27699
rect 1908 27679 1910 27699
rect 4476 27679 4478 27699
rect 18399 27696 18413 27699
rect 18423 27699 30365 27703
rect 18423 27696 18437 27699
rect 19644 27679 19646 27699
rect 21276 27679 21278 27699
rect 21985 27694 21988 27699
rect 21996 27694 21998 27699
rect 21995 27680 21998 27694
rect 23292 27679 23294 27699
rect 24207 27696 24221 27699
rect 24444 27679 24447 27696
rect 24924 27679 24926 27699
rect 27433 27694 27436 27699
rect 27516 27696 27518 27699
rect 30351 27696 30365 27699
rect 27443 27680 27446 27694
rect 27444 27679 27446 27680
rect 27516 27679 27519 27696
rect -5804 27675 -5732 27679
rect -5721 27675 20309 27679
rect -5721 27672 -5707 27675
rect -5148 27656 -5146 27675
rect -5159 27655 -5101 27656
rect -1164 27655 -1162 27675
rect 1908 27655 1910 27675
rect 4476 27655 4478 27675
rect 19537 27655 19595 27656
rect 19644 27655 19646 27675
rect 20295 27672 20309 27675
rect 20319 27675 22085 27679
rect 20319 27672 20333 27675
rect 21276 27655 21278 27675
rect 22071 27672 22085 27675
rect 22095 27675 24413 27679
rect 22095 27672 22109 27675
rect 23292 27655 23294 27675
rect 24399 27672 24413 27675
rect 24423 27675 27509 27679
rect 24423 27672 24437 27675
rect 24444 27672 24447 27675
rect 24444 27656 24446 27672
rect 24433 27655 24491 27656
rect 24924 27655 24926 27675
rect 27444 27656 27446 27675
rect 27495 27672 27509 27675
rect 27516 27675 29021 27679
rect 27516 27672 27533 27675
rect 29007 27672 29021 27675
rect 29031 27675 30485 27679
rect 29031 27672 29045 27675
rect 29751 27672 29765 27675
rect 30471 27672 30485 27675
rect 30495 27675 30820 27679
rect 30495 27672 30509 27675
rect 27433 27655 27491 27656
rect 30409 27655 30467 27656
rect 31057 27655 31091 27656
rect -6945 27651 -5804 27655
rect -5793 27651 31091 27655
rect -6945 27648 -6931 27651
rect -5793 27648 -5779 27651
rect -7020 27632 -7017 27648
rect -5159 27646 -5156 27651
rect -5148 27646 -5146 27651
rect -5149 27632 -5146 27646
rect -7031 27631 -6973 27632
rect -1164 27631 -1162 27651
rect 1908 27631 1910 27651
rect 4476 27631 4478 27651
rect 19644 27648 19646 27651
rect 19644 27631 19647 27648
rect 20545 27631 20603 27632
rect 21276 27631 21278 27651
rect 23292 27631 23294 27651
rect 24433 27646 24436 27651
rect 24444 27646 24446 27651
rect 24443 27632 24446 27646
rect 24564 27631 24567 27648
rect 24924 27631 24926 27651
rect 27433 27646 27436 27651
rect 27444 27646 27446 27651
rect 27443 27632 27446 27646
rect 31164 27648 31166 27747
rect -7041 27627 -5059 27631
rect -7041 27624 -7027 27627
rect -7020 27624 -7017 27627
rect -5073 27624 -5059 27627
rect -5049 27627 19637 27631
rect -5049 27624 -5035 27627
rect -7031 27622 -7028 27624
rect -7020 27622 -7018 27624
rect -7021 27608 -7018 27622
rect -2543 27607 -2485 27608
rect -1164 27607 -1162 27627
rect 1908 27607 1910 27627
rect 4249 27607 4307 27608
rect 4476 27607 4478 27627
rect 19623 27624 19637 27627
rect 19644 27627 24533 27631
rect 19644 27624 19661 27627
rect 20569 27622 20572 27627
rect 20579 27608 20582 27622
rect 20580 27607 20582 27608
rect 21276 27607 21278 27627
rect 21385 27607 21443 27608
rect 23292 27607 23294 27627
rect 24519 27624 24533 27627
rect 24543 27627 27533 27631
rect 24543 27624 24557 27627
rect 24564 27624 24567 27627
rect 24564 27607 24566 27624
rect 24924 27608 24926 27627
rect 27519 27624 27533 27627
rect 27543 27627 30509 27631
rect 27543 27624 27557 27627
rect 30495 27624 30509 27627
rect 30519 27627 31157 27631
rect 30519 27624 30533 27627
rect 31143 27624 31157 27627
rect 31164 27624 31167 27648
rect 24913 27607 24971 27608
rect 27457 27607 27491 27608
rect -10857 27603 -6931 27607
rect -10857 27600 -10843 27603
rect -6945 27600 -6931 27603
rect -6921 27603 20645 27607
rect -6921 27600 -6907 27603
rect -8975 27583 -8941 27584
rect -1799 27583 -1741 27584
rect -1164 27583 -1162 27603
rect -167 27583 -133 27584
rect 1908 27583 1910 27603
rect 4380 27583 4383 27600
rect 4476 27583 4478 27603
rect 20580 27583 20582 27603
rect 20631 27600 20645 27603
rect 20655 27603 27491 27607
rect 27505 27607 27539 27608
rect 28225 27607 28283 27608
rect 29689 27607 29747 27608
rect 31153 27607 31187 27608
rect 27505 27603 31187 27607
rect 20655 27600 20669 27603
rect 21169 27583 21227 27584
rect 21276 27583 21278 27603
rect 23292 27583 23294 27603
rect 24564 27583 24566 27603
rect 24913 27598 24916 27603
rect 24924 27598 24926 27603
rect 24923 27584 24926 27598
rect 31260 27600 31262 27747
rect -15465 27579 -2443 27583
rect -15465 27576 -15451 27579
rect -2457 27576 -2443 27579
rect -2433 27579 4349 27583
rect -2433 27576 -2419 27579
rect -17653 27560 -17649 27574
rect -17652 27559 -17649 27560
rect -14591 27559 -14557 27560
rect -2231 27559 -2173 27560
rect -1223 27559 -1165 27560
rect -1164 27559 -1162 27579
rect 1908 27559 1910 27579
rect 4335 27576 4349 27579
rect 4359 27579 21485 27583
rect 4359 27576 4373 27579
rect 4380 27576 4383 27579
rect 4380 27559 4382 27576
rect 4476 27559 4478 27579
rect 4777 27559 4811 27560
rect -18369 27555 -1699 27559
rect -18369 27552 -18355 27555
rect -17673 27552 -17659 27555
rect -17652 27552 -17649 27555
rect -17577 27552 -17563 27555
rect -8889 27552 -8875 27555
rect -1713 27552 -1699 27555
rect -1689 27555 4811 27559
rect 4825 27559 4859 27560
rect 20580 27559 20582 27579
rect 21276 27576 21278 27579
rect 21471 27576 21485 27579
rect 21495 27579 25013 27583
rect 21495 27576 21509 27579
rect 21276 27559 21279 27576
rect 23292 27559 23294 27579
rect 24564 27559 24566 27579
rect 24999 27576 25013 27579
rect 25023 27579 27557 27583
rect 25023 27576 25037 27579
rect 27543 27576 27557 27579
rect 27591 27579 28325 27583
rect 27591 27576 27605 27579
rect 28311 27576 28325 27579
rect 28335 27579 29789 27583
rect 28335 27576 28349 27579
rect 29775 27576 29789 27579
rect 29799 27579 31253 27583
rect 29799 27576 29813 27579
rect 31239 27576 31253 27579
rect 31260 27576 31263 27600
rect 31356 27559 31358 27747
rect 31668 27728 31670 27747
rect 31764 27728 31766 27747
rect 31849 27742 31852 27747
rect 31860 27742 31862 27747
rect 31859 27728 31862 27742
rect 31561 27723 31595 27728
rect 31657 27723 31691 27728
rect 31753 27723 31787 27728
rect 31657 27718 31660 27723
rect 31668 27720 31670 27723
rect 31668 27718 31671 27720
rect 31753 27718 31756 27723
rect 31764 27720 31766 27723
rect 31764 27718 31767 27720
rect 31667 27704 31671 27718
rect 31763 27704 31767 27718
rect 31670 27696 31671 27704
rect 31766 27696 31767 27704
rect 31753 27603 31756 27608
rect 31839 27576 31853 27583
rect 4825 27555 21269 27559
rect -1689 27552 -1675 27555
rect -17652 27535 -17650 27552
rect -15551 27535 -15493 27536
rect -7127 27535 -7069 27536
rect -6407 27535 -6373 27536
rect -1164 27535 -1162 27555
rect -81 27552 -67 27555
rect 1908 27535 1910 27555
rect 4380 27535 4382 27555
rect 4476 27535 4478 27555
rect 19633 27535 19691 27536
rect 20580 27535 20582 27555
rect 21255 27552 21269 27555
rect 21276 27555 32164 27559
rect 21276 27552 21293 27555
rect 23292 27535 23294 27555
rect 24564 27535 24566 27555
rect 27481 27535 27539 27536
rect 28969 27535 29027 27536
rect 31249 27535 31283 27536
rect -18513 27531 -2131 27535
rect -18513 27528 -18499 27531
rect -18588 27512 -18585 27528
rect -18599 27511 -18541 27512
rect -17652 27511 -17650 27531
rect -14505 27528 -14491 27531
rect -2145 27528 -2131 27531
rect -2121 27531 -1123 27535
rect -2121 27528 -2107 27531
rect -16991 27511 -16957 27512
rect -15503 27511 -15469 27512
rect -14951 27511 -14917 27512
rect -6996 27511 -6993 27528
rect -5255 27511 -5197 27512
rect -1164 27511 -1162 27531
rect -1137 27528 -1123 27531
rect -1113 27531 4877 27535
rect -1113 27528 -1099 27531
rect 1908 27511 1910 27531
rect 4380 27511 4382 27531
rect 4476 27511 4478 27531
rect 4863 27528 4877 27531
rect 4911 27531 31283 27535
rect 4911 27528 4925 27531
rect 19657 27526 19660 27531
rect 19667 27512 19670 27526
rect 6841 27511 6899 27512
rect 13513 27511 13571 27512
rect 19668 27511 19670 27512
rect 20580 27511 20582 27531
rect 23292 27511 23294 27531
rect 24564 27511 24566 27531
rect 31356 27528 31358 27555
rect 31753 27531 31787 27536
rect 32041 27531 32075 27536
rect -18609 27507 -15451 27511
rect -18609 27504 -18595 27507
rect -18588 27504 -18585 27507
rect -18599 27502 -18596 27504
rect -18588 27502 -18586 27504
rect -18589 27488 -18586 27502
rect -17652 27487 -17650 27507
rect -15465 27504 -15451 27507
rect -15441 27507 -7027 27511
rect -15441 27504 -15427 27507
rect -7041 27504 -7027 27507
rect -7017 27507 19733 27511
rect -7017 27504 -7003 27507
rect -6996 27504 -6993 27507
rect -6321 27504 -6307 27507
rect -6996 27487 -6994 27504
rect -5124 27487 -5121 27504
rect -1164 27487 -1162 27507
rect 1908 27487 1910 27507
rect 4380 27487 4382 27507
rect 4476 27487 4478 27507
rect 19668 27487 19670 27507
rect 19719 27504 19733 27507
rect 19743 27507 27581 27511
rect 19743 27504 19757 27507
rect 20580 27487 20582 27507
rect 23292 27487 23294 27507
rect 24564 27487 24566 27507
rect 27567 27504 27581 27507
rect 27591 27507 29069 27511
rect 27591 27504 27605 27507
rect 29055 27504 29069 27507
rect 29079 27507 31349 27511
rect 29079 27504 29093 27507
rect 31335 27504 31349 27507
rect 31356 27504 31359 27528
rect 27145 27487 27179 27488
rect -18897 27483 -18499 27487
rect -18897 27480 -18883 27483
rect -18513 27480 -18499 27483
rect -18489 27483 -5155 27487
rect -18489 27480 -18475 27483
rect -17652 27463 -17650 27483
rect -16905 27480 -16891 27483
rect -15417 27480 -15403 27483
rect -14865 27480 -14851 27483
rect -6996 27463 -6994 27483
rect -5169 27480 -5155 27483
rect -5145 27483 6941 27487
rect -5145 27480 -5131 27483
rect -5124 27480 -5121 27483
rect -5124 27463 -5122 27480
rect -1164 27463 -1162 27483
rect 1908 27463 1910 27483
rect 4380 27463 4382 27483
rect 4476 27463 4478 27483
rect 6927 27480 6941 27483
rect 6951 27483 13613 27487
rect 6951 27480 6965 27483
rect 13599 27480 13613 27483
rect 13623 27483 27179 27487
rect 27265 27487 27299 27488
rect 27337 27487 27395 27488
rect 31249 27487 31283 27488
rect 27265 27483 31283 27487
rect 31345 27483 31379 27488
rect 13623 27480 13637 27483
rect 19668 27463 19670 27483
rect 20580 27463 20582 27483
rect 23292 27463 23294 27483
rect 24169 27463 24203 27464
rect 24564 27463 24566 27483
rect 31356 27478 31359 27480
rect 27361 27470 27365 27478
rect 27351 27464 27361 27470
rect 27371 27464 27375 27478
rect 31355 27464 31359 27478
rect 25513 27463 25547 27464
rect 27372 27463 27375 27464
rect 27721 27463 27779 27464
rect 28249 27463 28283 27464
rect -18980 27459 27245 27463
rect -17916 27368 -17914 27388
rect -17868 27368 -17866 27388
rect -17820 27368 -17818 27388
rect -17772 27368 -17770 27388
rect -17652 27368 -17650 27459
rect -17532 27368 -17530 27388
rect -17436 27368 -17434 27388
rect -17412 27368 -17410 27388
rect -17364 27368 -17362 27388
rect -17316 27368 -17314 27388
rect -17220 27368 -17218 27388
rect -17196 27368 -17194 27388
rect -17124 27368 -17122 27388
rect -17028 27368 -17026 27388
rect -16980 27368 -16978 27390
rect -16894 27388 -16892 27398
rect -15430 27388 -15428 27398
rect -15406 27388 -15404 27398
rect -16884 27368 -16882 27388
rect -16860 27368 -16858 27388
rect -16812 27368 -16810 27388
rect -16788 27368 -16786 27388
rect -16764 27368 -16762 27388
rect -16716 27368 -16714 27388
rect -16692 27368 -16690 27388
rect -16668 27368 -16666 27388
rect -16596 27368 -16594 27388
rect -16500 27368 -16498 27388
rect -16404 27368 -16402 27388
rect -16380 27368 -16378 27388
rect -16332 27368 -16330 27388
rect -16308 27368 -16306 27388
rect -16284 27368 -16282 27388
rect -16236 27368 -16234 27388
rect -16212 27368 -16210 27388
rect -16188 27368 -16186 27388
rect -15591 27368 -15557 27370
rect -15420 27368 -15418 27388
rect -15396 27368 -15394 27388
rect -15372 27368 -15370 27388
rect -15300 27368 -15298 27388
rect -15084 27368 -15082 27388
rect -15036 27368 -15034 27388
rect -14940 27368 -14938 27390
rect -14494 27388 -14492 27398
rect -14916 27368 -14914 27388
rect -14868 27368 -14866 27388
rect -14820 27368 -14818 27388
rect -14724 27368 -14722 27388
rect -14700 27368 -14698 27388
rect -14652 27368 -14650 27388
rect -14604 27368 -14602 27388
rect -14508 27368 -14506 27388
rect -14484 27368 -14482 27388
rect -14436 27368 -14434 27388
rect -14388 27368 -14386 27388
rect -14268 27368 -14266 27388
rect -14172 27368 -14170 27388
rect -14076 27368 -14074 27388
rect -14028 27368 -14026 27388
rect -13980 27368 -13978 27388
rect -13956 27368 -13954 27388
rect -13932 27368 -13930 27388
rect -13860 27368 -13858 27388
rect -13764 27368 -13762 27388
rect -13716 27368 -13714 27388
rect -13644 27368 -13642 27388
rect -13596 27368 -13594 27388
rect -13500 27368 -13498 27388
rect -13404 27368 -13402 27388
rect -13356 27368 -13354 27388
rect -13284 27368 -13282 27388
rect -12828 27368 -12826 27388
rect -12780 27368 -12778 27388
rect -12684 27368 -12682 27388
rect -12660 27368 -12658 27388
rect -12612 27368 -12610 27388
rect -12588 27368 -12586 27388
rect -12564 27368 -12562 27388
rect -12492 27368 -12490 27388
rect -12396 27368 -12394 27388
rect -12348 27368 -12346 27388
rect -12276 27368 -12274 27388
rect -12252 27368 -12250 27388
rect -12228 27368 -12226 27388
rect -12156 27368 -12154 27388
rect -12060 27368 -12058 27388
rect -12012 27368 -12010 27388
rect -11916 27368 -11914 27388
rect -11892 27368 -11890 27388
rect -11844 27368 -11842 27388
rect -11796 27368 -11794 27388
rect -11676 27368 -11674 27388
rect -11580 27368 -11578 27388
rect -11556 27368 -11554 27388
rect -11484 27368 -11482 27388
rect -11460 27368 -11458 27388
rect -11436 27368 -11434 27388
rect -11388 27368 -11386 27388
rect -11364 27368 -11362 27388
rect -11340 27368 -11338 27388
rect -11268 27368 -11266 27388
rect -11172 27368 -11170 27388
rect -11124 27368 -11122 27388
rect -11076 27368 -11074 27388
rect -11028 27368 -11026 27388
rect -10932 27368 -10930 27390
rect -10846 27388 -10844 27398
rect -10836 27368 -10834 27388
rect -10788 27368 -10786 27388
rect -10668 27368 -10666 27388
rect -10047 27368 -10013 27370
rect -9876 27368 -9874 27388
rect -9828 27368 -9826 27388
rect -9732 27368 -9730 27388
rect -9708 27368 -9706 27388
rect -9612 27368 -9610 27388
rect -9516 27368 -9514 27388
rect -9468 27368 -9466 27388
rect -9420 27368 -9418 27388
rect -9396 27368 -9394 27388
rect -9372 27368 -9370 27388
rect -9300 27368 -9298 27388
rect -9252 27368 -9250 27388
rect -9156 27368 -9154 27388
rect -9132 27368 -9130 27388
rect -9084 27368 -9082 27388
rect -9060 27368 -9058 27388
rect -9036 27368 -9034 27388
rect -8988 27368 -8986 27388
rect -8964 27368 -8962 27390
rect -8940 27368 -8938 27388
rect -8892 27368 -8890 27388
rect -8844 27368 -8842 27388
rect -8796 27368 -8794 27388
rect -8700 27368 -8698 27388
rect -8604 27368 -8602 27388
rect -8556 27368 -8554 27388
rect -8508 27368 -8506 27388
rect -8484 27368 -8482 27388
rect -8460 27368 -8458 27388
rect -8412 27368 -8410 27388
rect -8388 27368 -8386 27388
rect -8364 27368 -8362 27388
rect -8316 27368 -8314 27388
rect -8292 27368 -8290 27388
rect -8268 27368 -8266 27388
rect -8196 27368 -8194 27388
rect -8100 27368 -8098 27388
rect -8052 27368 -8050 27388
rect -7932 27368 -7930 27388
rect -7836 27368 -7834 27388
rect -7740 27368 -7738 27388
rect -7692 27368 -7690 27388
rect -7620 27368 -7618 27388
rect -7356 27368 -7354 27388
rect -7284 27368 -7282 27388
rect -7212 27368 -7210 27388
rect -7188 27368 -7186 27388
rect -7116 27368 -7114 27388
rect -7092 27368 -7090 27390
rect -7068 27368 -7066 27388
rect -6996 27368 -6994 27459
rect -6910 27388 -6908 27398
rect -6972 27368 -6970 27388
rect -6948 27368 -6946 27388
rect -6900 27368 -6898 27388
rect -6876 27368 -6874 27388
rect -6852 27368 -6850 27388
rect -6804 27368 -6802 27388
rect -6780 27368 -6778 27388
rect -6756 27368 -6754 27388
rect -6708 27368 -6706 27388
rect -6684 27368 -6682 27388
rect -6660 27368 -6658 27388
rect -6612 27368 -6610 27388
rect -6588 27368 -6586 27388
rect -6564 27368 -6562 27388
rect -6516 27368 -6514 27388
rect -6492 27368 -6490 27388
rect -6468 27368 -6466 27388
rect -6420 27368 -6418 27388
rect -6396 27368 -6394 27390
rect -6310 27388 -6308 27398
rect -6372 27368 -6370 27388
rect -6324 27368 -6322 27388
rect -6300 27368 -6298 27388
rect -6276 27368 -6274 27388
rect -6228 27368 -6226 27388
rect -6180 27368 -6178 27388
rect -6060 27368 -6058 27388
rect -5964 27368 -5962 27388
rect -5940 27368 -5938 27388
rect -5868 27368 -5866 27390
rect -5796 27368 -5794 27390
rect -5652 27368 -5650 27388
rect -5316 27368 -5314 27388
rect -5268 27368 -5266 27388
rect -5220 27368 -5218 27390
rect -5196 27368 -5194 27388
rect -5172 27368 -5170 27388
rect -5124 27368 -5122 27459
rect -5038 27388 -5036 27398
rect -5100 27368 -5098 27388
rect -5076 27368 -5074 27388
rect -5028 27368 -5026 27388
rect -4980 27368 -4978 27388
rect -4884 27368 -4882 27388
rect -4860 27368 -4858 27388
rect -4788 27368 -4786 27388
rect -4692 27368 -4690 27388
rect -4644 27368 -4642 27388
rect -4596 27368 -4594 27388
rect -4548 27368 -4546 27388
rect -4428 27368 -4426 27388
rect -4332 27368 -4330 27388
rect -4308 27368 -4306 27388
rect -4260 27368 -4258 27388
rect -4212 27368 -4210 27388
rect -4116 27368 -4114 27388
rect -4092 27368 -4090 27388
rect -4020 27368 -4018 27388
rect -3876 27368 -3874 27388
rect -3804 27368 -3802 27388
rect -3732 27368 -3730 27388
rect -3588 27368 -3586 27388
rect -3564 27368 -3562 27388
rect -3516 27368 -3514 27388
rect -3492 27368 -3490 27388
rect -3468 27368 -3466 27388
rect -3420 27368 -3418 27388
rect -3372 27368 -3370 27390
rect -3252 27368 -3250 27388
rect -3156 27368 -3154 27388
rect -3132 27368 -3130 27388
rect -3060 27368 -3058 27388
rect -3012 27368 -3010 27388
rect -2916 27368 -2914 27388
rect -2892 27368 -2890 27388
rect -2844 27368 -2842 27388
rect -2820 27368 -2818 27388
rect -2796 27368 -2794 27388
rect -2748 27368 -2746 27388
rect -2700 27368 -2698 27388
rect -2604 27368 -2602 27388
rect -2580 27368 -2578 27388
rect -2508 27368 -2506 27390
rect -2422 27388 -2420 27398
rect -2412 27368 -2410 27388
rect -2364 27368 -2362 27388
rect -2292 27368 -2290 27388
rect -2268 27368 -2266 27388
rect -2244 27368 -2242 27388
rect -2196 27368 -2194 27390
rect -2110 27388 -2108 27398
rect -2172 27368 -2170 27388
rect -2148 27368 -2146 27388
rect -2100 27368 -2098 27388
rect -2076 27368 -2074 27388
rect -2052 27368 -2050 27388
rect -1980 27368 -1978 27388
rect -1884 27368 -1882 27388
rect -1836 27368 -1834 27388
rect -1716 27368 -1714 27388
rect -1596 27368 -1594 27388
rect -1476 27368 -1474 27388
rect -1380 27368 -1378 27388
rect -1356 27368 -1354 27388
rect -1308 27368 -1306 27388
rect -1260 27368 -1258 27390
rect -1164 27368 -1162 27459
rect -1078 27388 -1076 27398
rect -70 27388 -68 27398
rect -1140 27368 -1138 27388
rect -1068 27368 -1066 27388
rect -852 27368 -850 27388
rect -804 27368 -802 27388
rect -756 27368 -754 27388
rect -708 27368 -706 27388
rect -612 27368 -610 27388
rect -588 27368 -586 27388
rect -540 27368 -538 27388
rect -516 27368 -514 27388
rect -492 27368 -490 27388
rect -444 27368 -442 27388
rect -396 27368 -394 27388
rect -300 27368 -298 27388
rect -276 27368 -274 27388
rect -204 27368 -202 27388
rect -108 27368 -106 27388
rect -60 27368 -58 27388
rect 12 27368 14 27388
rect 108 27368 110 27388
rect 156 27368 158 27388
rect 204 27368 206 27388
rect 228 27368 230 27388
rect 252 27368 254 27388
rect 300 27368 302 27390
rect 348 27368 350 27388
rect 468 27368 470 27388
rect 564 27368 566 27388
rect 588 27368 590 27388
rect 636 27368 638 27388
rect 660 27368 662 27388
rect 684 27368 686 27388
rect 732 27368 734 27388
rect 756 27368 758 27388
rect 780 27368 782 27388
rect 876 27368 878 27388
rect 972 27368 974 27388
rect 1020 27368 1022 27388
rect 1068 27368 1070 27388
rect 1092 27368 1094 27388
rect 1116 27368 1118 27388
rect 1164 27368 1166 27388
rect 1212 27368 1214 27388
rect 1308 27368 1310 27388
rect 1332 27368 1334 27388
rect 1380 27368 1382 27388
rect 1428 27368 1430 27388
rect 1524 27368 1526 27388
rect 1548 27368 1550 27388
rect 1596 27368 1598 27388
rect 1620 27368 1622 27388
rect 1644 27368 1646 27388
rect 1692 27368 1694 27388
rect 1716 27368 1718 27388
rect 1740 27368 1742 27388
rect 1788 27368 1790 27388
rect 1812 27368 1814 27390
rect 1836 27368 1838 27388
rect 1884 27368 1886 27388
rect 1908 27368 1910 27459
rect 1994 27388 1996 27398
rect 1932 27368 1934 27388
rect 1980 27368 1982 27388
rect 2004 27368 2006 27388
rect 2028 27368 2030 27388
rect 2076 27368 2078 27388
rect 2100 27368 2102 27388
rect 2124 27368 2126 27388
rect 2172 27368 2174 27388
rect 2196 27368 2198 27388
rect 2220 27368 2222 27388
rect 2268 27368 2270 27388
rect 2292 27368 2294 27388
rect 2316 27368 2318 27388
rect 2364 27368 2366 27388
rect 2388 27368 2390 27390
rect 2474 27388 2476 27398
rect 3506 27388 3508 27398
rect 2412 27368 2414 27388
rect 2460 27368 2462 27388
rect 2484 27368 2486 27388
rect 2508 27368 2510 27388
rect 2556 27368 2558 27388
rect 2580 27368 2582 27388
rect 2604 27368 2606 27388
rect 2652 27368 2654 27388
rect 2676 27368 2678 27388
rect 2700 27368 2702 27388
rect 2748 27368 2750 27388
rect 2772 27368 2774 27388
rect 2796 27368 2798 27388
rect 2844 27368 2846 27388
rect 2868 27368 2870 27388
rect 2892 27368 2894 27388
rect 2940 27368 2942 27388
rect 3012 27368 3014 27388
rect 3108 27368 3110 27388
rect 3156 27368 3158 27388
rect 3252 27368 3254 27388
rect 3348 27368 3350 27388
rect 3396 27368 3398 27388
rect 3468 27368 3470 27388
rect 3492 27368 3494 27388
rect 3516 27368 3518 27388
rect 3588 27368 3590 27388
rect 3612 27368 3614 27388
rect 3636 27368 3638 27388
rect 3708 27368 3710 27388
rect 3732 27368 3734 27388
rect 3756 27368 3758 27388
rect 3804 27368 3806 27388
rect 3828 27368 3830 27388
rect 3852 27368 3854 27388
rect 3900 27368 3902 27390
rect 3986 27388 3988 27398
rect 3924 27368 3926 27388
rect 3948 27368 3950 27388
rect 3996 27368 3998 27388
rect 4020 27368 4022 27388
rect 4044 27368 4046 27388
rect 4092 27368 4094 27388
rect 4116 27368 4118 27388
rect 4140 27368 4142 27388
rect 4188 27368 4190 27388
rect 4212 27368 4214 27388
rect 4236 27368 4238 27388
rect 4284 27368 4286 27390
rect 4308 27368 4310 27388
rect 4332 27368 4334 27388
rect 4380 27368 4382 27459
rect 4404 27368 4406 27388
rect 4428 27368 4430 27388
rect 4476 27368 4478 27459
rect 4500 27368 4502 27388
rect 4524 27368 4526 27388
rect 4596 27368 4598 27388
rect 4812 27368 4814 27390
rect 4898 27388 4900 27398
rect 4860 27368 4862 27388
rect 4908 27368 4910 27388
rect 4956 27368 4958 27388
rect 4980 27368 4982 27388
rect 5004 27368 5006 27388
rect 5076 27368 5078 27388
rect 5100 27368 5102 27388
rect 5124 27368 5126 27388
rect 5172 27368 5174 27388
rect 5196 27368 5198 27388
rect 5220 27368 5222 27388
rect 5268 27368 5270 27388
rect 5292 27368 5294 27388
rect 5316 27368 5318 27390
rect 5402 27388 5404 27398
rect 5426 27388 5428 27398
rect 5388 27368 5390 27388
rect 5412 27368 5414 27388
rect 5436 27368 5438 27388
rect 5484 27368 5486 27388
rect 5508 27368 5510 27388
rect 5532 27368 5534 27388
rect 5580 27368 5582 27388
rect 5628 27368 5630 27388
rect 5724 27368 5726 27388
rect 5748 27368 5750 27388
rect 5796 27368 5798 27388
rect 5820 27368 5822 27388
rect 5844 27368 5846 27388
rect 5916 27368 5918 27388
rect 6132 27368 6134 27388
rect 6180 27368 6182 27388
rect 6228 27368 6230 27388
rect 6252 27368 6254 27388
rect 6276 27368 6278 27388
rect 6324 27368 6326 27388
rect 6372 27368 6374 27388
rect 6468 27368 6470 27390
rect 6554 27388 6556 27398
rect 6492 27368 6494 27388
rect 6564 27368 6566 27388
rect 6588 27368 6590 27388
rect 6612 27368 6614 27388
rect 6660 27368 6662 27388
rect 6684 27368 6686 27388
rect 6708 27368 6710 27388
rect 6780 27368 6782 27388
rect 6804 27368 6806 27388
rect 6828 27368 6830 27388
rect 6876 27368 6878 27390
rect 6962 27388 6964 27398
rect 6900 27368 6902 27388
rect 6924 27368 6926 27388
rect 6972 27368 6974 27388
rect 7020 27368 7022 27388
rect 7140 27368 7142 27388
rect 7236 27368 7238 27388
rect 7260 27368 7262 27388
rect 7332 27368 7334 27388
rect 7356 27368 7358 27388
rect 7380 27368 7382 27388
rect 7428 27368 7430 27388
rect 7452 27368 7454 27388
rect 7476 27368 7478 27388
rect 7524 27368 7526 27388
rect 7548 27368 7550 27388
rect 7572 27368 7574 27388
rect 7620 27368 7622 27388
rect 7644 27368 7646 27388
rect 7668 27368 7670 27388
rect 7716 27368 7718 27388
rect 7740 27368 7742 27388
rect 7764 27368 7766 27388
rect 7836 27368 7838 27388
rect 7860 27368 7862 27388
rect 7884 27368 7886 27388
rect 7932 27368 7934 27388
rect 7956 27368 7958 27388
rect 7980 27368 7982 27388
rect 8052 27368 8054 27388
rect 8148 27368 8150 27388
rect 8196 27368 8198 27388
rect 8244 27368 8246 27388
rect 8268 27368 8270 27388
rect 8292 27368 8294 27388
rect 8340 27368 8342 27388
rect 8364 27368 8366 27388
rect 8388 27368 8390 27388
rect 8436 27368 8438 27388
rect 8460 27368 8462 27388
rect 8484 27368 8486 27388
rect 8556 27368 8558 27388
rect 8580 27368 8582 27388
rect 8604 27368 8606 27388
rect 8676 27368 8678 27388
rect 8700 27368 8702 27388
rect 8724 27368 8726 27388
rect 8772 27368 8774 27388
rect 8820 27368 8822 27388
rect 8844 27368 8846 27388
rect 8868 27368 8870 27388
rect 9465 27368 9499 27370
rect 9660 27368 9662 27388
rect 9684 27368 9686 27388
rect 9708 27368 9710 27388
rect 9756 27368 9758 27388
rect 9780 27368 9782 27388
rect 9804 27368 9806 27388
rect 9852 27368 9854 27388
rect 9876 27368 9878 27388
rect 9900 27368 9902 27388
rect 9948 27368 9950 27388
rect 9972 27368 9974 27388
rect 9996 27368 9998 27388
rect 10068 27368 10070 27388
rect 10092 27368 10094 27388
rect 10116 27368 10118 27388
rect 10164 27368 10166 27388
rect 10188 27368 10190 27388
rect 10212 27368 10214 27388
rect 10260 27368 10262 27388
rect 10284 27368 10286 27388
rect 10308 27368 10310 27388
rect 10380 27368 10382 27388
rect 10404 27368 10406 27388
rect 10428 27368 10430 27388
rect 10476 27368 10478 27388
rect 10500 27368 10502 27388
rect 10524 27368 10526 27388
rect 10572 27368 10574 27388
rect 10596 27368 10598 27388
rect 10620 27368 10622 27388
rect 10668 27368 10670 27388
rect 10692 27368 10694 27388
rect 10716 27368 10718 27388
rect 10788 27368 10790 27388
rect 10836 27368 10838 27388
rect 10956 27368 10958 27388
rect 11052 27368 11054 27388
rect 11076 27368 11078 27388
rect 11124 27368 11126 27388
rect 11172 27368 11174 27388
rect 11220 27368 11222 27388
rect 11340 27368 11342 27388
rect 11436 27368 11438 27388
rect 11532 27368 11534 27388
rect 11580 27368 11582 27388
rect 11628 27368 11630 27388
rect 11652 27368 11654 27390
rect 11738 27388 11740 27398
rect 12002 27388 12004 27398
rect 11676 27368 11678 27388
rect 11748 27368 11750 27388
rect 11772 27368 11774 27388
rect 11796 27368 11798 27388
rect 11844 27368 11846 27388
rect 11892 27368 11894 27388
rect 11988 27368 11990 27388
rect 12012 27368 12014 27388
rect 12084 27368 12086 27388
rect 12132 27368 12134 27388
rect 12228 27368 12230 27388
rect 12252 27368 12254 27388
rect 12300 27368 12302 27388
rect 12324 27368 12326 27388
rect 12348 27368 12350 27388
rect 12396 27368 12398 27388
rect 12420 27368 12422 27388
rect 12444 27368 12446 27388
rect 12492 27368 12494 27388
rect 12516 27368 12518 27388
rect 12540 27368 12542 27388
rect 12588 27368 12590 27388
rect 12636 27368 12638 27388
rect 12732 27368 12734 27388
rect 12756 27368 12758 27388
rect 12804 27368 12806 27388
rect 12828 27368 12830 27388
rect 12852 27368 12854 27388
rect 12900 27368 12902 27388
rect 12924 27368 12926 27390
rect 13010 27388 13012 27398
rect 13178 27388 13180 27398
rect 13634 27388 13636 27398
rect 13682 27388 13684 27398
rect 12948 27368 12950 27388
rect 13020 27368 13022 27388
rect 13044 27368 13046 27388
rect 13068 27368 13070 27388
rect 13116 27368 13118 27388
rect 13188 27368 13190 27388
rect 13284 27368 13286 27388
rect 13332 27368 13334 27388
rect 13428 27368 13430 27388
rect 13524 27368 13526 27388
rect 13572 27368 13574 27388
rect 13644 27368 13646 27388
rect 13668 27368 13670 27388
rect 13692 27368 13694 27388
rect 13764 27368 13766 27388
rect 13788 27368 13790 27390
rect 13874 27388 13876 27398
rect 13812 27368 13814 27388
rect 13860 27368 13862 27388
rect 13884 27368 13886 27388
rect 13908 27368 13910 27388
rect 13956 27368 13958 27388
rect 14004 27368 14006 27388
rect 14100 27368 14102 27388
rect 14196 27368 14198 27388
rect 14244 27368 14246 27388
rect 14292 27368 14294 27388
rect 14889 27368 14923 27370
rect 15132 27368 15134 27388
rect 15228 27368 15230 27388
rect 15252 27368 15254 27388
rect 15300 27368 15302 27388
rect 15324 27368 15326 27388
rect 15348 27368 15350 27390
rect 15434 27388 15436 27398
rect 15396 27368 15398 27388
rect 15420 27368 15422 27388
rect 15444 27368 15446 27388
rect 15492 27368 15494 27388
rect 15540 27368 15542 27388
rect 15636 27368 15638 27388
rect 15660 27368 15662 27388
rect 15708 27368 15710 27388
rect 15732 27368 15734 27388
rect 15756 27368 15758 27388
rect 15804 27368 15806 27388
rect 15828 27368 15830 27388
rect 15852 27368 15854 27388
rect 15900 27368 15902 27388
rect 15924 27368 15926 27390
rect 16010 27388 16012 27398
rect 15948 27368 15950 27388
rect 15996 27368 15998 27388
rect 16020 27368 16022 27388
rect 16044 27368 16046 27388
rect 16092 27368 16094 27388
rect 16140 27368 16142 27388
rect 16236 27368 16238 27388
rect 16260 27368 16262 27388
rect 16308 27368 16310 27388
rect 16332 27368 16334 27388
rect 16356 27368 16358 27388
rect 16404 27368 16406 27388
rect 16452 27368 16454 27388
rect 16548 27368 16550 27388
rect 16572 27368 16574 27388
rect 16620 27368 16622 27388
rect 16644 27368 16646 27390
rect 16730 27388 16732 27398
rect 16668 27368 16670 27388
rect 16716 27368 16718 27388
rect 16740 27368 16742 27388
rect 16764 27368 16766 27388
rect 16836 27368 16838 27388
rect 16884 27368 16886 27388
rect 16980 27368 16982 27388
rect 17004 27368 17006 27388
rect 17052 27368 17054 27388
rect 17100 27368 17102 27388
rect 17196 27368 17198 27388
rect 17220 27368 17222 27388
rect 17268 27368 17270 27390
rect 17292 27368 17294 27388
rect 17316 27368 17318 27388
rect 17913 27368 17947 27370
rect 18084 27368 18086 27388
rect 18108 27368 18110 27390
rect 18132 27368 18134 27388
rect 18180 27368 18182 27390
rect 18252 27368 18254 27388
rect 18348 27368 18350 27390
rect 18396 27368 18398 27388
rect 18492 27368 18494 27388
rect 18516 27368 18518 27388
rect 18564 27368 18566 27388
rect 18588 27368 18590 27388
rect 18612 27368 18614 27388
rect 18660 27368 18662 27388
rect 18684 27368 18686 27388
rect 18708 27368 18710 27388
rect 18756 27368 18758 27388
rect 18780 27368 18782 27390
rect 18866 27388 18868 27398
rect 18804 27368 18806 27388
rect 18852 27368 18854 27388
rect 18876 27368 18878 27388
rect 18900 27368 18902 27388
rect 18948 27368 18950 27390
rect 19034 27388 19036 27398
rect 18996 27368 18998 27388
rect 19020 27368 19022 27388
rect 19044 27368 19046 27388
rect 19092 27368 19094 27388
rect 19116 27368 19118 27388
rect 19140 27368 19142 27388
rect 19188 27368 19190 27388
rect 19236 27368 19238 27388
rect 19332 27368 19334 27388
rect 19428 27368 19430 27390
rect 19514 27388 19516 27398
rect 19476 27368 19478 27388
rect 19524 27368 19526 27388
rect 19572 27368 19574 27390
rect 19596 27368 19598 27390
rect 19620 27368 19622 27388
rect 19668 27368 19670 27459
rect 19682 27388 19684 27398
rect 19754 27388 19756 27398
rect 19692 27368 19694 27388
rect 19716 27368 19718 27388
rect 19764 27368 19766 27388
rect 19812 27368 19814 27388
rect 19836 27368 19838 27388
rect 19860 27368 19862 27388
rect 19932 27368 19934 27388
rect 19956 27368 19958 27388
rect 19980 27368 19982 27388
rect 20028 27368 20030 27388
rect 20052 27368 20054 27388
rect 20076 27368 20078 27388
rect 20148 27368 20150 27388
rect 20172 27368 20174 27388
rect 20196 27368 20198 27388
rect 20244 27368 20246 27390
rect 20330 27388 20332 27398
rect 20268 27368 20270 27388
rect 20292 27368 20294 27388
rect 20340 27368 20342 27388
rect 20388 27368 20390 27388
rect 20484 27368 20486 27390
rect 20508 27368 20510 27388
rect 20556 27368 20558 27388
rect 20580 27368 20582 27459
rect 20604 27368 20606 27388
rect 20700 27368 20702 27390
rect 20916 27368 20918 27388
rect 20964 27368 20966 27388
rect 21012 27368 21014 27388
rect 21060 27368 21062 27388
rect 21084 27368 21086 27388
rect 21108 27368 21110 27388
rect 21156 27368 21158 27390
rect 21204 27368 21206 27390
rect 21290 27388 21292 27398
rect 21362 27388 21364 27398
rect 21300 27368 21302 27388
rect 21324 27368 21326 27388
rect 21372 27368 21374 27388
rect 21420 27368 21422 27390
rect 21506 27388 21508 27398
rect 21444 27368 21446 27388
rect 21468 27368 21470 27388
rect 21516 27368 21518 27388
rect 21540 27368 21542 27390
rect 21564 27368 21566 27388
rect 21612 27368 21614 27388
rect 21660 27368 21662 27390
rect 21684 27368 21686 27388
rect 21708 27368 21710 27388
rect 21780 27368 21782 27390
rect 21804 27368 21806 27388
rect 21828 27368 21830 27388
rect 21900 27368 21902 27390
rect 21924 27368 21926 27388
rect 21948 27368 21950 27388
rect 22020 27368 22022 27390
rect 22106 27388 22108 27398
rect 22044 27368 22046 27388
rect 22068 27368 22070 27388
rect 22116 27368 22118 27388
rect 22164 27368 22166 27390
rect 22188 27368 22190 27388
rect 22212 27368 22214 27388
rect 22833 27368 22867 27370
rect 23004 27368 23006 27388
rect 23052 27368 23054 27388
rect 23076 27368 23078 27388
rect 23100 27368 23102 27388
rect 23148 27368 23150 27388
rect 23196 27368 23198 27390
rect 23220 27368 23222 27388
rect 23244 27368 23246 27388
rect 23292 27368 23294 27459
rect 24193 27435 24206 27440
rect 24216 27435 24227 27440
rect 23378 27388 23380 27398
rect 23316 27368 23318 27388
rect 23340 27368 23342 27388
rect 23388 27368 23390 27388
rect 23412 27368 23414 27388
rect 23436 27368 23438 27390
rect 23484 27368 23486 27390
rect 23522 27388 23524 27398
rect 23570 27388 23572 27398
rect 24026 27388 24028 27398
rect 23532 27368 23534 27388
rect 23556 27368 23558 27388
rect 23580 27368 23582 27388
rect 23628 27368 23630 27388
rect 23652 27368 23654 27388
rect 23676 27368 23678 27388
rect 23724 27368 23726 27388
rect 23748 27368 23750 27388
rect 23772 27368 23774 27388
rect 23820 27368 23822 27388
rect 23868 27368 23870 27388
rect 23892 27368 23894 27388
rect 23916 27368 23918 27388
rect 23988 27368 23990 27388
rect 24012 27368 24014 27388
rect 24036 27368 24038 27388
rect 24084 27368 24086 27388
rect 24132 27368 24134 27390
rect 24218 27388 24220 27398
rect 24290 27388 24292 27398
rect 24228 27368 24230 27388
rect 24252 27368 24254 27388
rect 24300 27368 24302 27388
rect 24348 27368 24350 27390
rect 24372 27368 24374 27388
rect 24396 27368 24398 27388
rect 24468 27368 24470 27390
rect 24492 27368 24494 27388
rect 24516 27368 24518 27388
rect 24564 27368 24566 27459
rect 27231 27456 27245 27459
rect 27351 27459 27437 27463
rect 27351 27456 27365 27459
rect 27372 27456 27375 27459
rect 27423 27456 27437 27459
rect 27447 27459 31349 27463
rect 27447 27456 27461 27459
rect 31335 27456 31349 27459
rect 31358 27456 31359 27464
rect 25537 27435 25550 27440
rect 25560 27435 25571 27440
rect 24650 27388 24652 27398
rect 24588 27368 24590 27388
rect 24612 27368 24614 27388
rect 24660 27368 24662 27388
rect 24708 27368 24710 27388
rect 24732 27368 24734 27388
rect 24756 27368 24758 27388
rect 24828 27368 24830 27390
rect 24852 27368 24854 27388
rect 24876 27368 24878 27388
rect 24948 27368 24950 27390
rect 25034 27388 25036 27398
rect 24972 27368 24974 27388
rect 24996 27368 24998 27388
rect 25044 27368 25046 27388
rect 25092 27368 25094 27388
rect 25140 27368 25142 27390
rect 25260 27368 25262 27388
rect 25356 27368 25358 27388
rect 25380 27368 25382 27388
rect 25452 27368 25454 27388
rect 25476 27368 25478 27388
rect 25500 27368 25502 27388
rect 25548 27368 25550 27390
rect 25634 27388 25636 27398
rect 25572 27368 25574 27388
rect 25596 27368 25598 27388
rect 25644 27368 25646 27388
rect 26241 27368 26275 27370
rect 26865 27368 26899 27370
rect 27060 27368 27062 27388
rect 27108 27368 27110 27388
rect 27180 27368 27182 27388
rect 27276 27368 27278 27390
rect 27324 27368 27326 27388
rect 27372 27368 27374 27456
rect 32017 27445 32020 27450
rect 32089 27446 32093 27454
rect 32079 27440 32089 27446
rect 32102 27440 32103 27443
rect 28273 27435 28286 27440
rect 28296 27435 28307 27440
rect 32041 27435 32054 27440
rect 32064 27435 32075 27440
rect 32089 27433 32123 27440
rect 32089 27432 32093 27433
rect 32102 27432 32103 27433
rect 27458 27388 27460 27398
rect 27396 27368 27398 27388
rect 27420 27368 27422 27388
rect 27468 27368 27470 27388
rect 27516 27368 27518 27390
rect 30482 27388 30484 27398
rect 30530 27388 30532 27398
rect 27540 27368 27542 27388
rect 27564 27368 27566 27388
rect 28190 27368 28224 27370
rect 28910 27368 28944 27370
rect 29630 27368 29664 27370
rect 30350 27368 30384 27370
rect 30492 27368 30494 27388
rect 30540 27368 30542 27388
rect 30612 27368 30614 27390
rect 30698 27388 30700 27398
rect 30636 27368 30638 27388
rect 30660 27368 30662 27388
rect 30708 27368 30710 27388
rect 30756 27368 30758 27390
rect 30842 27388 30844 27398
rect 30780 27368 30782 27388
rect 30804 27368 30806 27388
rect 30852 27368 30854 27388
rect 30900 27368 30902 27390
rect 30986 27388 30988 27398
rect 30924 27368 30926 27388
rect 30948 27368 30950 27388
rect 30996 27368 30998 27388
rect 31044 27368 31046 27390
rect 31130 27388 31132 27398
rect 31068 27368 31070 27388
rect 31092 27368 31094 27388
rect 31140 27368 31142 27388
rect 31188 27368 31190 27388
rect 31236 27368 31238 27388
rect 31857 27368 31891 27370
rect 32076 27368 32078 27388
rect 32100 27368 32102 27390
rect 32138 27388 32140 27398
rect 32148 27368 32150 27388
rect -19052 27363 32194 27368
rect -17916 27345 -17914 27363
rect -17868 27345 -17866 27363
rect -17820 27345 -17818 27363
rect -17772 27345 -17770 27363
rect -17652 27345 -17650 27363
rect -17532 27345 -17530 27363
rect -17436 27345 -17434 27363
rect -17412 27345 -17410 27363
rect -17364 27345 -17362 27363
rect -17316 27345 -17314 27363
rect -17220 27345 -17218 27363
rect -17196 27345 -17194 27363
rect -17124 27345 -17122 27363
rect -17028 27345 -17026 27363
rect -16980 27345 -16978 27363
rect -16884 27345 -16882 27363
rect -16860 27345 -16858 27363
rect -16812 27345 -16810 27363
rect -16788 27345 -16786 27363
rect -16764 27345 -16762 27363
rect -16716 27345 -16714 27363
rect -16692 27345 -16690 27363
rect -16668 27345 -16666 27363
rect -16596 27345 -16594 27363
rect -16500 27345 -16498 27363
rect -16404 27345 -16402 27363
rect -16380 27345 -16378 27363
rect -16332 27345 -16330 27363
rect -16308 27345 -16306 27363
rect -16284 27345 -16282 27363
rect -16236 27345 -16234 27363
rect -16212 27345 -16210 27363
rect -16188 27345 -16186 27363
rect -15769 27360 -15753 27363
rect -15809 27345 -15773 27348
rect -15560 27346 -15557 27363
rect -15560 27345 -15558 27346
rect -15420 27345 -15418 27363
rect -15396 27345 -15394 27363
rect -15372 27345 -15370 27363
rect -15300 27345 -15298 27363
rect -15084 27345 -15082 27363
rect -15036 27345 -15034 27363
rect -14940 27345 -14938 27363
rect -14916 27345 -14914 27363
rect -14868 27345 -14866 27363
rect -14820 27345 -14818 27363
rect -14724 27345 -14722 27363
rect -14700 27345 -14698 27363
rect -14652 27345 -14650 27363
rect -14604 27345 -14602 27363
rect -14508 27345 -14506 27363
rect -14484 27345 -14482 27363
rect -14436 27345 -14434 27363
rect -14388 27345 -14386 27363
rect -14268 27345 -14266 27363
rect -14172 27345 -14170 27363
rect -14076 27345 -14074 27363
rect -14028 27345 -14026 27363
rect -13980 27345 -13978 27363
rect -13956 27345 -13954 27363
rect -13932 27345 -13930 27363
rect -13860 27345 -13858 27363
rect -13764 27345 -13762 27363
rect -13716 27345 -13714 27363
rect -13644 27345 -13642 27363
rect -13596 27345 -13594 27363
rect -13500 27345 -13498 27363
rect -13404 27345 -13402 27363
rect -13356 27345 -13354 27363
rect -13284 27345 -13282 27363
rect -12828 27345 -12826 27363
rect -12780 27345 -12778 27363
rect -12684 27345 -12682 27363
rect -12660 27345 -12658 27363
rect -12612 27345 -12610 27363
rect -12588 27345 -12586 27363
rect -12564 27345 -12562 27363
rect -12492 27345 -12490 27363
rect -12396 27345 -12394 27363
rect -12348 27345 -12346 27363
rect -12276 27345 -12274 27363
rect -12252 27345 -12250 27363
rect -12228 27345 -12226 27363
rect -12156 27345 -12154 27363
rect -12060 27345 -12058 27363
rect -12012 27345 -12010 27363
rect -11916 27345 -11914 27363
rect -11892 27345 -11890 27363
rect -11844 27345 -11842 27363
rect -11796 27345 -11794 27363
rect -11676 27345 -11674 27363
rect -11580 27345 -11578 27363
rect -11556 27345 -11554 27363
rect -11484 27345 -11482 27363
rect -11460 27345 -11458 27363
rect -11436 27345 -11434 27363
rect -11388 27345 -11386 27363
rect -11364 27345 -11362 27363
rect -11340 27345 -11338 27363
rect -11268 27345 -11266 27363
rect -11172 27345 -11170 27363
rect -11124 27345 -11122 27363
rect -11076 27345 -11074 27363
rect -11028 27345 -11026 27363
rect -10932 27345 -10930 27363
rect -10836 27345 -10834 27363
rect -10788 27345 -10786 27363
rect -10668 27345 -10666 27363
rect -10225 27360 -10209 27363
rect -10265 27345 -10229 27348
rect -10016 27346 -10013 27363
rect -10016 27345 -10014 27346
rect -9876 27345 -9874 27363
rect -9828 27345 -9826 27363
rect -9732 27345 -9730 27363
rect -9708 27345 -9706 27363
rect -9612 27345 -9610 27363
rect -9516 27345 -9514 27363
rect -9468 27345 -9466 27363
rect -9420 27345 -9418 27363
rect -9396 27345 -9394 27363
rect -9372 27345 -9370 27363
rect -9300 27345 -9298 27363
rect -9252 27345 -9250 27363
rect -9156 27345 -9154 27363
rect -9132 27345 -9130 27363
rect -9084 27345 -9082 27363
rect -9060 27345 -9058 27363
rect -9036 27345 -9034 27363
rect -8988 27345 -8986 27363
rect -8964 27345 -8962 27363
rect -8940 27345 -8938 27363
rect -8892 27345 -8890 27363
rect -8844 27345 -8842 27363
rect -8796 27345 -8794 27363
rect -8700 27345 -8698 27363
rect -8604 27345 -8602 27363
rect -8556 27345 -8554 27363
rect -8508 27345 -8506 27363
rect -8484 27345 -8482 27363
rect -8460 27345 -8458 27363
rect -8412 27345 -8410 27363
rect -8388 27345 -8386 27363
rect -8364 27345 -8362 27363
rect -8316 27345 -8314 27363
rect -8292 27345 -8290 27363
rect -8268 27345 -8266 27363
rect -8196 27345 -8194 27363
rect -8100 27345 -8098 27363
rect -8052 27345 -8050 27363
rect -7932 27345 -7930 27363
rect -7836 27345 -7834 27363
rect -7740 27345 -7738 27363
rect -7692 27345 -7690 27363
rect -7620 27345 -7618 27363
rect -7356 27345 -7354 27363
rect -7284 27345 -7282 27363
rect -7212 27345 -7210 27363
rect -7188 27345 -7186 27363
rect -7116 27345 -7114 27363
rect -7092 27345 -7090 27363
rect -7068 27345 -7066 27363
rect -6996 27345 -6994 27363
rect -6972 27345 -6970 27363
rect -6948 27345 -6946 27363
rect -6900 27345 -6898 27363
rect -6876 27345 -6874 27363
rect -6852 27345 -6850 27363
rect -6804 27345 -6802 27363
rect -6780 27345 -6778 27363
rect -6756 27345 -6754 27363
rect -6708 27345 -6706 27363
rect -6684 27345 -6682 27363
rect -6660 27345 -6658 27363
rect -6612 27345 -6610 27363
rect -6588 27345 -6586 27363
rect -6564 27345 -6562 27363
rect -6516 27345 -6514 27363
rect -6492 27345 -6490 27363
rect -6468 27345 -6466 27363
rect -6420 27345 -6418 27363
rect -6396 27345 -6394 27363
rect -6372 27345 -6370 27363
rect -6324 27345 -6322 27363
rect -6300 27345 -6298 27363
rect -6276 27345 -6274 27363
rect -6228 27345 -6226 27363
rect -6180 27345 -6178 27363
rect -6060 27345 -6058 27363
rect -5964 27345 -5962 27363
rect -5940 27345 -5938 27363
rect -5868 27345 -5866 27363
rect -5796 27345 -5794 27363
rect -5652 27345 -5650 27363
rect -5316 27345 -5314 27363
rect -5268 27345 -5266 27363
rect -5220 27345 -5218 27363
rect -5196 27345 -5194 27363
rect -5172 27345 -5170 27363
rect -5124 27345 -5122 27363
rect -5100 27345 -5098 27363
rect -5076 27345 -5074 27363
rect -5028 27345 -5026 27363
rect -4980 27345 -4978 27363
rect -4884 27345 -4882 27363
rect -4860 27345 -4858 27363
rect -4788 27345 -4786 27363
rect -4692 27345 -4690 27363
rect -4644 27345 -4642 27363
rect -4596 27345 -4594 27363
rect -4548 27345 -4546 27363
rect -4428 27345 -4426 27363
rect -4332 27345 -4330 27363
rect -4308 27345 -4306 27363
rect -4260 27345 -4258 27363
rect -4212 27345 -4210 27363
rect -4116 27345 -4114 27363
rect -4092 27345 -4090 27363
rect -4020 27345 -4018 27363
rect -3876 27345 -3874 27363
rect -3804 27345 -3802 27363
rect -3732 27345 -3730 27363
rect -3588 27345 -3586 27363
rect -3564 27345 -3562 27363
rect -3516 27345 -3514 27363
rect -3492 27345 -3490 27363
rect -3468 27345 -3466 27363
rect -3420 27345 -3418 27363
rect -3372 27345 -3370 27363
rect -3252 27345 -3250 27363
rect -3156 27345 -3154 27363
rect -3132 27345 -3130 27363
rect -3060 27345 -3058 27363
rect -3012 27345 -3010 27363
rect -2916 27345 -2914 27363
rect -2892 27345 -2890 27363
rect -2844 27345 -2842 27363
rect -2820 27345 -2818 27363
rect -2796 27345 -2794 27363
rect -2748 27345 -2746 27363
rect -2700 27345 -2698 27363
rect -2604 27345 -2602 27363
rect -2580 27345 -2578 27363
rect -2508 27345 -2506 27363
rect -2412 27345 -2410 27363
rect -2364 27345 -2362 27363
rect -2292 27345 -2290 27363
rect -2268 27345 -2266 27363
rect -2244 27345 -2242 27363
rect -2196 27345 -2194 27363
rect -2172 27345 -2170 27363
rect -2148 27345 -2146 27363
rect -2100 27345 -2098 27363
rect -2076 27345 -2074 27363
rect -2052 27345 -2050 27363
rect -1980 27345 -1978 27363
rect -1884 27345 -1882 27363
rect -1836 27345 -1834 27363
rect -1716 27345 -1714 27363
rect -1596 27345 -1594 27363
rect -1476 27345 -1474 27363
rect -1380 27345 -1378 27363
rect -1356 27345 -1354 27363
rect -1308 27345 -1306 27363
rect -1260 27345 -1258 27363
rect -1164 27345 -1162 27363
rect -1140 27345 -1138 27363
rect -1068 27345 -1066 27363
rect -852 27345 -850 27363
rect -804 27345 -802 27363
rect -756 27345 -754 27363
rect -708 27345 -706 27363
rect -612 27345 -610 27363
rect -588 27345 -586 27363
rect -540 27345 -538 27363
rect -516 27345 -514 27363
rect -492 27345 -490 27363
rect -444 27345 -442 27363
rect -396 27345 -394 27363
rect -300 27345 -298 27363
rect -276 27345 -274 27363
rect -204 27345 -202 27363
rect -108 27345 -106 27363
rect -60 27345 -58 27363
rect 12 27345 14 27363
rect 108 27345 110 27363
rect 156 27345 158 27363
rect 204 27345 206 27363
rect 228 27345 230 27363
rect 252 27345 254 27363
rect 300 27345 302 27363
rect 348 27345 350 27363
rect 468 27345 470 27363
rect 564 27345 566 27363
rect 588 27345 590 27363
rect 636 27345 638 27363
rect 660 27345 662 27363
rect 684 27345 686 27363
rect 732 27345 734 27363
rect 756 27345 758 27363
rect 780 27345 782 27363
rect 876 27345 878 27363
rect 972 27345 974 27363
rect 1020 27345 1022 27363
rect 1068 27345 1070 27363
rect 1092 27345 1094 27363
rect 1116 27345 1118 27363
rect 1164 27345 1166 27363
rect 1212 27345 1214 27363
rect 1308 27345 1310 27363
rect 1332 27345 1334 27363
rect 1380 27345 1382 27363
rect 1428 27345 1430 27363
rect 1524 27345 1526 27363
rect 1548 27345 1550 27363
rect 1596 27345 1598 27363
rect 1620 27345 1622 27363
rect 1644 27345 1646 27363
rect 1692 27345 1694 27363
rect 1716 27345 1718 27363
rect 1740 27345 1742 27363
rect 1788 27345 1790 27363
rect 1812 27345 1814 27363
rect 1836 27345 1838 27363
rect 1884 27345 1886 27363
rect 1908 27345 1910 27363
rect 1932 27345 1934 27363
rect 1980 27345 1982 27363
rect 2004 27345 2006 27363
rect 2028 27345 2030 27363
rect 2076 27345 2078 27363
rect 2100 27345 2102 27363
rect 2124 27345 2126 27363
rect 2172 27345 2174 27363
rect 2196 27345 2198 27363
rect 2220 27345 2222 27363
rect 2268 27345 2270 27363
rect 2292 27345 2294 27363
rect 2316 27345 2318 27363
rect 2364 27345 2366 27363
rect 2388 27345 2390 27363
rect 2412 27345 2414 27363
rect 2460 27345 2462 27363
rect 2484 27345 2486 27363
rect 2508 27345 2510 27363
rect 2556 27345 2558 27363
rect 2580 27345 2582 27363
rect 2604 27345 2606 27363
rect 2652 27345 2654 27363
rect 2676 27345 2678 27363
rect 2700 27345 2702 27363
rect 2748 27345 2750 27363
rect 2772 27345 2774 27363
rect 2796 27345 2798 27363
rect 2844 27345 2846 27363
rect 2868 27345 2870 27363
rect 2892 27345 2894 27363
rect 2940 27345 2942 27363
rect 3012 27345 3014 27363
rect 3108 27345 3110 27363
rect 3156 27345 3158 27363
rect 3252 27345 3254 27363
rect 3348 27345 3350 27363
rect 3396 27345 3398 27363
rect 3468 27345 3470 27363
rect 3492 27345 3494 27363
rect 3516 27345 3518 27363
rect 3588 27345 3590 27363
rect 3612 27345 3614 27363
rect 3636 27345 3638 27363
rect 3708 27345 3710 27363
rect 3732 27345 3734 27363
rect 3756 27345 3758 27363
rect 3804 27345 3806 27363
rect 3828 27345 3830 27363
rect 3852 27345 3854 27363
rect 3900 27345 3902 27363
rect 3924 27345 3926 27363
rect 3948 27345 3950 27363
rect 3996 27345 3998 27363
rect 4020 27345 4022 27363
rect 4044 27345 4046 27363
rect 4092 27345 4094 27363
rect 4116 27345 4118 27363
rect 4140 27345 4142 27363
rect 4188 27345 4190 27363
rect 4212 27345 4214 27363
rect 4236 27345 4238 27363
rect 4284 27345 4286 27363
rect 4308 27345 4310 27363
rect 4332 27345 4334 27363
rect 4380 27345 4382 27363
rect 4404 27345 4406 27363
rect 4428 27345 4430 27363
rect 4476 27345 4478 27363
rect 4500 27345 4502 27363
rect 4524 27345 4526 27363
rect 4596 27345 4598 27363
rect 4812 27345 4814 27363
rect 4860 27345 4862 27363
rect 4908 27345 4910 27363
rect 4956 27345 4958 27363
rect 4980 27345 4982 27363
rect 5004 27345 5006 27363
rect 5076 27345 5078 27363
rect 5100 27345 5102 27363
rect 5124 27345 5126 27363
rect 5172 27345 5174 27363
rect 5196 27345 5198 27363
rect 5220 27345 5222 27363
rect 5268 27345 5270 27363
rect 5292 27345 5294 27363
rect 5316 27345 5318 27363
rect 5388 27345 5390 27363
rect 5412 27345 5414 27363
rect 5436 27345 5438 27363
rect 5484 27345 5486 27363
rect 5508 27345 5510 27363
rect 5532 27345 5534 27363
rect 5580 27345 5582 27363
rect 5628 27345 5630 27363
rect 5724 27345 5726 27363
rect 5748 27345 5750 27363
rect 5796 27345 5798 27363
rect 5820 27345 5822 27363
rect 5844 27345 5846 27363
rect 5916 27345 5918 27363
rect 6132 27345 6134 27363
rect 6180 27345 6182 27363
rect 6228 27345 6230 27363
rect 6252 27345 6254 27363
rect 6276 27345 6278 27363
rect 6324 27345 6326 27363
rect 6372 27345 6374 27363
rect 6468 27345 6470 27363
rect 6492 27345 6494 27363
rect 6564 27345 6566 27363
rect 6588 27345 6590 27363
rect 6612 27345 6614 27363
rect 6660 27345 6662 27363
rect 6684 27345 6686 27363
rect 6708 27345 6710 27363
rect 6780 27345 6782 27363
rect 6804 27345 6806 27363
rect 6828 27345 6830 27363
rect 6876 27345 6878 27363
rect 6900 27345 6902 27363
rect 6924 27345 6926 27363
rect 6972 27345 6974 27363
rect 7020 27345 7022 27363
rect 7140 27345 7142 27363
rect 7236 27345 7238 27363
rect 7260 27345 7262 27363
rect 7332 27345 7334 27363
rect 7356 27345 7358 27363
rect 7380 27345 7382 27363
rect 7428 27345 7430 27363
rect 7452 27345 7454 27363
rect 7476 27345 7478 27363
rect 7524 27345 7526 27363
rect 7548 27345 7550 27363
rect 7572 27345 7574 27363
rect 7620 27345 7622 27363
rect 7644 27345 7646 27363
rect 7668 27345 7670 27363
rect 7716 27345 7718 27363
rect 7740 27345 7742 27363
rect 7764 27345 7766 27363
rect 7836 27345 7838 27363
rect 7860 27345 7862 27363
rect 7884 27345 7886 27363
rect 7932 27345 7934 27363
rect 7956 27345 7958 27363
rect 7980 27345 7982 27363
rect 8052 27345 8054 27363
rect 8148 27345 8150 27363
rect 8196 27345 8198 27363
rect 8244 27345 8246 27363
rect 8268 27345 8270 27363
rect 8292 27345 8294 27363
rect 8340 27345 8342 27363
rect 8364 27345 8366 27363
rect 8388 27345 8390 27363
rect 8436 27345 8438 27363
rect 8460 27345 8462 27363
rect 8484 27345 8486 27363
rect 8556 27345 8558 27363
rect 8580 27345 8582 27363
rect 8604 27345 8606 27363
rect 8676 27345 8678 27363
rect 8700 27345 8702 27363
rect 8724 27345 8726 27363
rect 8772 27345 8774 27363
rect 8820 27345 8822 27363
rect 8844 27345 8846 27363
rect 8868 27345 8870 27363
rect 9287 27360 9303 27363
rect 9247 27345 9283 27348
rect 9496 27346 9499 27363
rect 9496 27345 9498 27346
rect 9660 27345 9662 27363
rect 9684 27345 9686 27363
rect 9708 27345 9710 27363
rect 9756 27345 9758 27363
rect 9780 27345 9782 27363
rect 9804 27345 9806 27363
rect 9852 27345 9854 27363
rect 9876 27345 9878 27363
rect 9900 27345 9902 27363
rect 9948 27345 9950 27363
rect 9972 27345 9974 27363
rect 9996 27345 9998 27363
rect 10068 27345 10070 27363
rect 10092 27345 10094 27363
rect 10116 27345 10118 27363
rect 10164 27345 10166 27363
rect 10188 27345 10190 27363
rect 10212 27345 10214 27363
rect 10260 27345 10262 27363
rect 10284 27345 10286 27363
rect 10308 27345 10310 27363
rect 10380 27345 10382 27363
rect 10404 27345 10406 27363
rect 10428 27345 10430 27363
rect 10476 27345 10478 27363
rect 10500 27345 10502 27363
rect 10524 27345 10526 27363
rect 10572 27345 10574 27363
rect 10596 27345 10598 27363
rect 10620 27345 10622 27363
rect 10668 27345 10670 27363
rect 10692 27345 10694 27363
rect 10716 27345 10718 27363
rect 10788 27345 10790 27363
rect 10836 27345 10838 27363
rect 10956 27345 10958 27363
rect 11052 27345 11054 27363
rect 11076 27345 11078 27363
rect 11124 27345 11126 27363
rect 11172 27345 11174 27363
rect 11220 27345 11222 27363
rect 11340 27345 11342 27363
rect 11436 27345 11438 27363
rect 11532 27345 11534 27363
rect 11580 27345 11582 27363
rect 11628 27345 11630 27363
rect 11652 27345 11654 27363
rect 11676 27345 11678 27363
rect 11748 27345 11750 27363
rect 11772 27345 11774 27363
rect 11796 27345 11798 27363
rect 11844 27345 11846 27363
rect 11892 27345 11894 27363
rect 11988 27345 11990 27363
rect 12012 27345 12014 27363
rect 12084 27345 12086 27363
rect 12132 27345 12134 27363
rect 12228 27345 12230 27363
rect 12252 27345 12254 27363
rect 12300 27345 12302 27363
rect 12324 27345 12326 27363
rect 12348 27345 12350 27363
rect 12396 27345 12398 27363
rect 12420 27345 12422 27363
rect 12444 27345 12446 27363
rect 12492 27345 12494 27363
rect 12516 27345 12518 27363
rect 12540 27345 12542 27363
rect 12588 27345 12590 27363
rect 12636 27345 12638 27363
rect 12732 27345 12734 27363
rect 12756 27345 12758 27363
rect 12804 27345 12806 27363
rect 12828 27345 12830 27363
rect 12852 27345 12854 27363
rect 12900 27345 12902 27363
rect 12924 27345 12926 27363
rect 12948 27345 12950 27363
rect 13020 27345 13022 27363
rect 13044 27345 13046 27363
rect 13068 27345 13070 27363
rect 13116 27345 13118 27363
rect 13188 27345 13190 27363
rect 13284 27345 13286 27363
rect 13332 27345 13334 27363
rect 13428 27345 13430 27363
rect 13524 27345 13526 27363
rect 13572 27345 13574 27363
rect 13644 27345 13646 27363
rect 13668 27345 13670 27363
rect 13692 27345 13694 27363
rect 13764 27345 13766 27363
rect 13788 27345 13790 27363
rect 13812 27345 13814 27363
rect 13860 27345 13862 27363
rect 13884 27345 13886 27363
rect 13908 27345 13910 27363
rect 13956 27345 13958 27363
rect 14004 27345 14006 27363
rect 14100 27345 14102 27363
rect 14196 27345 14198 27363
rect 14244 27345 14246 27363
rect 14292 27345 14294 27363
rect 14711 27360 14727 27363
rect 14671 27345 14707 27348
rect 14920 27346 14923 27363
rect 14920 27345 14922 27346
rect 15132 27345 15134 27363
rect 15228 27345 15230 27363
rect 15252 27345 15254 27363
rect 15300 27345 15302 27363
rect 15324 27345 15326 27363
rect 15348 27345 15350 27363
rect 15396 27345 15398 27363
rect 15420 27345 15422 27363
rect 15444 27345 15446 27363
rect 15492 27345 15494 27363
rect 15540 27345 15542 27363
rect 15636 27345 15638 27363
rect 15660 27345 15662 27363
rect 15708 27345 15710 27363
rect 15732 27345 15734 27363
rect 15756 27345 15758 27363
rect 15804 27345 15806 27363
rect 15828 27345 15830 27363
rect 15852 27345 15854 27363
rect 15900 27345 15902 27363
rect 15924 27345 15926 27363
rect 15948 27345 15950 27363
rect 15996 27345 15998 27363
rect 16020 27345 16022 27363
rect 16044 27345 16046 27363
rect 16092 27345 16094 27363
rect 16140 27345 16142 27363
rect 16236 27345 16238 27363
rect 16260 27345 16262 27363
rect 16308 27345 16310 27363
rect 16332 27345 16334 27363
rect 16356 27345 16358 27363
rect 16404 27345 16406 27363
rect 16452 27345 16454 27363
rect 16548 27345 16550 27363
rect 16572 27345 16574 27363
rect 16620 27345 16622 27363
rect 16644 27345 16646 27363
rect 16668 27345 16670 27363
rect 16716 27345 16718 27363
rect 16740 27345 16742 27363
rect 16764 27345 16766 27363
rect 16836 27345 16838 27363
rect 16884 27345 16886 27363
rect 16980 27345 16982 27363
rect 17004 27345 17006 27363
rect 17052 27345 17054 27363
rect 17100 27345 17102 27363
rect 17196 27345 17198 27363
rect 17220 27345 17222 27363
rect 17268 27345 17270 27363
rect 17292 27345 17294 27363
rect 17316 27345 17318 27363
rect 17735 27360 17751 27363
rect 17695 27345 17731 27348
rect 17944 27346 17947 27363
rect 17944 27345 17946 27346
rect 18084 27345 18086 27363
rect 18108 27345 18110 27363
rect 18132 27345 18134 27363
rect 18180 27345 18182 27363
rect 18252 27345 18254 27363
rect 18348 27345 18350 27363
rect 18396 27345 18398 27363
rect 18492 27345 18494 27363
rect 18516 27345 18518 27363
rect 18564 27345 18566 27363
rect 18588 27345 18590 27363
rect 18612 27345 18614 27363
rect 18660 27345 18662 27363
rect 18684 27345 18686 27363
rect 18708 27345 18710 27363
rect 18756 27345 18758 27363
rect 18780 27345 18782 27363
rect 18804 27345 18806 27363
rect 18852 27345 18854 27363
rect 18876 27345 18878 27363
rect 18900 27345 18902 27363
rect 18948 27345 18950 27363
rect 18996 27345 18998 27363
rect 19020 27345 19022 27363
rect 19044 27345 19046 27363
rect 19092 27345 19094 27363
rect 19116 27345 19118 27363
rect 19140 27345 19142 27363
rect 19188 27345 19190 27363
rect 19236 27345 19238 27363
rect 19332 27345 19334 27363
rect 19428 27345 19430 27363
rect 19476 27345 19478 27363
rect 19524 27345 19526 27363
rect 19572 27345 19574 27363
rect 19596 27345 19598 27363
rect 19620 27345 19622 27363
rect 19668 27345 19670 27363
rect 19692 27345 19694 27363
rect 19716 27345 19718 27363
rect 19764 27345 19766 27363
rect 19812 27345 19814 27363
rect 19836 27345 19838 27363
rect 19860 27345 19862 27363
rect 19932 27345 19934 27363
rect 19956 27345 19958 27363
rect 19980 27345 19982 27363
rect 20028 27345 20030 27363
rect 20052 27345 20054 27363
rect 20076 27345 20078 27363
rect 20148 27345 20150 27363
rect 20172 27345 20174 27363
rect 20196 27345 20198 27363
rect 20244 27345 20246 27363
rect 20268 27345 20270 27363
rect 20292 27345 20294 27363
rect 20340 27345 20342 27363
rect 20388 27345 20390 27363
rect 20484 27345 20486 27363
rect 20508 27345 20510 27363
rect 20556 27345 20558 27363
rect 20580 27345 20582 27363
rect 20604 27345 20606 27363
rect 20700 27345 20702 27363
rect 20916 27345 20918 27363
rect 20964 27345 20966 27363
rect 21012 27345 21014 27363
rect 21060 27345 21062 27363
rect 21084 27345 21086 27363
rect 21108 27345 21110 27363
rect 21156 27345 21158 27363
rect 21204 27345 21206 27363
rect 21300 27345 21302 27363
rect 21324 27345 21326 27363
rect 21372 27345 21374 27363
rect 21420 27345 21422 27363
rect 21444 27345 21446 27363
rect 21468 27345 21470 27363
rect 21516 27345 21518 27363
rect 21540 27345 21542 27363
rect 21564 27345 21566 27363
rect 21612 27345 21614 27363
rect 21660 27345 21662 27363
rect 21684 27345 21686 27363
rect 21708 27345 21710 27363
rect 21780 27345 21782 27363
rect 21804 27345 21806 27363
rect 21828 27345 21830 27363
rect 21900 27345 21902 27363
rect 21924 27345 21926 27363
rect 21948 27345 21950 27363
rect 22020 27345 22022 27363
rect 22044 27345 22046 27363
rect 22068 27345 22070 27363
rect 22116 27345 22118 27363
rect 22164 27345 22166 27363
rect 22188 27345 22190 27363
rect 22212 27345 22214 27363
rect 22655 27360 22671 27363
rect 22615 27345 22651 27348
rect 22864 27346 22867 27363
rect 22864 27345 22866 27346
rect 23004 27345 23006 27363
rect 23052 27345 23054 27363
rect 23076 27345 23078 27363
rect 23100 27345 23102 27363
rect 23148 27345 23150 27363
rect 23196 27345 23198 27363
rect 23220 27345 23222 27363
rect 23244 27345 23246 27363
rect 23292 27345 23294 27363
rect 23316 27345 23318 27363
rect 23340 27345 23342 27363
rect 23388 27345 23390 27363
rect 23412 27345 23414 27363
rect 23436 27345 23438 27363
rect 23484 27345 23486 27363
rect 23532 27345 23534 27363
rect 23556 27345 23558 27363
rect 23580 27345 23582 27363
rect 23628 27345 23630 27363
rect 23652 27345 23654 27363
rect 23676 27345 23678 27363
rect 23724 27345 23726 27363
rect 23748 27345 23750 27363
rect 23772 27345 23774 27363
rect 23820 27345 23822 27363
rect 23868 27345 23870 27363
rect 23892 27345 23894 27363
rect 23916 27345 23918 27363
rect 23988 27345 23990 27363
rect 24012 27345 24014 27363
rect 24036 27345 24038 27363
rect 24084 27345 24086 27363
rect 24132 27345 24134 27363
rect 24228 27345 24230 27363
rect 24252 27345 24254 27363
rect 24300 27345 24302 27363
rect 24348 27345 24350 27363
rect 24372 27345 24374 27363
rect 24396 27345 24398 27363
rect 24468 27345 24470 27363
rect 24492 27345 24494 27363
rect 24516 27345 24518 27363
rect 24564 27345 24566 27363
rect 24588 27345 24590 27363
rect 24612 27345 24614 27363
rect 24660 27345 24662 27363
rect 24708 27345 24710 27363
rect 24732 27345 24734 27363
rect 24756 27345 24758 27363
rect 24828 27345 24830 27363
rect 24852 27345 24854 27363
rect 24876 27345 24878 27363
rect 24948 27345 24950 27363
rect 24972 27345 24974 27363
rect 24996 27345 24998 27363
rect 25044 27345 25046 27363
rect 25092 27345 25094 27363
rect 25140 27345 25142 27363
rect 25260 27345 25262 27363
rect 25356 27345 25358 27363
rect 25380 27345 25382 27363
rect 25452 27345 25454 27363
rect 25476 27345 25478 27363
rect 25500 27345 25502 27363
rect 25548 27345 25550 27363
rect 25572 27345 25574 27363
rect 25596 27345 25598 27363
rect 25644 27345 25646 27363
rect 26063 27360 26079 27363
rect 26023 27345 26059 27348
rect 26272 27346 26275 27363
rect 26687 27360 26703 27363
rect 26272 27345 26274 27346
rect 26647 27345 26683 27348
rect 26896 27346 26899 27363
rect 26896 27345 26898 27346
rect 27060 27345 27062 27363
rect 27108 27345 27110 27363
rect 27180 27345 27182 27363
rect 27276 27345 27278 27363
rect 27324 27345 27326 27363
rect 27372 27345 27374 27363
rect 27396 27345 27398 27363
rect 27420 27345 27422 27363
rect 27468 27345 27470 27363
rect 27516 27345 27518 27363
rect 27540 27345 27542 27363
rect 27564 27345 27566 27363
rect 27983 27360 27999 27363
rect 28703 27360 28719 27363
rect 29423 27360 29439 27363
rect 30143 27360 30159 27363
rect 27943 27345 27979 27348
rect 28663 27345 28699 27348
rect 29383 27345 29419 27348
rect 30103 27345 30139 27348
rect 30492 27345 30494 27363
rect 30540 27345 30542 27363
rect 30612 27345 30614 27363
rect 30636 27345 30638 27363
rect 30660 27345 30662 27363
rect 30708 27345 30710 27363
rect 30756 27345 30758 27363
rect 30780 27345 30782 27363
rect 30804 27345 30806 27363
rect 30852 27345 30854 27363
rect 30900 27345 30902 27363
rect 30924 27345 30926 27363
rect 30948 27345 30950 27363
rect 30996 27345 30998 27363
rect 31044 27345 31046 27363
rect 31068 27345 31070 27363
rect 31092 27345 31094 27363
rect 31140 27345 31142 27363
rect 31188 27345 31190 27363
rect 31236 27345 31238 27363
rect 31679 27360 31695 27363
rect 31639 27345 31675 27348
rect 31888 27346 31891 27363
rect 31888 27345 31890 27346
rect 32076 27345 32078 27363
rect 32100 27345 32102 27363
rect 32148 27345 32150 27363
rect -19052 27340 32194 27345
rect -17916 27322 -17914 27340
rect -17868 27322 -17866 27340
rect -17820 27322 -17818 27340
rect -17772 27322 -17770 27340
rect -17652 27322 -17650 27340
rect -17532 27322 -17530 27340
rect -17436 27322 -17434 27340
rect -17412 27322 -17410 27340
rect -17364 27322 -17362 27340
rect -17316 27322 -17314 27340
rect -17220 27322 -17218 27340
rect -17196 27322 -17194 27340
rect -17124 27322 -17122 27340
rect -17028 27322 -17026 27340
rect -16980 27322 -16978 27340
rect -16884 27322 -16882 27340
rect -16860 27322 -16858 27340
rect -16812 27322 -16810 27340
rect -16788 27322 -16786 27340
rect -16764 27322 -16762 27340
rect -16716 27322 -16714 27340
rect -16692 27322 -16690 27340
rect -16668 27322 -16666 27340
rect -16596 27322 -16594 27340
rect -16500 27322 -16498 27340
rect -16404 27322 -16402 27340
rect -16380 27322 -16378 27340
rect -16332 27322 -16330 27340
rect -16308 27322 -16306 27340
rect -16284 27322 -16282 27340
rect -16236 27322 -16234 27340
rect -16212 27322 -16210 27340
rect -16188 27322 -16186 27340
rect -15560 27322 -15558 27340
rect -15505 27338 -15491 27340
rect -15420 27322 -15418 27340
rect -15396 27322 -15394 27340
rect -15372 27322 -15370 27340
rect -15300 27322 -15298 27340
rect -15084 27322 -15082 27340
rect -15036 27322 -15034 27340
rect -14940 27322 -14938 27340
rect -14916 27322 -14914 27340
rect -14868 27322 -14866 27340
rect -14820 27322 -14818 27340
rect -14724 27322 -14722 27340
rect -14700 27322 -14698 27340
rect -14652 27322 -14650 27340
rect -14604 27322 -14602 27340
rect -14508 27322 -14506 27340
rect -14484 27322 -14482 27340
rect -14436 27322 -14434 27340
rect -14388 27322 -14386 27340
rect -14268 27322 -14266 27340
rect -14172 27322 -14170 27340
rect -14076 27322 -14074 27340
rect -14028 27322 -14026 27340
rect -13980 27322 -13978 27340
rect -13956 27322 -13954 27340
rect -13932 27322 -13930 27340
rect -13860 27322 -13858 27340
rect -13764 27322 -13762 27340
rect -13716 27322 -13714 27340
rect -13644 27322 -13642 27340
rect -13596 27322 -13594 27340
rect -13500 27322 -13498 27340
rect -13404 27322 -13402 27340
rect -13356 27322 -13354 27340
rect -13284 27322 -13282 27340
rect -12828 27322 -12826 27340
rect -12780 27322 -12778 27340
rect -12684 27322 -12682 27340
rect -12660 27322 -12658 27340
rect -12612 27322 -12610 27340
rect -12588 27322 -12586 27340
rect -12564 27322 -12562 27340
rect -12492 27322 -12490 27340
rect -12396 27322 -12394 27340
rect -12348 27322 -12346 27340
rect -12276 27322 -12274 27340
rect -12252 27322 -12250 27340
rect -12228 27322 -12226 27340
rect -12156 27322 -12154 27340
rect -12060 27322 -12058 27340
rect -12012 27322 -12010 27340
rect -11916 27322 -11914 27340
rect -11892 27322 -11890 27340
rect -11844 27322 -11842 27340
rect -11796 27322 -11794 27340
rect -11676 27322 -11674 27340
rect -11580 27322 -11578 27340
rect -11556 27322 -11554 27340
rect -11484 27322 -11482 27340
rect -11460 27322 -11458 27340
rect -11436 27322 -11434 27340
rect -11388 27322 -11386 27340
rect -11364 27322 -11362 27340
rect -11340 27322 -11338 27340
rect -11268 27322 -11266 27340
rect -11172 27322 -11170 27340
rect -11124 27322 -11122 27340
rect -11076 27322 -11074 27340
rect -11028 27322 -11026 27340
rect -10932 27322 -10930 27340
rect -10836 27322 -10834 27340
rect -10788 27322 -10786 27340
rect -10668 27322 -10666 27340
rect -10016 27322 -10014 27340
rect -9961 27338 -9947 27340
rect -9876 27322 -9874 27340
rect -9828 27322 -9826 27340
rect -9732 27322 -9730 27340
rect -9708 27322 -9706 27340
rect -9612 27322 -9610 27340
rect -9516 27322 -9514 27340
rect -9468 27322 -9466 27340
rect -9420 27322 -9418 27340
rect -9396 27322 -9394 27340
rect -9372 27322 -9370 27340
rect -9300 27322 -9298 27340
rect -9252 27322 -9250 27340
rect -9156 27322 -9154 27340
rect -9132 27322 -9130 27340
rect -9084 27322 -9082 27340
rect -9060 27322 -9058 27340
rect -9036 27322 -9034 27340
rect -8988 27322 -8986 27340
rect -8964 27322 -8962 27340
rect -8940 27322 -8938 27340
rect -8892 27322 -8890 27340
rect -8844 27322 -8842 27340
rect -8796 27322 -8794 27340
rect -8700 27322 -8698 27340
rect -8604 27322 -8602 27340
rect -8556 27322 -8554 27340
rect -8508 27322 -8506 27340
rect -8484 27322 -8482 27340
rect -8460 27322 -8458 27340
rect -8412 27322 -8410 27340
rect -8388 27322 -8386 27340
rect -8364 27322 -8362 27340
rect -8316 27322 -8314 27340
rect -8292 27322 -8290 27340
rect -8268 27322 -8266 27340
rect -8196 27322 -8194 27340
rect -8100 27322 -8098 27340
rect -8052 27322 -8050 27340
rect -7932 27322 -7930 27340
rect -7836 27322 -7834 27340
rect -7740 27322 -7738 27340
rect -7692 27322 -7690 27340
rect -7620 27322 -7618 27340
rect -7356 27322 -7354 27340
rect -7284 27322 -7282 27340
rect -7212 27322 -7210 27340
rect -7188 27322 -7186 27340
rect -7116 27322 -7114 27340
rect -7092 27322 -7090 27340
rect -7068 27322 -7066 27340
rect -6996 27322 -6994 27340
rect -6972 27322 -6970 27340
rect -6948 27322 -6946 27340
rect -6900 27322 -6898 27340
rect -6876 27322 -6874 27340
rect -6852 27322 -6850 27340
rect -6804 27322 -6802 27340
rect -6780 27322 -6778 27340
rect -6756 27322 -6754 27340
rect -6708 27322 -6706 27340
rect -6684 27322 -6682 27340
rect -6660 27322 -6658 27340
rect -6612 27322 -6610 27340
rect -6588 27322 -6586 27340
rect -6564 27322 -6562 27340
rect -6516 27322 -6514 27340
rect -6492 27322 -6490 27340
rect -6468 27322 -6466 27340
rect -6420 27322 -6418 27340
rect -6396 27322 -6394 27340
rect -6372 27322 -6370 27340
rect -6324 27322 -6322 27340
rect -6300 27322 -6298 27340
rect -6276 27322 -6274 27340
rect -6228 27322 -6226 27340
rect -6180 27322 -6178 27340
rect -6060 27322 -6058 27340
rect -5964 27322 -5962 27340
rect -5940 27322 -5938 27340
rect -5868 27322 -5866 27340
rect -5796 27322 -5794 27340
rect -5652 27322 -5650 27340
rect -5316 27322 -5314 27340
rect -5268 27322 -5266 27340
rect -5220 27322 -5218 27340
rect -5196 27322 -5194 27340
rect -5172 27322 -5170 27340
rect -5124 27322 -5122 27340
rect -5100 27322 -5098 27340
rect -5076 27322 -5074 27340
rect -5028 27322 -5026 27340
rect -4980 27322 -4978 27340
rect -4884 27322 -4882 27340
rect -4860 27322 -4858 27340
rect -4788 27322 -4786 27340
rect -4692 27322 -4690 27340
rect -4644 27322 -4642 27340
rect -4596 27322 -4594 27340
rect -4548 27322 -4546 27340
rect -4428 27322 -4426 27340
rect -4332 27322 -4330 27340
rect -4308 27322 -4306 27340
rect -4260 27322 -4258 27340
rect -4212 27322 -4210 27340
rect -4116 27322 -4114 27340
rect -4092 27322 -4090 27340
rect -4020 27322 -4018 27340
rect -3876 27322 -3874 27340
rect -3804 27322 -3802 27340
rect -3732 27322 -3730 27340
rect -3588 27322 -3586 27340
rect -3564 27322 -3562 27340
rect -3516 27322 -3514 27340
rect -3492 27322 -3490 27340
rect -3468 27322 -3466 27340
rect -3420 27322 -3418 27340
rect -3372 27322 -3370 27340
rect -3252 27322 -3250 27340
rect -3156 27322 -3154 27340
rect -3132 27322 -3130 27340
rect -3060 27322 -3058 27340
rect -3012 27322 -3010 27340
rect -2916 27322 -2914 27340
rect -2892 27322 -2890 27340
rect -2844 27322 -2842 27340
rect -2820 27322 -2818 27340
rect -2796 27322 -2794 27340
rect -2748 27322 -2746 27340
rect -2700 27322 -2698 27340
rect -2604 27322 -2602 27340
rect -2580 27322 -2578 27340
rect -2508 27322 -2506 27340
rect -2412 27322 -2410 27340
rect -2364 27322 -2362 27340
rect -2292 27322 -2290 27340
rect -2268 27322 -2266 27340
rect -2244 27322 -2242 27340
rect -2196 27322 -2194 27340
rect -2172 27322 -2170 27340
rect -2148 27322 -2146 27340
rect -2100 27322 -2098 27340
rect -2076 27322 -2074 27340
rect -2052 27322 -2050 27340
rect -1980 27322 -1978 27340
rect -1884 27322 -1882 27340
rect -1836 27322 -1834 27340
rect -1716 27322 -1714 27340
rect -1596 27322 -1594 27340
rect -1476 27322 -1474 27340
rect -1380 27322 -1378 27340
rect -1356 27322 -1354 27340
rect -1308 27322 -1306 27340
rect -1260 27322 -1258 27340
rect -1164 27322 -1162 27340
rect -1140 27322 -1138 27340
rect -1068 27322 -1066 27340
rect -852 27322 -850 27340
rect -804 27322 -802 27340
rect -756 27322 -754 27340
rect -708 27322 -706 27340
rect -612 27322 -610 27340
rect -588 27322 -586 27340
rect -540 27322 -538 27340
rect -516 27322 -514 27340
rect -492 27322 -490 27340
rect -444 27322 -442 27340
rect -396 27322 -394 27340
rect -300 27322 -298 27340
rect -276 27322 -274 27340
rect -204 27322 -202 27340
rect -108 27322 -106 27340
rect -60 27322 -58 27340
rect 12 27322 14 27340
rect 108 27322 110 27340
rect 156 27322 158 27340
rect 204 27322 206 27340
rect 228 27322 230 27340
rect 252 27322 254 27340
rect 300 27322 302 27340
rect 348 27322 350 27340
rect 468 27322 470 27340
rect 564 27322 566 27340
rect 588 27322 590 27340
rect 636 27322 638 27340
rect 660 27322 662 27340
rect 684 27322 686 27340
rect 732 27322 734 27340
rect 756 27322 758 27340
rect 780 27322 782 27340
rect 876 27322 878 27340
rect 972 27322 974 27340
rect 1020 27322 1022 27340
rect 1068 27322 1070 27340
rect 1092 27322 1094 27340
rect 1116 27322 1118 27340
rect 1164 27322 1166 27340
rect 1212 27322 1214 27340
rect 1308 27322 1310 27340
rect 1332 27322 1334 27340
rect 1380 27322 1382 27340
rect 1428 27322 1430 27340
rect 1524 27322 1526 27340
rect 1548 27322 1550 27340
rect 1596 27322 1598 27340
rect 1620 27322 1622 27340
rect 1644 27322 1646 27340
rect 1692 27322 1694 27340
rect 1716 27322 1718 27340
rect 1740 27322 1742 27340
rect 1788 27322 1790 27340
rect 1812 27322 1814 27340
rect 1836 27322 1838 27340
rect 1884 27322 1886 27340
rect 1908 27322 1910 27340
rect 1932 27322 1934 27340
rect 1980 27322 1982 27340
rect 2004 27322 2006 27340
rect 2028 27322 2030 27340
rect 2076 27322 2078 27340
rect 2100 27322 2102 27340
rect 2124 27322 2126 27340
rect 2172 27322 2174 27340
rect 2196 27322 2198 27340
rect 2220 27322 2222 27340
rect 2268 27322 2270 27340
rect 2292 27322 2294 27340
rect 2316 27322 2318 27340
rect 2364 27322 2366 27340
rect 2388 27322 2390 27340
rect 2412 27322 2414 27340
rect 2460 27322 2462 27340
rect 2484 27322 2486 27340
rect 2508 27322 2510 27340
rect 2556 27322 2558 27340
rect 2580 27322 2582 27340
rect 2604 27322 2606 27340
rect 2652 27322 2654 27340
rect 2676 27322 2678 27340
rect 2700 27322 2702 27340
rect 2748 27322 2750 27340
rect 2772 27322 2774 27340
rect 2796 27322 2798 27340
rect 2844 27322 2846 27340
rect 2868 27322 2870 27340
rect 2892 27322 2894 27340
rect 2940 27322 2942 27340
rect 3012 27322 3014 27340
rect 3108 27322 3110 27340
rect 3156 27322 3158 27340
rect 3252 27322 3254 27340
rect 3348 27322 3350 27340
rect 3396 27322 3398 27340
rect 3468 27322 3470 27340
rect 3492 27322 3494 27340
rect 3516 27322 3518 27340
rect 3588 27322 3590 27340
rect 3612 27322 3614 27340
rect 3636 27322 3638 27340
rect 3708 27322 3710 27340
rect 3732 27322 3734 27340
rect 3756 27322 3758 27340
rect 3804 27322 3806 27340
rect 3828 27322 3830 27340
rect 3852 27322 3854 27340
rect 3900 27322 3902 27340
rect 3924 27322 3926 27340
rect 3948 27322 3950 27340
rect 3996 27322 3998 27340
rect 4020 27322 4022 27340
rect 4044 27322 4046 27340
rect 4092 27322 4094 27340
rect 4116 27322 4118 27340
rect 4140 27322 4142 27340
rect 4188 27322 4190 27340
rect 4212 27322 4214 27340
rect 4236 27322 4238 27340
rect 4284 27322 4286 27340
rect 4308 27322 4310 27340
rect 4332 27322 4334 27340
rect 4380 27322 4382 27340
rect 4404 27322 4406 27340
rect 4428 27322 4430 27340
rect 4476 27322 4478 27340
rect 4500 27322 4502 27340
rect 4524 27322 4526 27340
rect 4596 27322 4598 27340
rect 4812 27322 4814 27340
rect 4860 27322 4862 27340
rect 4908 27322 4910 27340
rect 4956 27322 4958 27340
rect 4980 27322 4982 27340
rect 5004 27322 5006 27340
rect 5076 27322 5078 27340
rect 5100 27322 5102 27340
rect 5124 27322 5126 27340
rect 5172 27322 5174 27340
rect 5196 27322 5198 27340
rect 5220 27322 5222 27340
rect 5268 27322 5270 27340
rect 5292 27322 5294 27340
rect 5316 27322 5318 27340
rect 5388 27322 5390 27340
rect 5412 27322 5414 27340
rect 5436 27322 5438 27340
rect 5484 27322 5486 27340
rect 5508 27322 5510 27340
rect 5532 27322 5534 27340
rect 5580 27322 5582 27340
rect 5628 27322 5630 27340
rect 5724 27322 5726 27340
rect 5748 27322 5750 27340
rect 5796 27322 5798 27340
rect 5820 27322 5822 27340
rect 5844 27322 5846 27340
rect 5916 27322 5918 27340
rect 6132 27322 6134 27340
rect 6180 27322 6182 27340
rect 6228 27322 6230 27340
rect 6252 27322 6254 27340
rect 6276 27322 6278 27340
rect 6324 27322 6326 27340
rect 6372 27322 6374 27340
rect 6468 27322 6470 27340
rect 6492 27322 6494 27340
rect 6564 27322 6566 27340
rect 6588 27322 6590 27340
rect 6612 27322 6614 27340
rect 6660 27322 6662 27340
rect 6684 27322 6686 27340
rect 6708 27322 6710 27340
rect 6780 27322 6782 27340
rect 6804 27322 6806 27340
rect 6828 27322 6830 27340
rect 6876 27322 6878 27340
rect 6900 27322 6902 27340
rect 6924 27322 6926 27340
rect 6972 27322 6974 27340
rect 7020 27322 7022 27340
rect 7140 27322 7142 27340
rect 7236 27322 7238 27340
rect 7260 27322 7262 27340
rect 7332 27322 7334 27340
rect 7356 27322 7358 27340
rect 7380 27322 7382 27340
rect 7428 27322 7430 27340
rect 7452 27322 7454 27340
rect 7476 27322 7478 27340
rect 7524 27322 7526 27340
rect 7548 27322 7550 27340
rect 7572 27322 7574 27340
rect 7620 27322 7622 27340
rect 7644 27322 7646 27340
rect 7668 27322 7670 27340
rect 7716 27322 7718 27340
rect 7740 27322 7742 27340
rect 7764 27322 7766 27340
rect 7836 27322 7838 27340
rect 7860 27322 7862 27340
rect 7884 27322 7886 27340
rect 7932 27322 7934 27340
rect 7956 27322 7958 27340
rect 7980 27322 7982 27340
rect 8052 27322 8054 27340
rect 8148 27322 8150 27340
rect 8196 27322 8198 27340
rect 8244 27322 8246 27340
rect 8268 27322 8270 27340
rect 8292 27322 8294 27340
rect 8340 27322 8342 27340
rect 8364 27322 8366 27340
rect 8388 27322 8390 27340
rect 8436 27322 8438 27340
rect 8460 27322 8462 27340
rect 8484 27322 8486 27340
rect 8556 27322 8558 27340
rect 8580 27322 8582 27340
rect 8604 27322 8606 27340
rect 8676 27322 8678 27340
rect 8700 27322 8702 27340
rect 8724 27322 8726 27340
rect 8772 27322 8774 27340
rect 8820 27322 8822 27340
rect 8844 27322 8846 27340
rect 8868 27322 8870 27340
rect 9496 27322 9498 27340
rect 9551 27338 9565 27340
rect 9660 27322 9662 27340
rect 9684 27322 9686 27340
rect 9708 27322 9710 27340
rect 9756 27322 9758 27340
rect 9780 27322 9782 27340
rect 9804 27322 9806 27340
rect 9852 27322 9854 27340
rect 9876 27322 9878 27340
rect 9900 27322 9902 27340
rect 9948 27322 9950 27340
rect 9972 27322 9974 27340
rect 9996 27322 9998 27340
rect 10068 27322 10070 27340
rect 10092 27322 10094 27340
rect 10116 27322 10118 27340
rect 10164 27322 10166 27340
rect 10188 27322 10190 27340
rect 10212 27322 10214 27340
rect 10260 27322 10262 27340
rect 10284 27322 10286 27340
rect 10308 27322 10310 27340
rect 10380 27322 10382 27340
rect 10404 27322 10406 27340
rect 10428 27322 10430 27340
rect 10476 27322 10478 27340
rect 10500 27322 10502 27340
rect 10524 27322 10526 27340
rect 10572 27322 10574 27340
rect 10596 27322 10598 27340
rect 10620 27322 10622 27340
rect 10668 27322 10670 27340
rect 10692 27322 10694 27340
rect 10716 27322 10718 27340
rect 10788 27322 10790 27340
rect 10836 27322 10838 27340
rect 10956 27322 10958 27340
rect 11052 27322 11054 27340
rect 11076 27322 11078 27340
rect 11124 27322 11126 27340
rect 11172 27322 11174 27340
rect 11220 27322 11222 27340
rect 11340 27322 11342 27340
rect 11436 27322 11438 27340
rect 11532 27322 11534 27340
rect 11580 27322 11582 27340
rect 11628 27322 11630 27340
rect 11652 27322 11654 27340
rect 11676 27322 11678 27340
rect 11748 27322 11750 27340
rect 11772 27322 11774 27340
rect 11796 27322 11798 27340
rect 11844 27322 11846 27340
rect 11892 27322 11894 27340
rect 11988 27322 11990 27340
rect 12012 27322 12014 27340
rect 12084 27322 12086 27340
rect 12132 27322 12134 27340
rect 12228 27322 12230 27340
rect 12252 27322 12254 27340
rect 12300 27322 12302 27340
rect 12324 27322 12326 27340
rect 12348 27322 12350 27340
rect 12396 27322 12398 27340
rect 12420 27322 12422 27340
rect 12444 27322 12446 27340
rect 12492 27322 12494 27340
rect 12516 27322 12518 27340
rect 12540 27322 12542 27340
rect 12588 27322 12590 27340
rect 12636 27322 12638 27340
rect 12732 27322 12734 27340
rect 12756 27322 12758 27340
rect 12804 27322 12806 27340
rect 12828 27322 12830 27340
rect 12852 27322 12854 27340
rect 12900 27322 12902 27340
rect 12924 27322 12926 27340
rect 12948 27322 12950 27340
rect 13020 27322 13022 27340
rect 13044 27322 13046 27340
rect 13068 27322 13070 27340
rect 13116 27322 13118 27340
rect 13188 27322 13190 27340
rect 13284 27322 13286 27340
rect 13332 27322 13334 27340
rect 13428 27322 13430 27340
rect 13524 27322 13526 27340
rect 13572 27322 13574 27340
rect 13644 27322 13646 27340
rect 13668 27322 13670 27340
rect 13692 27322 13694 27340
rect 13764 27322 13766 27340
rect 13788 27322 13790 27340
rect 13812 27322 13814 27340
rect 13860 27322 13862 27340
rect 13884 27322 13886 27340
rect 13908 27322 13910 27340
rect 13956 27322 13958 27340
rect 14004 27322 14006 27340
rect 14100 27322 14102 27340
rect 14196 27322 14198 27340
rect 14244 27322 14246 27340
rect 14292 27322 14294 27340
rect 14920 27322 14922 27340
rect 14975 27338 14989 27340
rect 15132 27322 15134 27340
rect 15228 27322 15230 27340
rect 15252 27322 15254 27340
rect 15300 27322 15302 27340
rect 15324 27322 15326 27340
rect 15348 27322 15350 27340
rect 15396 27322 15398 27340
rect 15420 27322 15422 27340
rect 15444 27322 15446 27340
rect 15492 27322 15494 27340
rect 15540 27322 15542 27340
rect 15636 27322 15638 27340
rect 15660 27322 15662 27340
rect 15708 27322 15710 27340
rect 15732 27322 15734 27340
rect 15756 27322 15758 27340
rect 15804 27322 15806 27340
rect 15828 27322 15830 27340
rect 15852 27322 15854 27340
rect 15900 27322 15902 27340
rect 15924 27322 15926 27340
rect 15948 27322 15950 27340
rect 15996 27322 15998 27340
rect 16020 27322 16022 27340
rect 16044 27322 16046 27340
rect 16092 27322 16094 27340
rect 16140 27322 16142 27340
rect 16236 27322 16238 27340
rect 16260 27322 16262 27340
rect 16308 27322 16310 27340
rect 16332 27322 16334 27340
rect 16356 27322 16358 27340
rect 16404 27322 16406 27340
rect 16452 27322 16454 27340
rect 16548 27322 16550 27340
rect 16572 27322 16574 27340
rect 16620 27322 16622 27340
rect 16644 27322 16646 27340
rect 16668 27322 16670 27340
rect 16716 27322 16718 27340
rect 16740 27322 16742 27340
rect 16764 27322 16766 27340
rect 16836 27322 16838 27340
rect 16884 27322 16886 27340
rect 16980 27322 16982 27340
rect 17004 27322 17006 27340
rect 17052 27322 17054 27340
rect 17100 27322 17102 27340
rect 17196 27322 17198 27340
rect 17220 27322 17222 27340
rect 17268 27322 17270 27340
rect 17292 27322 17294 27340
rect 17316 27322 17318 27340
rect 17944 27322 17946 27340
rect 17999 27338 18013 27340
rect 18084 27322 18086 27340
rect 18108 27322 18110 27340
rect 18132 27322 18134 27340
rect 18180 27322 18182 27340
rect 18252 27322 18254 27340
rect 18348 27322 18350 27340
rect 18396 27322 18398 27340
rect 18492 27322 18494 27340
rect 18516 27322 18518 27340
rect 18564 27322 18566 27340
rect 18588 27322 18590 27340
rect 18612 27322 18614 27340
rect 18660 27322 18662 27340
rect 18684 27322 18686 27340
rect 18708 27322 18710 27340
rect 18756 27322 18758 27340
rect 18780 27322 18782 27340
rect 18804 27322 18806 27340
rect 18852 27322 18854 27340
rect 18876 27322 18878 27340
rect 18900 27322 18902 27340
rect 18948 27322 18950 27340
rect 18996 27322 18998 27340
rect 19020 27322 19022 27340
rect 19044 27322 19046 27340
rect 19092 27322 19094 27340
rect 19116 27322 19118 27340
rect 19140 27322 19142 27340
rect 19188 27322 19190 27340
rect 19236 27322 19238 27340
rect 19332 27322 19334 27340
rect 19428 27322 19430 27340
rect 19476 27322 19478 27340
rect 19524 27322 19526 27340
rect 19572 27322 19574 27340
rect 19596 27322 19598 27340
rect 19620 27322 19622 27340
rect 19668 27322 19670 27340
rect 19692 27322 19694 27340
rect 19716 27322 19718 27340
rect 19764 27322 19766 27340
rect 19812 27322 19814 27340
rect 19836 27322 19838 27340
rect 19860 27322 19862 27340
rect 19932 27322 19934 27340
rect 19956 27322 19958 27340
rect 19980 27322 19982 27340
rect 20028 27322 20030 27340
rect 20052 27322 20054 27340
rect 20076 27322 20078 27340
rect 20148 27322 20150 27340
rect 20172 27322 20174 27340
rect 20196 27322 20198 27340
rect 20244 27322 20246 27340
rect 20268 27322 20270 27340
rect 20292 27322 20294 27340
rect 20340 27322 20342 27340
rect 20388 27322 20390 27340
rect 20484 27322 20486 27340
rect 20508 27322 20510 27340
rect 20556 27322 20558 27340
rect 20580 27322 20582 27340
rect 20604 27322 20606 27340
rect 20700 27322 20702 27340
rect 20916 27322 20918 27340
rect 20964 27322 20966 27340
rect 21012 27322 21014 27340
rect 21060 27322 21062 27340
rect 21084 27322 21086 27340
rect 21108 27322 21110 27340
rect 21156 27322 21158 27340
rect 21204 27322 21206 27340
rect 21300 27322 21302 27340
rect 21324 27322 21326 27340
rect 21372 27322 21374 27340
rect 21420 27322 21422 27340
rect 21444 27322 21446 27340
rect 21468 27322 21470 27340
rect 21516 27322 21518 27340
rect 21540 27322 21542 27340
rect 21564 27322 21566 27340
rect 21612 27322 21614 27340
rect 21660 27322 21662 27340
rect 21684 27322 21686 27340
rect 21708 27322 21710 27340
rect 21780 27322 21782 27340
rect 21804 27322 21806 27340
rect 21828 27322 21830 27340
rect 21900 27322 21902 27340
rect 21924 27322 21926 27340
rect 21948 27322 21950 27340
rect 22020 27322 22022 27340
rect 22044 27322 22046 27340
rect 22068 27322 22070 27340
rect 22116 27322 22118 27340
rect 22164 27322 22166 27340
rect 22188 27322 22190 27340
rect 22212 27322 22214 27340
rect 22864 27322 22866 27340
rect 22919 27338 22933 27340
rect 23004 27322 23006 27340
rect 23052 27322 23054 27340
rect 23076 27322 23078 27340
rect 23100 27322 23102 27340
rect 23148 27322 23150 27340
rect 23196 27322 23198 27340
rect 23220 27322 23222 27340
rect 23244 27322 23246 27340
rect 23292 27322 23294 27340
rect 23316 27322 23318 27340
rect 23340 27322 23342 27340
rect 23388 27322 23390 27340
rect 23412 27322 23414 27340
rect 23436 27322 23438 27340
rect 23484 27322 23486 27340
rect 23532 27322 23534 27340
rect 23556 27322 23558 27340
rect 23580 27322 23582 27340
rect 23628 27322 23630 27340
rect 23652 27322 23654 27340
rect 23676 27322 23678 27340
rect 23724 27322 23726 27340
rect 23748 27322 23750 27340
rect 23772 27322 23774 27340
rect 23820 27322 23822 27340
rect 23868 27322 23870 27340
rect 23892 27322 23894 27340
rect 23916 27322 23918 27340
rect 23988 27322 23990 27340
rect 24012 27322 24014 27340
rect 24036 27322 24038 27340
rect 24084 27322 24086 27340
rect 24132 27322 24134 27340
rect 24228 27322 24230 27340
rect 24252 27322 24254 27340
rect 24300 27322 24302 27340
rect 24348 27322 24350 27340
rect 24372 27322 24374 27340
rect 24396 27322 24398 27340
rect 24468 27322 24470 27340
rect 24492 27322 24494 27340
rect 24516 27322 24518 27340
rect 24564 27322 24566 27340
rect 24588 27322 24590 27340
rect 24612 27322 24614 27340
rect 24660 27322 24662 27340
rect 24708 27322 24710 27340
rect 24732 27322 24734 27340
rect 24756 27322 24758 27340
rect 24828 27322 24830 27340
rect 24852 27322 24854 27340
rect 24876 27322 24878 27340
rect 24948 27322 24950 27340
rect 24972 27322 24974 27340
rect 24996 27322 24998 27340
rect 25044 27322 25046 27340
rect 25092 27322 25094 27340
rect 25140 27322 25142 27340
rect 25260 27322 25262 27340
rect 25356 27322 25358 27340
rect 25380 27322 25382 27340
rect 25452 27322 25454 27340
rect 25476 27322 25478 27340
rect 25500 27322 25502 27340
rect 25548 27322 25550 27340
rect 25572 27322 25574 27340
rect 25596 27322 25598 27340
rect 25644 27322 25646 27340
rect 26272 27322 26274 27340
rect 26327 27338 26341 27340
rect 26896 27322 26898 27340
rect 26951 27338 26965 27340
rect 27060 27322 27062 27340
rect 27108 27322 27110 27340
rect 27180 27322 27182 27340
rect 27276 27322 27278 27340
rect 27324 27322 27326 27340
rect 27372 27322 27374 27340
rect 27396 27322 27398 27340
rect 27420 27322 27422 27340
rect 27468 27322 27470 27340
rect 27516 27322 27518 27340
rect 27540 27322 27542 27340
rect 27564 27322 27566 27340
rect 28276 27338 28290 27340
rect 28996 27338 29010 27340
rect 29716 27338 29730 27340
rect 30436 27338 30450 27340
rect 30492 27322 30494 27340
rect 30540 27322 30542 27340
rect 30612 27322 30614 27340
rect 30636 27322 30638 27340
rect 30660 27322 30662 27340
rect 30708 27322 30710 27340
rect 30756 27322 30758 27340
rect 30780 27322 30782 27340
rect 30804 27322 30806 27340
rect 30852 27322 30854 27340
rect 30900 27322 30902 27340
rect 30924 27322 30926 27340
rect 30948 27322 30950 27340
rect 30996 27322 30998 27340
rect 31044 27322 31046 27340
rect 31068 27322 31070 27340
rect 31092 27322 31094 27340
rect 31140 27322 31142 27340
rect 31188 27322 31190 27340
rect 31236 27322 31238 27340
rect 31888 27322 31890 27340
rect 31943 27338 31957 27340
rect 32076 27322 32078 27340
rect 32100 27322 32102 27340
rect 32148 27322 32150 27340
rect -19052 27317 32194 27322
rect -17916 27312 -17914 27317
rect -17868 27312 -17866 27317
rect -19038 27304 -19030 27312
rect -19010 27304 -18994 27312
rect -18978 27304 -18966 27312
rect -18950 27304 -18938 27312
rect -18918 27304 -18910 27312
rect -18890 27304 -18874 27312
rect -18858 27304 -18846 27312
rect -18830 27304 -18818 27312
rect -18798 27304 -18790 27312
rect -18770 27304 -18754 27312
rect -18738 27304 -18726 27312
rect -18710 27304 -18698 27312
rect -18678 27304 -18670 27312
rect -18650 27304 -18634 27312
rect -18618 27304 -18606 27312
rect -18590 27304 -18578 27312
rect -18558 27304 -18550 27312
rect -18530 27304 -18514 27312
rect -18498 27304 -18486 27312
rect -18470 27304 -18458 27312
rect -18438 27304 -18430 27312
rect -18410 27304 -18394 27312
rect -18378 27304 -18366 27312
rect -18350 27304 -18338 27312
rect -18318 27304 -18310 27312
rect -18290 27304 -18274 27312
rect -18258 27304 -18246 27312
rect -18230 27304 -18218 27312
rect -18198 27304 -18190 27312
rect -18170 27304 -18154 27312
rect -18138 27304 -18126 27312
rect -18110 27304 -18098 27312
rect -18078 27304 -18070 27312
rect -18050 27304 -18034 27312
rect -18018 27304 -18006 27312
rect -17990 27304 -17978 27312
rect -17958 27304 -17950 27312
rect -17930 27304 -17914 27312
rect -17900 27304 -17888 27312
rect -17872 27304 -17860 27312
rect -19030 27296 -19022 27304
rect -18982 27296 -18978 27304
rect -18954 27296 -18950 27304
rect -18910 27296 -18902 27304
rect -18862 27296 -18858 27304
rect -18834 27296 -18830 27304
rect -18790 27296 -18782 27304
rect -18742 27296 -18738 27304
rect -18714 27296 -18710 27304
rect -18670 27296 -18662 27304
rect -18622 27296 -18618 27304
rect -18594 27296 -18590 27304
rect -18550 27296 -18542 27304
rect -18502 27296 -18498 27304
rect -18474 27296 -18470 27304
rect -18430 27296 -18422 27304
rect -18382 27296 -18378 27304
rect -18354 27296 -18350 27304
rect -18310 27296 -18302 27304
rect -18262 27296 -18258 27304
rect -18234 27296 -18230 27304
rect -18190 27296 -18182 27304
rect -18142 27296 -18138 27304
rect -18114 27296 -18110 27304
rect -18070 27296 -18062 27304
rect -18022 27296 -18018 27304
rect -17994 27296 -17990 27304
rect -17950 27296 -17942 27304
rect -19052 27294 -19041 27296
rect -19052 27279 -19043 27287
rect -18980 27078 -18977 27090
rect -19028 27071 -19011 27078
rect -18968 27071 -18965 27078
rect -18968 27028 -18964 27068
rect -18952 27058 -18947 27064
rect -18963 27048 -18952 27058
rect -18950 27028 -18947 27058
rect -18941 27048 -18937 27111
rect -18860 27083 -18849 27090
rect -18740 27083 -18729 27090
rect -18620 27083 -18609 27090
rect -18500 27083 -18489 27090
rect -18380 27083 -18369 27090
rect -18260 27083 -18249 27090
rect -18140 27083 -18129 27090
rect -18020 27083 -18009 27090
rect -18858 27078 -18849 27083
rect -18738 27078 -18729 27083
rect -18618 27078 -18609 27083
rect -18498 27078 -18489 27083
rect -18378 27078 -18369 27083
rect -18258 27078 -18249 27083
rect -18138 27078 -18129 27083
rect -18018 27078 -18009 27083
rect -18848 27048 -18837 27078
rect -18728 27048 -18717 27078
rect -18608 27048 -18597 27078
rect -18488 27048 -18477 27078
rect -18368 27048 -18357 27078
rect -18248 27048 -18237 27078
rect -18128 27048 -18117 27078
rect -18008 27048 -17997 27078
rect -17916 27059 -17914 27304
rect -17902 27296 -17900 27304
rect -17888 27296 -17886 27304
rect -17874 27296 -17872 27304
rect -17905 27083 -17889 27091
rect -17923 27049 -17914 27059
rect -17912 27049 -17906 27079
rect -17905 27077 -17894 27079
rect -17905 27049 -17896 27070
rect -18848 27040 -18839 27048
rect -18728 27040 -18719 27048
rect -18608 27040 -18599 27048
rect -18488 27040 -18479 27048
rect -18368 27040 -18359 27048
rect -18248 27040 -18239 27048
rect -18128 27040 -18119 27048
rect -18008 27040 -17999 27048
rect -17916 27015 -17914 27049
rect -17913 27040 -17906 27049
rect -17894 27040 -17889 27070
rect -17913 27015 -17912 27040
rect -17880 27039 -17876 27049
rect -17868 27039 -17866 27304
rect -17860 27296 -17858 27304
rect -17846 27079 -17842 27081
rect -17848 27071 -17842 27079
rect -17847 27049 -17842 27051
rect -17836 27049 -17830 27071
rect -17820 27056 -17818 27317
rect -17772 27312 -17770 27317
rect -17652 27312 -17650 27317
rect -17532 27312 -17530 27317
rect -17436 27312 -17434 27317
rect -17412 27312 -17410 27317
rect -17806 27304 -17796 27312
rect -17778 27304 -17768 27312
rect -17746 27304 -17738 27312
rect -17682 27304 -17674 27312
rect -17654 27304 -17646 27312
rect -17622 27304 -17614 27312
rect -17594 27304 -17578 27312
rect -17562 27304 -17550 27312
rect -17534 27304 -17522 27312
rect -17502 27304 -17494 27312
rect -17474 27304 -17460 27312
rect -17444 27304 -17432 27312
rect -17416 27304 -17404 27312
rect -17812 27296 -17806 27304
rect -17784 27296 -17778 27304
rect -17815 27083 -17806 27084
rect -17796 27083 -17789 27084
rect -17782 27083 -17781 27279
rect -17772 27083 -17770 27304
rect -17738 27296 -17730 27304
rect -17690 27296 -17682 27304
rect -17662 27296 -17654 27304
rect -17672 27116 -17658 27132
rect -17815 27082 -17784 27083
rect -17782 27082 -17754 27083
rect -17739 27082 -17729 27104
rect -17822 27046 -17818 27056
rect -18848 27013 -18846 27015
rect -18728 27013 -18726 27015
rect -18608 27013 -18606 27015
rect -18488 27013 -18486 27015
rect -18368 27013 -18366 27015
rect -18248 27013 -18246 27015
rect -18128 27013 -18126 27015
rect -18008 27013 -18006 27015
rect -19016 26998 -19014 27010
rect -18856 27004 -18846 27013
rect -18736 27004 -18726 27013
rect -18616 27004 -18606 27013
rect -18496 27004 -18486 27013
rect -18376 27004 -18366 27013
rect -18256 27004 -18246 27013
rect -18136 27004 -18126 27013
rect -18016 27004 -18006 27013
rect -18972 26999 -18968 27002
rect -19024 26992 -19014 26998
rect -18948 26997 -18938 27002
rect -18852 26999 -18842 27004
rect -18732 26999 -18722 27004
rect -18612 26999 -18602 27004
rect -18492 26999 -18482 27004
rect -18372 26999 -18362 27004
rect -18252 26999 -18242 27004
rect -18132 26999 -18122 27004
rect -18012 26999 -18002 27004
rect -19028 26987 -19024 26992
rect -17916 26991 -17912 27015
rect -17906 27004 -17904 27014
rect -17894 27004 -17887 27015
rect -17870 27009 -17866 27039
rect -18848 26989 -18846 26990
rect -18728 26989 -18726 26990
rect -18608 26989 -18606 26990
rect -18488 26989 -18486 26990
rect -18368 26989 -18366 26990
rect -18248 26989 -18246 26990
rect -18128 26989 -18126 26990
rect -18008 26989 -18006 26990
rect -17916 26987 -17914 26991
rect -17913 26987 -17912 26991
rect -17896 26991 -17887 27004
rect -17882 26991 -17878 27004
rect -17896 26990 -17882 26991
rect -17894 26989 -17886 26990
rect -17868 26987 -17866 27009
rect -17820 26987 -17818 27046
rect -17812 27041 -17810 27046
rect -17792 27041 -17788 27056
rect -17784 27041 -17782 27071
rect -17772 27041 -17770 27082
rect -17767 27041 -17766 27071
rect -17806 27036 -17770 27041
rect -17736 27038 -17722 27046
rect -17806 27032 -17798 27036
rect -17792 27032 -17788 27036
rect -17806 27031 -17802 27032
rect -17796 27015 -17792 27031
rect -17794 27012 -17792 27015
rect -17786 27012 -17780 27020
rect -17794 27001 -17780 27012
rect -17772 27010 -17770 27036
rect -17686 27027 -17681 27057
rect -17672 27029 -17660 27038
rect -17652 27034 -17650 27304
rect -17614 27296 -17606 27304
rect -17566 27296 -17562 27304
rect -17538 27296 -17534 27304
rect -17589 27057 -17580 27067
rect -17674 27027 -17655 27029
rect -17776 26996 -17770 27010
rect -17699 27002 -17690 27014
rect -17654 27008 -17650 27034
rect -17623 27019 -17620 27049
rect -17618 27027 -17607 27049
rect -17605 27027 -17602 27057
rect -17596 27019 -17592 27027
rect -17579 27019 -17570 27057
rect -17551 27027 -17544 27057
rect -17532 27049 -17530 27304
rect -17494 27296 -17486 27304
rect -17460 27296 -17458 27304
rect -17446 27296 -17444 27304
rect -17466 27079 -17460 27089
rect -17542 27027 -17536 27049
rect -17561 27019 -17554 27027
rect -17534 27019 -17527 27049
rect -17503 27019 -17500 27049
rect -17498 27027 -17487 27049
rect -17485 27027 -17482 27057
rect -17467 27049 -17460 27059
rect -17456 27049 -17450 27079
rect -17436 27049 -17434 27304
rect -17432 27296 -17430 27304
rect -17418 27296 -17416 27304
rect -17431 27049 -17424 27057
rect -17412 27049 -17410 27304
rect -17404 27296 -17402 27304
rect -17390 27079 -17386 27081
rect -17392 27071 -17386 27079
rect -17402 27049 -17396 27059
rect -17391 27049 -17386 27051
rect -17380 27049 -17374 27071
rect -17364 27056 -17362 27317
rect -17316 27312 -17314 27317
rect -17220 27312 -17218 27317
rect -17196 27312 -17194 27317
rect -17124 27312 -17122 27317
rect -17028 27312 -17026 27317
rect -16980 27312 -16978 27317
rect -16884 27312 -16882 27317
rect -16860 27312 -16858 27317
rect -17350 27304 -17340 27312
rect -17322 27304 -17312 27312
rect -17290 27304 -17282 27312
rect -17228 27304 -17218 27312
rect -17200 27304 -17190 27312
rect -17130 27304 -17122 27312
rect -17102 27304 -17096 27312
rect -17070 27304 -17062 27312
rect -17042 27304 -17026 27312
rect -17010 27304 -16998 27312
rect -16982 27304 -16970 27312
rect -16950 27304 -16942 27312
rect -16922 27304 -16908 27312
rect -16892 27304 -16880 27312
rect -16864 27304 -16852 27312
rect -17356 27296 -17350 27304
rect -17328 27296 -17322 27304
rect -17359 27083 -17350 27084
rect -17340 27083 -17333 27084
rect -17326 27083 -17325 27279
rect -17316 27083 -17314 27304
rect -17282 27296 -17274 27304
rect -17234 27296 -17228 27304
rect -17359 27082 -17328 27083
rect -17326 27082 -17298 27083
rect -17283 27082 -17273 27104
rect -17476 27019 -17472 27027
rect -17457 27019 -17450 27049
rect -17438 27019 -17431 27049
rect -17424 27039 -17420 27049
rect -17412 27039 -17406 27049
rect -17366 27046 -17362 27056
rect -17416 27023 -17406 27039
rect -17414 27019 -17406 27023
rect -17772 26987 -17770 26996
rect -17652 26987 -17650 27008
rect -17612 26987 -17603 27019
rect -17551 26987 -17544 27019
rect -17532 26987 -17530 27019
rect -17492 26987 -17483 27019
rect -17436 26987 -17434 27019
rect -17414 27009 -17410 27019
rect -17412 27001 -17410 27009
rect -17416 26987 -17410 27001
rect -17364 26987 -17362 27046
rect -17356 27041 -17354 27046
rect -17336 27041 -17332 27056
rect -17328 27041 -17326 27071
rect -17316 27041 -17314 27082
rect -17232 27079 -17224 27090
rect -17220 27087 -17218 27304
rect -17206 27296 -17200 27304
rect -17240 27074 -17232 27079
rect -17230 27074 -17224 27079
rect -17222 27074 -17215 27087
rect -17200 27079 -17197 27092
rect -17311 27041 -17310 27071
rect -17230 27049 -17223 27074
rect -17220 27049 -17218 27074
rect -17350 27036 -17314 27041
rect -17280 27038 -17266 27046
rect -17350 27032 -17342 27036
rect -17336 27032 -17332 27036
rect -17350 27031 -17346 27032
rect -17340 27015 -17336 27031
rect -17338 27012 -17336 27015
rect -17330 27012 -17324 27020
rect -17338 27001 -17324 27012
rect -17316 27010 -17314 27036
rect -17222 27024 -17215 27049
rect -17208 27039 -17204 27049
rect -17196 27039 -17194 27304
rect -17140 27296 -17130 27304
rect -17174 27079 -17170 27081
rect -17176 27071 -17170 27079
rect -17175 27049 -17170 27051
rect -17164 27049 -17158 27071
rect -17320 26996 -17314 27010
rect -17241 27002 -17234 27014
rect -17220 27008 -17218 27024
rect -17200 27023 -17194 27039
rect -17198 27009 -17194 27023
rect -17316 26987 -17314 26996
rect -17222 26987 -17215 27008
rect -17196 26987 -17194 27009
rect -17124 27013 -17122 27304
rect -17112 27296 -17102 27304
rect -17062 27296 -17054 27304
rect -17119 27048 -17112 27078
rect -17110 27048 -17104 27071
rect -17102 27041 -17095 27071
rect -17093 27048 -17084 27279
rect -17028 27067 -17026 27304
rect -17014 27296 -17010 27304
rect -16986 27296 -16982 27304
rect -17037 27057 -17026 27067
rect -17110 27013 -17108 27023
rect -17102 27015 -17098 27041
rect -17028 27040 -17018 27057
rect -17017 27040 -17011 27057
rect -17009 27040 -17002 27065
rect -17000 27040 -16991 27279
rect -17028 27027 -17019 27040
rect -17124 27001 -17110 27013
rect -17100 27001 -17098 27013
rect -17124 26993 -17122 27001
rect -17124 26987 -17120 26993
rect -17028 26987 -17024 27027
rect -17018 27004 -17016 27014
rect -17008 26990 -17006 27004
rect -16980 26987 -16978 27304
rect -16942 27296 -16934 27304
rect -16908 27296 -16906 27304
rect -16894 27296 -16892 27304
rect -16914 27079 -16908 27089
rect -16951 27019 -16948 27049
rect -16946 27027 -16935 27049
rect -16933 27027 -16930 27057
rect -16915 27049 -16908 27059
rect -16904 27049 -16898 27079
rect -16884 27049 -16882 27304
rect -16880 27296 -16878 27304
rect -16866 27296 -16864 27304
rect -16879 27049 -16872 27057
rect -16860 27049 -16858 27304
rect -16852 27296 -16850 27304
rect -16838 27079 -16834 27081
rect -16840 27071 -16834 27079
rect -16850 27049 -16844 27059
rect -16839 27049 -16834 27051
rect -16828 27049 -16822 27071
rect -16812 27059 -16810 27317
rect -16788 27312 -16786 27317
rect -16764 27312 -16762 27317
rect -16796 27304 -16786 27312
rect -16768 27304 -16760 27312
rect -16804 27296 -16796 27304
rect -16819 27049 -16810 27059
rect -16808 27049 -16802 27079
rect -16788 27049 -16786 27304
rect -16776 27296 -16768 27304
rect -16783 27071 -16776 27079
rect -16764 27071 -16762 27304
rect -16754 27149 -16748 27279
rect -16754 27133 -16746 27149
rect -16764 27049 -16758 27071
rect -16754 27049 -16748 27133
rect -16742 27079 -16738 27081
rect -16744 27071 -16738 27079
rect -16743 27049 -16738 27051
rect -16732 27049 -16726 27071
rect -16716 27059 -16714 27317
rect -16692 27312 -16690 27317
rect -16668 27312 -16666 27317
rect -16700 27304 -16690 27312
rect -16672 27304 -16664 27312
rect -16612 27304 -16607 27312
rect -16596 27304 -16594 27317
rect -16500 27312 -16498 27317
rect -16404 27312 -16402 27317
rect -16380 27312 -16378 27317
rect -16584 27304 -16579 27312
rect -16531 27304 -16523 27312
rect -16503 27304 -16495 27312
rect -16475 27304 -16467 27312
rect -16412 27304 -16402 27312
rect -16384 27304 -16375 27312
rect -16708 27296 -16700 27304
rect -16723 27049 -16714 27059
rect -16712 27049 -16706 27079
rect -16692 27049 -16690 27304
rect -16680 27296 -16672 27304
rect -16687 27071 -16680 27079
rect -16668 27071 -16666 27304
rect -16607 27296 -16594 27304
rect -16579 27296 -16568 27304
rect -16523 27296 -16515 27304
rect -16634 27294 -16594 27296
rect -16634 27288 -16624 27294
rect -16612 27288 -16594 27294
rect -16658 27149 -16652 27279
rect -16658 27133 -16650 27149
rect -16668 27049 -16662 27071
rect -16658 27049 -16652 27133
rect -16646 27079 -16642 27081
rect -16648 27071 -16642 27079
rect -16647 27049 -16642 27051
rect -16636 27049 -16630 27071
rect -16622 27053 -16620 27071
rect -16618 27053 -16611 27079
rect -16924 27019 -16920 27027
rect -16905 27019 -16898 27049
rect -16886 27019 -16879 27049
rect -16872 27039 -16868 27049
rect -16860 27039 -16854 27049
rect -16864 27023 -16854 27039
rect -16862 27019 -16854 27023
rect -16940 26987 -16931 27019
rect -16884 26987 -16882 27019
rect -16862 27009 -16858 27019
rect -16860 27001 -16858 27009
rect -16864 26987 -16858 27001
rect -16812 26987 -16810 27049
rect -16809 27041 -16802 27049
rect -16790 27041 -16783 27049
rect -16778 27041 -16758 27049
rect -16809 27023 -16808 27041
rect -16788 26993 -16786 27041
rect -16778 27039 -16772 27041
rect -16764 27039 -16762 27041
rect -16768 27023 -16762 27039
rect -16766 27009 -16762 27023
rect -16788 26987 -16784 26993
rect -16764 26987 -16762 27009
rect -16716 26987 -16714 27049
rect -16713 27041 -16706 27049
rect -16694 27041 -16687 27049
rect -16682 27041 -16662 27049
rect -16713 27023 -16712 27041
rect -16692 26993 -16690 27041
rect -16682 27039 -16676 27041
rect -16668 27039 -16666 27041
rect -16672 27023 -16666 27039
rect -16670 27009 -16666 27023
rect -16604 27031 -16597 27053
rect -16596 27031 -16594 27288
rect -16577 27126 -16574 27128
rect -16582 27125 -16574 27126
rect -16570 27125 -16566 27137
rect -16540 27131 -16533 27133
rect -16540 27125 -16530 27131
rect -16546 27120 -16530 27125
rect -16558 27095 -16556 27101
rect -16527 27100 -16520 27279
rect -16517 27100 -16501 27117
rect -16528 27095 -16501 27100
rect -16575 27083 -16566 27093
rect -16528 27083 -16520 27095
rect -16508 27083 -16502 27093
rect -16500 27085 -16498 27304
rect -16495 27296 -16487 27304
rect -16467 27296 -16459 27304
rect -16419 27296 -16412 27304
rect -16482 27087 -16475 27117
rect -16472 27095 -16466 27117
rect -16464 27095 -16457 27125
rect -16591 27053 -16584 27079
rect -16565 27075 -16549 27083
rect -16528 27075 -16523 27083
rect -16500 27075 -16490 27085
rect -16482 27075 -16481 27087
rect -16451 27075 -16446 27279
rect -16404 27091 -16402 27304
rect -16391 27296 -16384 27304
rect -16380 27092 -16378 27304
rect -16384 27091 -16378 27092
rect -16436 27087 -16378 27091
rect -16582 27053 -16578 27071
rect -16574 27053 -16567 27071
rect -16565 27053 -16556 27075
rect -16546 27053 -16533 27075
rect -16582 27041 -16567 27053
rect -16546 27045 -16530 27053
rect -16527 27052 -16518 27061
rect -16527 27045 -16520 27052
rect -16518 27045 -16511 27052
rect -16509 27045 -16502 27075
rect -16500 27045 -16492 27075
rect -16489 27045 -16475 27075
rect -16424 27056 -16421 27079
rect -16404 27056 -16402 27087
rect -16380 27056 -16378 27087
rect -16358 27079 -16354 27081
rect -16360 27071 -16354 27079
rect -16472 27052 -16463 27056
rect -16461 27052 -16456 27054
rect -16472 27045 -16456 27052
rect -16424 27049 -16368 27056
rect -16359 27049 -16354 27051
rect -16348 27049 -16342 27071
rect -16332 27059 -16330 27317
rect -16308 27312 -16306 27317
rect -16284 27312 -16282 27317
rect -16316 27304 -16306 27312
rect -16288 27304 -16280 27312
rect -16324 27296 -16316 27304
rect -16339 27049 -16330 27059
rect -16328 27049 -16322 27079
rect -16308 27049 -16306 27304
rect -16296 27296 -16288 27304
rect -16303 27071 -16296 27079
rect -16284 27071 -16282 27304
rect -16274 27149 -16268 27279
rect -16274 27133 -16266 27149
rect -16284 27049 -16278 27071
rect -16274 27049 -16268 27133
rect -16262 27079 -16258 27081
rect -16264 27071 -16258 27079
rect -16263 27049 -16258 27051
rect -16252 27049 -16246 27071
rect -16236 27059 -16234 27317
rect -16212 27312 -16210 27317
rect -16188 27312 -16186 27317
rect -15723 27314 -15707 27317
rect -16220 27304 -16210 27312
rect -16192 27304 -16184 27312
rect -16125 27304 -16116 27312
rect -16096 27304 -16088 27312
rect -16065 27304 -16055 27312
rect -16036 27304 -16027 27312
rect -16007 27304 -15999 27312
rect -15979 27304 -15971 27312
rect -15951 27304 -15942 27312
rect -15923 27304 -15914 27312
rect -15894 27304 -15886 27312
rect -15866 27304 -15858 27312
rect -15838 27304 -15830 27312
rect -15810 27304 -15802 27312
rect -15782 27304 -15774 27312
rect -15754 27304 -15746 27312
rect -15560 27309 -15558 27317
rect -15698 27304 -15690 27309
rect -15670 27304 -15662 27309
rect -16228 27296 -16220 27304
rect -16243 27049 -16234 27059
rect -16232 27049 -16226 27079
rect -16212 27049 -16210 27304
rect -16200 27296 -16192 27304
rect -16207 27071 -16200 27079
rect -16188 27071 -16186 27304
rect -16132 27296 -16125 27304
rect -16104 27296 -16096 27304
rect -16055 27296 -16049 27304
rect -16027 27296 -16020 27304
rect -15999 27296 -15991 27304
rect -15971 27296 -15963 27304
rect -15942 27296 -15935 27304
rect -15914 27296 -15907 27304
rect -15886 27296 -15878 27304
rect -15858 27296 -15850 27304
rect -15830 27296 -15822 27304
rect -15802 27296 -15794 27304
rect -15774 27296 -15766 27304
rect -15746 27296 -15738 27304
rect -15690 27293 -15682 27304
rect -15662 27294 -15654 27304
rect -15614 27301 -15606 27309
rect -15586 27301 -15578 27309
rect -15560 27301 -15550 27309
rect -15530 27301 -15516 27312
rect -15500 27301 -15488 27312
rect -15472 27301 -15460 27312
rect -15606 27294 -15598 27301
rect -15578 27294 -15570 27301
rect -15670 27293 -15654 27294
rect -15614 27293 -15598 27294
rect -15586 27293 -15570 27294
rect -15560 27294 -15558 27301
rect -15550 27294 -15542 27301
rect -15516 27296 -15514 27301
rect -15502 27296 -15500 27301
rect -15488 27296 -15486 27301
rect -15474 27296 -15472 27301
rect -15460 27296 -15458 27301
rect -15560 27293 -15542 27294
rect -15530 27293 -15522 27294
rect -16010 27279 -15877 27287
rect -15872 27279 -15819 27287
rect -16178 27149 -16172 27279
rect -15862 27261 -15858 27270
rect -15794 27269 -15787 27278
rect -15811 27257 -15805 27262
rect -15786 27257 -15777 27269
rect -15815 27252 -15811 27257
rect -15786 27253 -15770 27257
rect -15769 27253 -15766 27257
rect -16178 27133 -16170 27149
rect -16188 27049 -16182 27071
rect -16178 27049 -16172 27133
rect -16166 27079 -16162 27081
rect -16102 27080 -16096 27248
rect -16037 27238 -16031 27246
rect -16000 27238 -15989 27242
rect -16027 27230 -16021 27238
rect -16046 27210 -16031 27230
rect -16000 27227 -15987 27238
rect -15962 27230 -15955 27238
rect -15971 27227 -15955 27230
rect -15924 27227 -15914 27249
rect -16046 27200 -16027 27210
rect -16020 27200 -16001 27210
rect -16027 27198 -16021 27200
rect -15980 27198 -15977 27227
rect -15971 27208 -15963 27227
rect -15897 27219 -15891 27249
rect -15856 27219 -15851 27249
rect -15815 27227 -15814 27252
rect -15782 27227 -15775 27253
rect -15975 27200 -15962 27208
rect -16027 27192 -16020 27198
rect -16027 27190 -16013 27192
rect -16027 27185 -16004 27190
rect -16038 27160 -16031 27170
rect -16020 27168 -16004 27185
rect -15994 27168 -15987 27198
rect -15973 27195 -15955 27198
rect -15980 27166 -15973 27190
rect -15965 27168 -15955 27195
rect -15782 27193 -15777 27227
rect -15745 27221 -15736 27222
rect -15739 27219 -15736 27221
rect -15904 27190 -15898 27193
rect -16020 27160 -15966 27166
rect -15965 27160 -15956 27168
rect -15939 27163 -15923 27190
rect -15904 27163 -15901 27190
rect -15898 27163 -15897 27190
rect -15863 27185 -15858 27193
rect -15863 27163 -15847 27185
rect -15841 27163 -15833 27185
rect -15939 27160 -15932 27163
rect -15897 27160 -15891 27163
rect -16030 27153 -16021 27160
rect -15863 27155 -15825 27163
rect -15794 27155 -15787 27185
rect -15782 27163 -15775 27193
rect -15560 27186 -15558 27293
rect -15773 27163 -15766 27185
rect -15761 27163 -15757 27185
rect -15773 27155 -15756 27163
rect -15672 27156 -15660 27172
rect -16092 27125 -16086 27130
rect -16168 27071 -16162 27079
rect -16167 27049 -16162 27051
rect -16156 27049 -16150 27071
rect -16591 27031 -16587 27041
rect -16604 27020 -16601 27031
rect -16607 27010 -16601 27020
rect -16596 27015 -16587 27031
rect -16574 27015 -16570 27041
rect -16528 27022 -16521 27045
rect -16500 27022 -16491 27045
rect -16464 27044 -16456 27045
rect -16404 27044 -16402 27049
rect -16464 27035 -16457 27044
rect -16473 27022 -16457 27035
rect -16451 27022 -16444 27044
rect -16406 27041 -16399 27044
rect -16596 27010 -16594 27015
rect -16591 27010 -16587 27015
rect -16692 26987 -16688 26993
rect -16668 26987 -16666 27009
rect -16604 26987 -16601 27010
rect -16597 27001 -16581 27010
rect -16597 26994 -16594 27001
rect -16596 26993 -16594 26994
rect -16596 26987 -16592 26993
rect -16591 26987 -16587 27001
rect -16528 26987 -16523 27022
rect -16500 26987 -16492 27022
rect -16482 26987 -16481 27022
rect -16473 27017 -16465 27022
rect -16473 27014 -16452 27017
rect -16404 26991 -16402 27041
rect -16392 27039 -16388 27049
rect -16380 27044 -16378 27049
rect -16384 27014 -16378 27044
rect -16382 27009 -16378 27014
rect -16464 26987 -16463 26991
rect -16404 26987 -16390 26991
rect -16380 26987 -16376 27009
rect -16332 26987 -16330 27049
rect -16329 27041 -16322 27049
rect -16310 27041 -16303 27049
rect -16298 27041 -16278 27049
rect -16329 27023 -16328 27041
rect -16308 26993 -16306 27041
rect -16298 27039 -16292 27041
rect -16284 27039 -16282 27041
rect -16288 27023 -16282 27039
rect -16286 27009 -16282 27023
rect -16308 26987 -16304 26993
rect -16284 26987 -16282 27009
rect -16236 26987 -16234 27049
rect -16233 27041 -16226 27049
rect -16214 27041 -16207 27049
rect -16202 27041 -16182 27049
rect -16104 27041 -16099 27071
rect -16030 27070 -16023 27153
rect -15980 27122 -15977 27133
rect -15898 27132 -15891 27148
rect -15889 27133 -15859 27140
rect -15782 27130 -15777 27155
rect -15581 27148 -15580 27164
rect -15565 27162 -15557 27186
rect -15766 27133 -15752 27140
rect -15980 27092 -15973 27122
rect -15863 27100 -15858 27130
rect -15822 27100 -15815 27130
rect -15794 27100 -15793 27122
rect -15782 27100 -15775 27130
rect -15809 27092 -15787 27100
rect -15761 27092 -15754 27122
rect -15703 27106 -15690 27122
rect -15685 27106 -15681 27136
rect -15603 27110 -15587 27126
rect -15594 27101 -15587 27110
rect -15582 27106 -15580 27128
rect -15565 27106 -15556 27146
rect -15458 27140 -15453 27279
rect -15458 27133 -15451 27140
rect -15611 27098 -15607 27101
rect -15596 27098 -15580 27101
rect -15458 27098 -15453 27133
rect -15980 27070 -15977 27092
rect -15782 27083 -15777 27092
rect -16046 27062 -15994 27070
rect -15987 27062 -15975 27070
rect -15931 27062 -15895 27070
rect -16233 27023 -16232 27041
rect -16212 26993 -16210 27041
rect -16202 27039 -16196 27041
rect -16188 27039 -16186 27041
rect -16192 27023 -16186 27039
rect -16190 27009 -16186 27023
rect -16212 26987 -16208 26993
rect -16188 26987 -16186 27009
rect -16030 26987 -16023 27062
rect -15980 27060 -15977 27062
rect -15994 27052 -15987 27060
rect -15994 27030 -15978 27052
rect -15962 27030 -15955 27060
rect -15904 27052 -15898 27060
rect -15863 27052 -15858 27060
rect -15782 27057 -15775 27083
rect -15782 27052 -15777 27057
rect -15921 27030 -15909 27052
rect -15904 27030 -15903 27052
rect -15898 27030 -15897 27052
rect -15858 27030 -15856 27052
rect -15845 27030 -15830 27052
rect -15897 27027 -15891 27030
rect -15925 27022 -15891 27027
rect -15856 27022 -15851 27030
rect -15794 27022 -15787 27052
rect -15761 27026 -15754 27052
rect -15752 27047 -15744 27082
rect -15673 27027 -15669 27043
rect -15668 27041 -15657 27043
rect -15621 27041 -15615 27098
rect -15602 27071 -15601 27073
rect -15594 27071 -15588 27098
rect -15545 27083 -15542 27091
rect -15535 27081 -15532 27083
rect -15605 27041 -15598 27071
rect -15592 27041 -15587 27063
rect -15582 27041 -15576 27063
rect -15574 27041 -15567 27071
rect -15565 27041 -15556 27081
rect -15555 27041 -15549 27063
rect -15547 27041 -15540 27071
rect -15535 27041 -15529 27081
rect -15512 27049 -15511 27079
rect -15496 27063 -15490 27065
rect -15487 27063 -15481 27079
rect -15458 27073 -15456 27093
rect -15446 27079 -15442 27081
rect -15506 27049 -15496 27063
rect -15494 27049 -15490 27063
rect -15488 27049 -15487 27063
rect -15658 27035 -15657 27041
rect -15594 27033 -15587 27041
rect -15565 27033 -15557 27041
rect -15494 27033 -15488 27049
rect -15467 27043 -15463 27063
rect -15458 27049 -15453 27073
rect -15448 27071 -15442 27079
rect -15447 27049 -15442 27051
rect -15436 27049 -15430 27071
rect -15420 27059 -15418 27317
rect -15396 27312 -15394 27317
rect -15372 27312 -15370 27317
rect -15300 27312 -15298 27317
rect -15404 27304 -15394 27312
rect -15376 27304 -15368 27312
rect -15306 27304 -15298 27312
rect -15278 27304 -15272 27312
rect -15246 27304 -15238 27312
rect -15218 27304 -15202 27312
rect -15186 27304 -15174 27312
rect -15158 27304 -15146 27312
rect -15126 27304 -15118 27312
rect -15098 27304 -15086 27312
rect -15084 27304 -15082 27317
rect -15036 27312 -15034 27317
rect -14940 27312 -14938 27317
rect -14916 27312 -14914 27317
rect -15070 27304 -15058 27312
rect -15042 27304 -15030 27312
rect -15010 27304 -15002 27312
rect -14948 27304 -14938 27312
rect -14920 27304 -14910 27312
rect -15412 27296 -15404 27304
rect -15427 27049 -15418 27059
rect -15416 27049 -15410 27079
rect -15396 27049 -15394 27304
rect -15384 27296 -15376 27304
rect -15391 27071 -15384 27079
rect -15372 27071 -15370 27304
rect -15316 27296 -15306 27304
rect -15362 27149 -15356 27279
rect -15362 27133 -15354 27149
rect -15372 27049 -15366 27071
rect -15362 27049 -15356 27133
rect -15350 27079 -15346 27081
rect -15352 27071 -15346 27079
rect -15351 27049 -15346 27051
rect -15340 27049 -15334 27071
rect -15467 27039 -15462 27043
rect -15472 27033 -15463 27039
rect -15770 27022 -15754 27026
rect -15980 26987 -15977 27022
rect -15909 26999 -15905 27015
rect -15904 26987 -15901 26995
rect -15845 26991 -15829 26993
rect -15782 26987 -15777 27022
rect -15594 27018 -15588 27033
rect -15695 27008 -15687 27018
rect -15594 27013 -15579 27018
rect -15685 27008 -15676 27011
rect -15685 26992 -15677 27008
rect -15676 26995 -15669 27008
rect -15594 27003 -15588 27013
rect -15564 26987 -15557 27033
rect -15472 27023 -15471 27033
rect -15502 26991 -15493 27001
rect -15492 26990 -15483 26991
rect -15420 26987 -15418 27049
rect -15417 27041 -15410 27049
rect -15398 27041 -15391 27049
rect -15386 27041 -15366 27049
rect -15417 27023 -15416 27041
rect -15396 26993 -15394 27041
rect -15386 27039 -15380 27041
rect -15372 27039 -15370 27041
rect -15376 27023 -15370 27039
rect -15374 27009 -15370 27023
rect -15396 26987 -15392 26993
rect -15372 26987 -15370 27009
rect -15300 27013 -15298 27304
rect -15288 27296 -15278 27304
rect -15238 27296 -15230 27304
rect -15190 27296 -15186 27304
rect -15162 27296 -15158 27304
rect -15118 27296 -15110 27304
rect -15086 27296 -15082 27304
rect -15058 27296 -15054 27304
rect -15295 27048 -15288 27078
rect -15286 27048 -15280 27071
rect -15278 27041 -15271 27071
rect -15269 27048 -15260 27279
rect -15188 27083 -15177 27090
rect -15186 27078 -15177 27083
rect -15176 27048 -15165 27078
rect -15084 27056 -15082 27296
rect -15073 27083 -15057 27099
rect -15079 27082 -15070 27083
rect -15286 27013 -15284 27023
rect -15278 27015 -15274 27041
rect -15176 27040 -15167 27048
rect -15086 27046 -15082 27056
rect -15084 27015 -15082 27046
rect -15076 27040 -15074 27046
rect -15073 27040 -15062 27046
rect -15058 27040 -15057 27070
rect -15056 27032 -15052 27040
rect -15176 27013 -15174 27015
rect -15300 27001 -15286 27013
rect -15276 27001 -15274 27013
rect -15184 27004 -15174 27013
rect -15300 26993 -15298 27001
rect -15180 26999 -15170 27004
rect -15300 26987 -15296 26993
rect -15084 26991 -15080 27015
rect -15074 27004 -15072 27014
rect -15056 27006 -15054 27012
rect -15050 27010 -15044 27020
rect -15036 27010 -15034 27304
rect -15030 27296 -15026 27304
rect -15002 27296 -14994 27304
rect -14954 27296 -14948 27304
rect -15003 27082 -14993 27104
rect -14952 27079 -14944 27090
rect -14940 27087 -14938 27304
rect -14926 27296 -14920 27304
rect -14960 27074 -14952 27079
rect -14950 27074 -14944 27079
rect -14942 27074 -14935 27087
rect -14920 27079 -14917 27092
rect -14950 27049 -14943 27074
rect -14940 27049 -14938 27074
rect -15000 27038 -14986 27046
rect -14942 27024 -14935 27049
rect -14928 27039 -14924 27049
rect -14916 27039 -14914 27304
rect -14894 27079 -14890 27081
rect -14896 27071 -14890 27079
rect -14895 27049 -14890 27051
rect -14884 27049 -14878 27071
rect -14868 27056 -14866 27317
rect -14820 27312 -14818 27317
rect -14724 27312 -14722 27317
rect -14700 27312 -14698 27317
rect -14854 27304 -14844 27312
rect -14826 27304 -14816 27312
rect -14794 27304 -14786 27312
rect -14732 27304 -14722 27312
rect -14704 27304 -14694 27312
rect -14860 27296 -14854 27304
rect -14832 27296 -14826 27304
rect -14863 27083 -14854 27084
rect -14844 27083 -14837 27084
rect -14830 27083 -14829 27279
rect -14820 27083 -14818 27304
rect -14786 27296 -14778 27304
rect -14738 27296 -14732 27304
rect -14863 27082 -14832 27083
rect -14830 27082 -14802 27083
rect -14787 27082 -14777 27104
rect -14870 27046 -14866 27056
rect -15060 27004 -15054 27006
rect -15176 26989 -15174 26990
rect -15084 26987 -15082 26991
rect -15064 26990 -15062 27004
rect -15056 26996 -15050 27004
rect -15040 26996 -15034 27010
rect -14961 27002 -14954 27014
rect -14940 27008 -14938 27024
rect -14920 27023 -14914 27039
rect -14918 27009 -14914 27023
rect -15036 26987 -15034 26996
rect -14942 26987 -14935 27008
rect -14916 26987 -14914 27009
rect -14868 26987 -14866 27046
rect -14860 27041 -14858 27046
rect -14840 27041 -14836 27056
rect -14832 27041 -14830 27071
rect -14820 27041 -14818 27082
rect -14736 27079 -14728 27090
rect -14724 27087 -14722 27304
rect -14710 27296 -14704 27304
rect -14744 27074 -14736 27079
rect -14734 27074 -14728 27079
rect -14726 27074 -14719 27087
rect -14704 27079 -14701 27092
rect -14815 27041 -14814 27071
rect -14734 27049 -14727 27074
rect -14724 27049 -14722 27074
rect -14854 27036 -14818 27041
rect -14784 27038 -14770 27046
rect -14854 27032 -14846 27036
rect -14840 27032 -14836 27036
rect -14854 27031 -14850 27032
rect -14844 27015 -14840 27031
rect -14842 27012 -14840 27015
rect -14834 27012 -14828 27020
rect -14842 27001 -14828 27012
rect -14820 27010 -14818 27036
rect -14726 27024 -14719 27049
rect -14712 27039 -14708 27049
rect -14700 27039 -14698 27304
rect -14678 27079 -14674 27081
rect -14680 27071 -14674 27079
rect -14679 27049 -14674 27051
rect -14668 27049 -14662 27071
rect -14652 27067 -14650 27317
rect -14604 27312 -14602 27317
rect -14508 27312 -14506 27317
rect -14484 27312 -14482 27317
rect -14634 27304 -14628 27312
rect -14606 27304 -14600 27312
rect -14574 27304 -14566 27312
rect -14546 27304 -14532 27312
rect -14516 27304 -14504 27312
rect -14488 27304 -14476 27312
rect -14644 27296 -14634 27304
rect -14616 27296 -14606 27304
rect -14624 27132 -14614 27141
rect -14614 27125 -14608 27132
rect -14661 27057 -14650 27067
rect -14604 27065 -14602 27304
rect -14566 27296 -14558 27304
rect -14532 27296 -14530 27304
rect -14518 27296 -14516 27304
rect -14538 27079 -14532 27089
rect -14633 27057 -14626 27065
rect -14824 26996 -14818 27010
rect -14745 27002 -14738 27014
rect -14724 27008 -14722 27024
rect -14704 27023 -14698 27039
rect -14702 27009 -14698 27023
rect -14820 26987 -14818 26996
rect -14726 26987 -14719 27008
rect -14700 26987 -14698 27009
rect -14652 27041 -14642 27057
rect -14652 27027 -14643 27041
rect -14638 27031 -14635 27041
rect -14623 27031 -14616 27057
rect -14614 27041 -14608 27057
rect -14606 27041 -14599 27065
rect -14628 27027 -14612 27031
rect -14604 27027 -14602 27041
rect -14652 27023 -14648 27027
rect -14652 26987 -14649 27023
rect -14606 27015 -14602 27027
rect -14575 27019 -14572 27049
rect -14570 27027 -14559 27049
rect -14557 27027 -14554 27057
rect -14539 27049 -14532 27059
rect -14528 27049 -14522 27079
rect -14508 27049 -14506 27304
rect -14504 27296 -14502 27304
rect -14490 27296 -14488 27304
rect -14503 27049 -14496 27057
rect -14484 27049 -14482 27304
rect -14476 27296 -14474 27304
rect -14462 27079 -14458 27081
rect -14464 27071 -14458 27079
rect -14474 27049 -14468 27059
rect -14463 27049 -14458 27051
rect -14452 27049 -14446 27071
rect -14436 27067 -14434 27317
rect -14388 27312 -14386 27317
rect -14268 27312 -14266 27317
rect -14172 27312 -14170 27317
rect -14076 27312 -14074 27317
rect -14028 27312 -14026 27317
rect -14418 27304 -14412 27312
rect -14390 27304 -14384 27312
rect -14358 27304 -14350 27312
rect -14330 27304 -14314 27312
rect -14298 27304 -14286 27312
rect -14270 27304 -14258 27312
rect -14238 27304 -14230 27312
rect -14210 27304 -14194 27312
rect -14178 27304 -14166 27312
rect -14150 27304 -14138 27312
rect -14118 27304 -14110 27312
rect -14090 27304 -14074 27312
rect -14060 27304 -14048 27312
rect -14032 27304 -14020 27312
rect -14428 27296 -14418 27304
rect -14400 27296 -14390 27304
rect -14408 27132 -14398 27141
rect -14398 27125 -14392 27132
rect -14445 27057 -14434 27067
rect -14388 27065 -14386 27304
rect -14350 27296 -14342 27304
rect -14302 27296 -14298 27304
rect -14274 27296 -14270 27304
rect -14417 27057 -14410 27065
rect -14548 27019 -14544 27027
rect -14529 27019 -14522 27049
rect -14510 27019 -14503 27049
rect -14496 27039 -14492 27049
rect -14484 27039 -14478 27049
rect -14488 27023 -14478 27039
rect -14486 27019 -14478 27023
rect -14436 27041 -14426 27057
rect -14436 27027 -14427 27041
rect -14422 27031 -14419 27041
rect -14407 27031 -14400 27057
rect -14398 27041 -14392 27057
rect -14390 27041 -14383 27065
rect -14325 27057 -14316 27067
rect -14412 27027 -14396 27031
rect -14388 27027 -14386 27041
rect -14436 27023 -14432 27027
rect -14623 26987 -14616 27015
rect -14604 26987 -14602 27015
rect -14564 26987 -14555 27019
rect -14508 26987 -14506 27019
rect -14486 27009 -14482 27019
rect -14484 27001 -14482 27009
rect -14488 26987 -14482 27001
rect -14436 26987 -14433 27023
rect -14390 27015 -14386 27027
rect -14359 27019 -14356 27049
rect -14354 27027 -14343 27049
rect -14341 27027 -14338 27057
rect -14332 27019 -14328 27027
rect -14315 27019 -14306 27057
rect -14287 27027 -14280 27057
rect -14268 27049 -14266 27304
rect -14230 27296 -14222 27304
rect -14182 27296 -14178 27304
rect -14278 27027 -14272 27049
rect -14297 27019 -14290 27027
rect -14270 27019 -14263 27049
rect -14239 27019 -14236 27049
rect -14234 27027 -14223 27049
rect -14221 27027 -14218 27057
rect -14212 27019 -14208 27027
rect -14407 26987 -14400 27015
rect -14388 26987 -14386 27015
rect -14348 26987 -14339 27019
rect -14287 26987 -14280 27019
rect -14268 26987 -14266 27019
rect -14228 26987 -14219 27019
rect -14172 26987 -14170 27304
rect -14154 27296 -14150 27304
rect -14110 27296 -14102 27304
rect -14167 27048 -14160 27057
rect -14152 27049 -14142 27064
rect -14076 27059 -14074 27304
rect -14062 27296 -14060 27304
rect -14048 27296 -14046 27304
rect -14034 27296 -14032 27304
rect -14065 27083 -14049 27091
rect -14158 27048 -14152 27049
rect -14150 27019 -14143 27049
rect -14141 27048 -14132 27059
rect -14083 27049 -14074 27059
rect -14072 27049 -14066 27079
rect -14065 27077 -14054 27079
rect -14065 27049 -14056 27070
rect -14152 26987 -14148 27019
rect -14076 27015 -14074 27049
rect -14073 27040 -14066 27049
rect -14054 27040 -14049 27070
rect -14073 27015 -14072 27040
rect -14040 27039 -14036 27049
rect -14028 27039 -14026 27304
rect -14020 27296 -14018 27304
rect -14006 27079 -14002 27081
rect -14008 27071 -14002 27079
rect -14007 27049 -14002 27051
rect -13996 27049 -13990 27071
rect -13980 27059 -13978 27317
rect -13956 27312 -13954 27317
rect -13932 27312 -13930 27317
rect -13860 27312 -13858 27317
rect -13964 27304 -13954 27312
rect -13936 27304 -13928 27312
rect -13866 27304 -13858 27312
rect -13838 27304 -13832 27312
rect -13806 27304 -13798 27312
rect -13778 27304 -13766 27312
rect -13764 27304 -13762 27317
rect -13716 27312 -13714 27317
rect -13750 27304 -13738 27312
rect -13722 27304 -13710 27312
rect -13690 27304 -13682 27312
rect -13972 27296 -13964 27304
rect -13987 27049 -13978 27059
rect -13976 27049 -13970 27079
rect -13956 27049 -13954 27304
rect -13944 27296 -13936 27304
rect -13951 27071 -13944 27079
rect -13932 27071 -13930 27304
rect -13876 27296 -13866 27304
rect -13922 27149 -13916 27279
rect -13922 27133 -13914 27149
rect -13932 27049 -13926 27071
rect -13922 27049 -13916 27133
rect -13910 27079 -13906 27081
rect -13912 27071 -13906 27079
rect -13911 27049 -13906 27051
rect -13900 27049 -13894 27071
rect -14076 26991 -14072 27015
rect -14066 27004 -14064 27014
rect -14054 27004 -14047 27015
rect -14030 27009 -14026 27039
rect -14076 26987 -14074 26991
rect -14073 26987 -14072 26991
rect -14056 26991 -14047 27004
rect -14042 26991 -14038 27004
rect -14056 26990 -14042 26991
rect -14054 26989 -14046 26990
rect -14028 26987 -14026 27009
rect -13980 26987 -13978 27049
rect -13977 27041 -13970 27049
rect -13958 27041 -13951 27049
rect -13946 27041 -13926 27049
rect -13977 27023 -13976 27041
rect -13956 26993 -13954 27041
rect -13946 27039 -13940 27041
rect -13932 27039 -13930 27041
rect -13936 27023 -13930 27039
rect -13934 27009 -13930 27023
rect -13956 26987 -13952 26993
rect -13932 26987 -13930 27009
rect -13860 27013 -13858 27304
rect -13848 27296 -13838 27304
rect -13798 27296 -13790 27304
rect -13766 27296 -13762 27304
rect -13738 27296 -13734 27304
rect -13855 27048 -13848 27078
rect -13846 27048 -13840 27071
rect -13838 27041 -13831 27071
rect -13829 27048 -13820 27279
rect -13764 27056 -13762 27296
rect -13764 27055 -13753 27056
rect -13846 27013 -13844 27023
rect -13838 27015 -13834 27041
rect -13764 27025 -13755 27055
rect -13753 27040 -13747 27055
rect -13745 27040 -13738 27063
rect -13860 27001 -13846 27013
rect -13836 27001 -13834 27013
rect -13860 26993 -13858 27001
rect -13860 26987 -13856 26993
rect -13764 26987 -13760 27025
rect -13754 27004 -13752 27014
rect -13744 27002 -13742 27004
rect -13730 27002 -13728 27004
rect -13744 26998 -13730 27002
rect -13754 26990 -13730 26998
rect -13754 26989 -13744 26990
rect -13742 26989 -13734 26990
rect -13716 26987 -13714 27304
rect -13710 27296 -13706 27304
rect -13682 27296 -13674 27304
rect -13644 27055 -13642 27317
rect -13596 27312 -13594 27317
rect -13500 27312 -13498 27317
rect -13404 27312 -13402 27317
rect -13356 27312 -13354 27317
rect -13284 27312 -13282 27317
rect -13626 27304 -13618 27312
rect -13598 27304 -13590 27312
rect -13566 27304 -13558 27312
rect -13538 27304 -13522 27312
rect -13506 27304 -13494 27312
rect -13478 27304 -13466 27312
rect -13446 27304 -13438 27312
rect -13418 27304 -13402 27312
rect -13388 27304 -13376 27312
rect -13360 27304 -13348 27312
rect -13290 27304 -13282 27312
rect -13262 27304 -13256 27312
rect -13230 27304 -13222 27312
rect -13202 27304 -13186 27312
rect -13170 27304 -13158 27312
rect -13142 27304 -13130 27312
rect -13110 27304 -13102 27312
rect -13082 27304 -13066 27312
rect -13050 27304 -13038 27312
rect -13022 27304 -13010 27312
rect -12990 27304 -12982 27312
rect -12962 27304 -12946 27312
rect -12930 27304 -12918 27312
rect -12902 27304 -12890 27312
rect -12870 27304 -12862 27312
rect -12842 27304 -12830 27312
rect -12828 27304 -12826 27317
rect -12780 27312 -12778 27317
rect -12684 27312 -12682 27317
rect -12660 27312 -12658 27317
rect -12814 27304 -12802 27312
rect -12786 27304 -12774 27312
rect -12754 27304 -12746 27312
rect -12692 27304 -12682 27312
rect -12664 27304 -12654 27312
rect -13634 27296 -13626 27304
rect -13606 27296 -13598 27304
rect -13616 27116 -13600 27123
rect -13687 27020 -13684 27047
rect -13682 27025 -13671 27047
rect -13669 27025 -13666 27055
rect -13644 27027 -13635 27055
rect -13615 27027 -13608 27055
rect -13596 27047 -13594 27304
rect -13558 27296 -13550 27304
rect -13510 27296 -13506 27304
rect -13606 27027 -13600 27047
rect -13687 27017 -13675 27020
rect -13644 26987 -13642 27027
rect -13625 27017 -13618 27027
rect -13598 27017 -13591 27047
rect -13567 27019 -13564 27049
rect -13562 27027 -13551 27049
rect -13549 27027 -13546 27057
rect -13540 27019 -13536 27027
rect -13615 27007 -13608 27017
rect -13598 26991 -13594 27017
rect -13615 26987 -13608 26991
rect -13596 26987 -13594 26991
rect -13556 26987 -13547 27019
rect -13500 26987 -13498 27304
rect -13482 27296 -13478 27304
rect -13438 27296 -13430 27304
rect -13495 27048 -13488 27057
rect -13480 27049 -13470 27064
rect -13404 27059 -13402 27304
rect -13390 27296 -13388 27304
rect -13376 27296 -13374 27304
rect -13362 27296 -13360 27304
rect -13393 27083 -13377 27091
rect -13486 27048 -13480 27049
rect -13478 27019 -13471 27049
rect -13469 27048 -13460 27059
rect -13411 27049 -13402 27059
rect -13400 27049 -13394 27079
rect -13393 27077 -13382 27079
rect -13393 27049 -13384 27070
rect -13480 26987 -13476 27019
rect -13404 27015 -13402 27049
rect -13401 27040 -13394 27049
rect -13382 27040 -13377 27070
rect -13401 27015 -13400 27040
rect -13368 27039 -13364 27049
rect -13356 27039 -13354 27304
rect -13348 27296 -13346 27304
rect -13300 27296 -13290 27304
rect -13334 27079 -13330 27081
rect -13336 27071 -13330 27079
rect -13335 27049 -13330 27051
rect -13324 27049 -13318 27071
rect -13404 26991 -13400 27015
rect -13394 27004 -13392 27014
rect -13382 27004 -13375 27015
rect -13358 27009 -13354 27039
rect -13404 26987 -13402 26991
rect -13401 26987 -13400 26991
rect -13384 26991 -13375 27004
rect -13370 26991 -13366 27004
rect -13384 26990 -13370 26991
rect -13382 26989 -13374 26990
rect -13356 26987 -13354 27009
rect -13284 27013 -13282 27304
rect -13272 27296 -13262 27304
rect -13222 27296 -13214 27304
rect -13174 27296 -13170 27304
rect -13146 27296 -13142 27304
rect -13102 27296 -13094 27304
rect -13054 27296 -13050 27304
rect -13026 27296 -13022 27304
rect -12982 27296 -12974 27304
rect -12934 27296 -12930 27304
rect -12906 27296 -12902 27304
rect -12862 27296 -12854 27304
rect -12830 27296 -12826 27304
rect -12802 27296 -12798 27304
rect -13279 27048 -13272 27078
rect -13270 27048 -13264 27071
rect -13262 27041 -13255 27071
rect -13253 27048 -13244 27279
rect -13172 27083 -13161 27090
rect -13052 27083 -13041 27090
rect -12932 27083 -12921 27090
rect -13170 27078 -13161 27083
rect -13050 27078 -13041 27083
rect -12930 27078 -12921 27083
rect -13160 27048 -13149 27078
rect -13040 27048 -13029 27078
rect -12920 27048 -12909 27078
rect -12828 27056 -12826 27296
rect -12817 27083 -12801 27099
rect -12823 27082 -12814 27083
rect -13270 27013 -13268 27023
rect -13262 27015 -13258 27041
rect -13160 27040 -13151 27048
rect -13040 27040 -13031 27048
rect -12920 27040 -12911 27048
rect -12830 27046 -12826 27056
rect -12828 27015 -12826 27046
rect -12820 27040 -12818 27046
rect -12817 27040 -12806 27046
rect -12802 27040 -12801 27070
rect -12800 27032 -12796 27040
rect -13160 27013 -13158 27015
rect -13040 27013 -13038 27015
rect -12920 27013 -12918 27015
rect -13284 27001 -13270 27013
rect -13260 27001 -13258 27013
rect -13168 27004 -13158 27013
rect -13048 27004 -13038 27013
rect -12928 27004 -12918 27013
rect -13284 26993 -13282 27001
rect -13164 26999 -13154 27004
rect -13044 26999 -13034 27004
rect -12924 26999 -12914 27004
rect -13284 26987 -13280 26993
rect -12828 26991 -12824 27015
rect -12818 27004 -12816 27014
rect -12800 27006 -12798 27012
rect -12794 27010 -12788 27020
rect -12780 27010 -12778 27304
rect -12774 27296 -12770 27304
rect -12746 27296 -12738 27304
rect -12698 27296 -12692 27304
rect -12747 27082 -12737 27104
rect -12696 27079 -12688 27090
rect -12684 27087 -12682 27304
rect -12670 27296 -12664 27304
rect -12704 27074 -12696 27079
rect -12694 27074 -12688 27079
rect -12686 27074 -12679 27087
rect -12664 27079 -12661 27092
rect -12694 27049 -12687 27074
rect -12684 27049 -12682 27074
rect -12744 27038 -12730 27046
rect -12686 27024 -12679 27049
rect -12672 27039 -12668 27049
rect -12660 27039 -12658 27304
rect -12638 27079 -12634 27081
rect -12640 27071 -12634 27079
rect -12639 27049 -12634 27051
rect -12628 27049 -12622 27071
rect -12612 27059 -12610 27317
rect -12588 27312 -12586 27317
rect -12564 27312 -12562 27317
rect -12492 27312 -12490 27317
rect -12596 27304 -12586 27312
rect -12568 27304 -12560 27312
rect -12498 27304 -12490 27312
rect -12470 27304 -12464 27312
rect -12438 27304 -12430 27312
rect -12410 27304 -12398 27312
rect -12396 27304 -12394 27317
rect -12348 27312 -12346 27317
rect -12382 27304 -12370 27312
rect -12354 27304 -12342 27312
rect -12322 27304 -12314 27312
rect -12604 27296 -12596 27304
rect -12619 27049 -12610 27059
rect -12608 27049 -12602 27079
rect -12588 27049 -12586 27304
rect -12576 27296 -12568 27304
rect -12583 27071 -12576 27079
rect -12564 27071 -12562 27304
rect -12508 27296 -12498 27304
rect -12554 27149 -12548 27279
rect -12554 27133 -12546 27149
rect -12564 27049 -12558 27071
rect -12554 27049 -12548 27133
rect -12542 27079 -12538 27081
rect -12544 27071 -12538 27079
rect -12543 27049 -12538 27051
rect -12532 27049 -12526 27071
rect -12804 27004 -12798 27006
rect -13160 26989 -13158 26990
rect -13040 26989 -13038 26990
rect -12920 26989 -12918 26990
rect -12828 26987 -12826 26991
rect -12808 26990 -12806 27004
rect -12800 26996 -12794 27004
rect -12784 26996 -12778 27010
rect -12705 27002 -12698 27014
rect -12684 27008 -12682 27024
rect -12664 27023 -12658 27039
rect -12662 27009 -12658 27023
rect -12780 26987 -12778 26996
rect -12686 26987 -12679 27008
rect -12660 26987 -12658 27009
rect -12612 26987 -12610 27049
rect -12609 27041 -12602 27049
rect -12590 27041 -12583 27049
rect -12578 27041 -12558 27049
rect -12609 27023 -12608 27041
rect -12588 26993 -12586 27041
rect -12578 27039 -12572 27041
rect -12564 27039 -12562 27041
rect -12568 27023 -12562 27039
rect -12566 27009 -12562 27023
rect -12588 26987 -12584 26993
rect -12564 26987 -12562 27009
rect -12492 27013 -12490 27304
rect -12480 27296 -12470 27304
rect -12430 27296 -12422 27304
rect -12398 27296 -12394 27304
rect -12370 27296 -12366 27304
rect -12487 27048 -12480 27078
rect -12478 27048 -12472 27071
rect -12470 27041 -12463 27071
rect -12461 27048 -12452 27279
rect -12396 27056 -12394 27296
rect -12396 27055 -12385 27056
rect -12478 27013 -12476 27023
rect -12470 27015 -12466 27041
rect -12396 27025 -12387 27055
rect -12385 27040 -12379 27055
rect -12377 27040 -12370 27063
rect -12492 27001 -12478 27013
rect -12468 27001 -12466 27013
rect -12492 26993 -12490 27001
rect -12492 26987 -12488 26993
rect -12396 26987 -12392 27025
rect -12386 27004 -12384 27014
rect -12376 27002 -12374 27004
rect -12362 27002 -12360 27004
rect -12376 26998 -12362 27002
rect -12386 26990 -12362 26998
rect -12386 26989 -12376 26990
rect -12374 26989 -12366 26990
rect -12348 26987 -12346 27304
rect -12342 27296 -12338 27304
rect -12314 27296 -12306 27304
rect -12319 27020 -12316 27047
rect -12314 27025 -12303 27047
rect -12301 27025 -12298 27055
rect -12319 27017 -12307 27020
rect -12276 26987 -12274 27317
rect -12252 27312 -12250 27317
rect -12228 27312 -12226 27317
rect -12156 27312 -12154 27317
rect -12260 27304 -12250 27312
rect -12232 27304 -12222 27312
rect -12162 27304 -12154 27312
rect -12134 27304 -12128 27312
rect -12102 27304 -12094 27312
rect -12074 27304 -12062 27312
rect -12060 27304 -12058 27317
rect -12012 27312 -12010 27317
rect -11916 27312 -11914 27317
rect -11892 27312 -11890 27317
rect -12046 27304 -12034 27312
rect -12018 27304 -12006 27312
rect -11986 27304 -11978 27312
rect -11924 27304 -11914 27312
rect -11896 27304 -11886 27312
rect -12266 27296 -12260 27304
rect -12272 27049 -12254 27059
rect -12252 27047 -12250 27304
rect -12238 27296 -12232 27304
rect -12228 27059 -12226 27304
rect -12172 27296 -12162 27304
rect -12247 27049 -12226 27059
rect -12218 27049 -12212 27279
rect -12206 27079 -12202 27081
rect -12208 27071 -12202 27079
rect -12207 27049 -12202 27051
rect -12196 27049 -12190 27071
rect -12254 27017 -12247 27047
rect -12240 27039 -12236 27049
rect -12228 27047 -12226 27049
rect -12228 27039 -12222 27047
rect -12232 27023 -12222 27039
rect -12230 27017 -12222 27023
rect -12252 26991 -12250 27017
rect -12230 27009 -12226 27017
rect -12252 26987 -12238 26991
rect -12228 26987 -12226 27009
rect -12156 27013 -12154 27304
rect -12144 27296 -12134 27304
rect -12094 27296 -12086 27304
rect -12062 27296 -12058 27304
rect -12034 27296 -12030 27304
rect -12151 27048 -12144 27078
rect -12142 27048 -12136 27071
rect -12134 27041 -12127 27071
rect -12125 27048 -12116 27279
rect -12060 27056 -12058 27296
rect -12049 27083 -12033 27099
rect -12055 27082 -12046 27083
rect -12062 27046 -12058 27056
rect -12142 27013 -12140 27023
rect -12134 27015 -12130 27041
rect -12060 27015 -12058 27046
rect -12052 27040 -12050 27046
rect -12049 27040 -12038 27046
rect -12034 27040 -12033 27070
rect -12032 27032 -12028 27040
rect -12156 27001 -12142 27013
rect -12132 27001 -12130 27013
rect -12156 26993 -12154 27001
rect -12156 26987 -12152 26993
rect -12060 26991 -12056 27015
rect -12050 27004 -12048 27014
rect -12032 27006 -12030 27012
rect -12026 27010 -12020 27020
rect -12012 27010 -12010 27304
rect -12006 27296 -12002 27304
rect -11978 27296 -11970 27304
rect -11930 27296 -11924 27304
rect -11979 27082 -11969 27104
rect -11928 27079 -11920 27090
rect -11916 27087 -11914 27304
rect -11902 27296 -11896 27304
rect -11936 27074 -11928 27079
rect -11926 27074 -11920 27079
rect -11918 27074 -11911 27087
rect -11896 27079 -11893 27092
rect -11926 27049 -11919 27074
rect -11916 27049 -11914 27074
rect -11976 27038 -11962 27046
rect -11918 27024 -11911 27049
rect -11904 27039 -11900 27049
rect -11892 27039 -11890 27304
rect -11870 27079 -11866 27081
rect -11872 27071 -11866 27079
rect -11871 27049 -11866 27051
rect -11860 27049 -11854 27071
rect -11844 27056 -11842 27317
rect -11796 27312 -11794 27317
rect -11676 27312 -11674 27317
rect -11580 27312 -11578 27317
rect -11556 27312 -11554 27317
rect -11830 27304 -11820 27312
rect -11802 27304 -11792 27312
rect -11770 27304 -11762 27312
rect -11742 27304 -11726 27312
rect -11710 27304 -11698 27312
rect -11682 27304 -11670 27312
rect -11650 27304 -11642 27312
rect -11622 27304 -11606 27312
rect -11590 27304 -11578 27312
rect -11562 27304 -11550 27312
rect -11530 27304 -11522 27312
rect -11836 27296 -11830 27304
rect -11808 27296 -11802 27304
rect -11839 27083 -11830 27084
rect -11820 27083 -11813 27084
rect -11806 27083 -11805 27279
rect -11796 27083 -11794 27304
rect -11762 27296 -11754 27304
rect -11714 27296 -11710 27304
rect -11686 27296 -11682 27304
rect -11698 27116 -11682 27124
rect -11839 27082 -11808 27083
rect -11806 27082 -11778 27083
rect -11763 27082 -11753 27104
rect -11719 27082 -11712 27104
rect -11710 27082 -11703 27112
rect -11698 27110 -11693 27112
rect -11686 27110 -11682 27112
rect -11701 27082 -11695 27104
rect -11846 27046 -11842 27056
rect -12036 27004 -12030 27006
rect -12060 26987 -12058 26991
rect -12040 26990 -12038 27004
rect -12032 26996 -12026 27004
rect -12016 26996 -12010 27010
rect -11937 27002 -11930 27014
rect -11916 27008 -11914 27024
rect -11896 27023 -11890 27039
rect -11894 27009 -11890 27023
rect -12012 26987 -12010 26996
rect -11918 26987 -11911 27008
rect -11892 26987 -11890 27009
rect -11844 26987 -11842 27046
rect -11836 27041 -11834 27046
rect -11816 27041 -11812 27056
rect -11808 27041 -11806 27071
rect -11796 27041 -11794 27082
rect -11693 27074 -11686 27104
rect -11684 27082 -11677 27104
rect -11791 27041 -11790 27071
rect -11726 27046 -11718 27056
rect -11830 27036 -11794 27041
rect -11760 27038 -11746 27046
rect -11716 27038 -11702 27046
rect -11696 27038 -11692 27056
rect -11830 27032 -11822 27036
rect -11816 27032 -11812 27036
rect -11830 27031 -11826 27032
rect -11820 27015 -11816 27031
rect -11818 27012 -11816 27015
rect -11810 27012 -11804 27020
rect -11818 27001 -11804 27012
rect -11796 27010 -11794 27036
rect -11716 27034 -11708 27038
rect -11716 27032 -11702 27034
rect -11698 27032 -11692 27038
rect -11716 27028 -11706 27032
rect -11710 27024 -11706 27028
rect -11698 27024 -11696 27032
rect -11800 26996 -11794 27010
rect -11716 27002 -11714 27014
rect -11700 27012 -11696 27024
rect -11684 27020 -11680 27024
rect -11690 27012 -11680 27020
rect -11700 27008 -11684 27012
rect -11676 27010 -11674 27304
rect -11642 27296 -11634 27304
rect -11594 27296 -11590 27304
rect -11643 27082 -11633 27104
rect -11640 27038 -11626 27046
rect -11590 27025 -11585 27055
rect -11580 27029 -11578 27304
rect -11566 27296 -11562 27304
rect -11556 27034 -11554 27304
rect -11522 27296 -11514 27304
rect -11580 27027 -11559 27029
rect -11583 27025 -11559 27027
rect -11580 27012 -11578 27025
rect -11696 26996 -11693 27008
rect -11680 26996 -11674 27010
rect -11592 27002 -11588 27012
rect -11580 27008 -11564 27012
rect -11558 27008 -11554 27034
rect -11527 27020 -11524 27047
rect -11522 27025 -11511 27047
rect -11509 27025 -11506 27055
rect -11527 27017 -11515 27020
rect -11580 27002 -11578 27008
rect -11796 26987 -11794 26996
rect -11676 26987 -11674 26996
rect -11594 26988 -11590 26998
rect -11582 26988 -11578 27002
rect -11581 26987 -11578 26988
rect -11556 26987 -11554 27008
rect -11484 26987 -11482 27317
rect -11460 27312 -11458 27317
rect -11436 27312 -11434 27317
rect -11468 27304 -11458 27312
rect -11440 27304 -11430 27312
rect -11474 27296 -11468 27304
rect -11480 27049 -11462 27059
rect -11460 27047 -11458 27304
rect -11446 27296 -11440 27304
rect -11436 27059 -11434 27304
rect -11455 27049 -11434 27059
rect -11426 27049 -11420 27279
rect -11414 27079 -11410 27081
rect -11416 27071 -11410 27079
rect -11415 27049 -11410 27051
rect -11404 27049 -11398 27071
rect -11388 27059 -11386 27317
rect -11364 27312 -11362 27317
rect -11340 27312 -11338 27317
rect -11268 27312 -11266 27317
rect -11172 27312 -11170 27317
rect -11124 27312 -11122 27317
rect -11372 27304 -11362 27312
rect -11344 27304 -11336 27312
rect -11274 27304 -11266 27312
rect -11246 27304 -11240 27312
rect -11214 27304 -11206 27312
rect -11186 27304 -11170 27312
rect -11156 27304 -11144 27312
rect -11128 27304 -11116 27312
rect -11380 27296 -11372 27304
rect -11395 27049 -11386 27059
rect -11384 27049 -11378 27079
rect -11364 27049 -11362 27304
rect -11352 27296 -11344 27304
rect -11359 27071 -11352 27079
rect -11340 27071 -11338 27304
rect -11284 27296 -11274 27304
rect -11330 27149 -11324 27279
rect -11330 27133 -11322 27149
rect -11340 27049 -11334 27071
rect -11330 27049 -11324 27133
rect -11318 27079 -11314 27081
rect -11320 27071 -11314 27079
rect -11319 27049 -11314 27051
rect -11308 27049 -11302 27071
rect -11462 27017 -11455 27047
rect -11448 27039 -11444 27049
rect -11436 27047 -11434 27049
rect -11436 27039 -11430 27047
rect -11440 27023 -11430 27039
rect -11438 27017 -11430 27023
rect -11460 26991 -11458 27017
rect -11438 27009 -11434 27017
rect -11460 26987 -11446 26991
rect -11436 26987 -11434 27009
rect -11388 26987 -11386 27049
rect -11385 27041 -11378 27049
rect -11366 27041 -11359 27049
rect -11354 27041 -11334 27049
rect -11385 27023 -11384 27041
rect -11364 26993 -11362 27041
rect -11354 27039 -11348 27041
rect -11340 27039 -11338 27041
rect -11344 27023 -11338 27039
rect -11342 27009 -11338 27023
rect -11364 26987 -11360 26993
rect -11340 26987 -11338 27009
rect -11268 27013 -11266 27304
rect -11256 27296 -11246 27304
rect -11206 27296 -11198 27304
rect -11263 27048 -11256 27078
rect -11254 27048 -11248 27071
rect -11246 27041 -11239 27071
rect -11237 27048 -11228 27279
rect -11172 27059 -11170 27304
rect -11158 27296 -11156 27304
rect -11144 27296 -11142 27304
rect -11130 27296 -11128 27304
rect -11161 27083 -11145 27091
rect -11179 27049 -11170 27059
rect -11168 27049 -11162 27079
rect -11161 27077 -11150 27079
rect -11161 27049 -11152 27070
rect -11254 27013 -11252 27023
rect -11246 27015 -11242 27041
rect -11172 27015 -11170 27049
rect -11169 27040 -11162 27049
rect -11150 27040 -11145 27070
rect -11169 27015 -11168 27040
rect -11136 27039 -11132 27049
rect -11124 27039 -11122 27304
rect -11116 27296 -11114 27304
rect -11102 27079 -11098 27081
rect -11104 27071 -11098 27079
rect -11103 27049 -11098 27051
rect -11092 27049 -11086 27071
rect -11076 27067 -11074 27317
rect -11028 27312 -11026 27317
rect -10932 27312 -10930 27317
rect -11058 27304 -11052 27312
rect -11030 27304 -11024 27312
rect -10998 27304 -10990 27312
rect -10970 27304 -10954 27312
rect -10938 27304 -10926 27312
rect -10910 27304 -10898 27312
rect -10878 27304 -10870 27312
rect -10850 27304 -10838 27312
rect -10836 27304 -10834 27317
rect -10788 27312 -10786 27317
rect -10668 27312 -10666 27317
rect -10179 27314 -10163 27317
rect -10822 27304 -10810 27312
rect -10794 27304 -10782 27312
rect -10762 27304 -10754 27312
rect -10734 27304 -10718 27312
rect -10702 27304 -10690 27312
rect -10674 27304 -10662 27312
rect -10642 27304 -10634 27312
rect -10614 27304 -10598 27312
rect -10581 27304 -10570 27312
rect -10552 27304 -10542 27312
rect -10521 27304 -10511 27312
rect -10492 27304 -10483 27312
rect -10463 27304 -10455 27312
rect -10435 27304 -10427 27312
rect -10407 27304 -10398 27312
rect -10379 27304 -10370 27312
rect -10350 27304 -10342 27312
rect -10322 27304 -10314 27312
rect -10294 27304 -10286 27312
rect -10266 27304 -10258 27312
rect -10238 27304 -10230 27312
rect -10210 27304 -10202 27312
rect -10016 27309 -10014 27317
rect -10154 27304 -10146 27309
rect -10126 27304 -10118 27309
rect -11068 27296 -11058 27304
rect -11040 27296 -11030 27304
rect -11048 27132 -11038 27141
rect -11038 27125 -11032 27132
rect -11085 27057 -11074 27067
rect -11028 27065 -11026 27304
rect -10990 27296 -10982 27304
rect -10942 27296 -10938 27304
rect -11057 27057 -11050 27065
rect -11268 27001 -11254 27013
rect -11244 27001 -11242 27013
rect -11268 26993 -11266 27001
rect -11268 26987 -11264 26993
rect -11172 26991 -11168 27015
rect -11162 27004 -11160 27014
rect -11150 27004 -11143 27015
rect -11126 27009 -11122 27039
rect -11172 26987 -11170 26991
rect -11169 26987 -11168 26991
rect -11152 26991 -11143 27004
rect -11138 26991 -11134 27004
rect -11152 26990 -11138 26991
rect -11150 26989 -11142 26990
rect -11124 26987 -11122 27009
rect -11076 27041 -11066 27057
rect -11076 27027 -11067 27041
rect -11062 27031 -11059 27041
rect -11047 27031 -11040 27057
rect -11038 27041 -11032 27057
rect -11030 27041 -11023 27065
rect -11052 27027 -11036 27031
rect -11028 27027 -11026 27041
rect -11076 27023 -11072 27027
rect -11076 26987 -11073 27023
rect -11030 27015 -11026 27027
rect -10999 27019 -10996 27049
rect -10994 27027 -10983 27049
rect -10981 27027 -10978 27057
rect -10972 27019 -10968 27027
rect -11047 26987 -11040 27015
rect -11028 26987 -11026 27015
rect -10988 26987 -10979 27019
rect -10932 26987 -10930 27304
rect -10914 27296 -10910 27304
rect -10870 27296 -10862 27304
rect -10838 27296 -10834 27304
rect -10810 27296 -10806 27304
rect -10927 27048 -10920 27057
rect -10912 27049 -10902 27064
rect -10918 27048 -10912 27049
rect -10910 27019 -10903 27049
rect -10901 27048 -10892 27059
rect -10836 27056 -10834 27296
rect -10825 27083 -10809 27099
rect -10831 27082 -10822 27083
rect -10838 27046 -10834 27056
rect -10912 26987 -10908 27019
rect -10836 27015 -10834 27046
rect -10828 27040 -10826 27046
rect -10825 27040 -10814 27046
rect -10810 27040 -10809 27070
rect -10808 27032 -10804 27040
rect -10836 26991 -10832 27015
rect -10826 27004 -10824 27014
rect -10808 27006 -10806 27012
rect -10802 27010 -10796 27020
rect -10788 27010 -10786 27304
rect -10782 27296 -10778 27304
rect -10754 27296 -10746 27304
rect -10706 27296 -10702 27304
rect -10678 27296 -10674 27304
rect -10690 27116 -10674 27124
rect -10755 27082 -10745 27104
rect -10711 27082 -10704 27104
rect -10702 27082 -10695 27112
rect -10690 27110 -10685 27112
rect -10678 27110 -10674 27112
rect -10693 27082 -10687 27104
rect -10685 27074 -10678 27104
rect -10676 27082 -10669 27104
rect -10718 27046 -10710 27056
rect -10752 27038 -10738 27046
rect -10708 27038 -10694 27046
rect -10688 27038 -10684 27056
rect -10708 27034 -10700 27038
rect -10708 27032 -10694 27034
rect -10690 27032 -10684 27038
rect -10708 27028 -10698 27032
rect -10702 27024 -10698 27028
rect -10690 27024 -10688 27032
rect -10812 27004 -10806 27006
rect -10836 26987 -10834 26991
rect -10816 26990 -10814 27004
rect -10808 26996 -10802 27004
rect -10792 26996 -10786 27010
rect -10708 27002 -10706 27014
rect -10692 27012 -10688 27024
rect -10676 27020 -10672 27024
rect -10682 27012 -10672 27020
rect -10692 27008 -10676 27012
rect -10668 27010 -10666 27304
rect -10634 27296 -10626 27304
rect -10586 27296 -10581 27304
rect -10558 27296 -10552 27304
rect -10511 27296 -10505 27304
rect -10483 27296 -10476 27304
rect -10455 27296 -10447 27304
rect -10427 27296 -10419 27304
rect -10398 27296 -10391 27304
rect -10370 27296 -10363 27304
rect -10342 27296 -10334 27304
rect -10314 27296 -10306 27304
rect -10286 27296 -10278 27304
rect -10258 27296 -10250 27304
rect -10230 27296 -10222 27304
rect -10202 27296 -10194 27304
rect -10146 27293 -10138 27304
rect -10118 27294 -10110 27304
rect -10070 27301 -10062 27309
rect -10042 27301 -10034 27309
rect -10016 27301 -10006 27309
rect -9986 27301 -9972 27312
rect -9956 27301 -9944 27312
rect -9928 27301 -9916 27312
rect -10062 27294 -10054 27301
rect -10034 27294 -10026 27301
rect -10126 27293 -10110 27294
rect -10070 27293 -10054 27294
rect -10042 27293 -10026 27294
rect -10016 27294 -10014 27301
rect -10006 27294 -9998 27301
rect -9972 27296 -9970 27301
rect -9958 27296 -9956 27301
rect -9944 27296 -9942 27301
rect -9930 27296 -9928 27301
rect -9916 27296 -9914 27301
rect -10016 27293 -9998 27294
rect -9986 27293 -9978 27294
rect -10466 27279 -10333 27287
rect -10328 27279 -10275 27287
rect -10318 27261 -10314 27270
rect -10250 27269 -10243 27278
rect -10267 27257 -10261 27262
rect -10242 27257 -10233 27269
rect -10271 27252 -10267 27257
rect -10242 27253 -10226 27257
rect -10225 27253 -10222 27257
rect -10493 27238 -10487 27246
rect -10456 27238 -10445 27242
rect -10483 27230 -10477 27238
rect -10502 27210 -10487 27230
rect -10456 27227 -10443 27238
rect -10418 27230 -10411 27238
rect -10427 27227 -10411 27230
rect -10380 27227 -10370 27249
rect -10502 27200 -10483 27210
rect -10476 27200 -10457 27210
rect -10483 27198 -10477 27200
rect -10436 27198 -10433 27227
rect -10427 27208 -10419 27227
rect -10353 27219 -10347 27249
rect -10312 27219 -10307 27249
rect -10271 27227 -10270 27252
rect -10238 27227 -10231 27253
rect -10431 27200 -10418 27208
rect -10483 27192 -10476 27198
rect -10483 27190 -10469 27192
rect -10483 27185 -10460 27190
rect -10558 27156 -10549 27166
rect -10494 27160 -10487 27170
rect -10476 27168 -10460 27185
rect -10450 27168 -10443 27198
rect -10429 27195 -10411 27198
rect -10436 27166 -10429 27190
rect -10421 27168 -10411 27195
rect -10238 27193 -10233 27227
rect -10201 27221 -10192 27222
rect -10195 27219 -10192 27221
rect -10360 27190 -10354 27193
rect -10476 27160 -10422 27166
rect -10421 27160 -10412 27168
rect -10395 27163 -10379 27190
rect -10360 27163 -10357 27190
rect -10354 27163 -10353 27190
rect -10319 27185 -10314 27193
rect -10319 27163 -10303 27185
rect -10297 27163 -10289 27185
rect -10395 27160 -10388 27163
rect -10353 27160 -10347 27163
rect -10562 27130 -10554 27132
rect -10562 27116 -10555 27130
rect -10548 27116 -10539 27156
rect -10486 27153 -10477 27160
rect -10319 27155 -10281 27163
rect -10250 27155 -10243 27185
rect -10238 27163 -10231 27193
rect -10016 27186 -10014 27293
rect -10229 27163 -10222 27185
rect -10217 27163 -10213 27185
rect -10229 27155 -10212 27163
rect -10128 27156 -10116 27172
rect -10635 27082 -10625 27104
rect -10578 27074 -10574 27114
rect -10562 27074 -10555 27104
rect -10548 27100 -10537 27116
rect -10486 27070 -10479 27153
rect -10436 27122 -10433 27133
rect -10354 27132 -10347 27148
rect -10345 27133 -10315 27140
rect -10238 27130 -10233 27155
rect -10037 27148 -10036 27164
rect -10021 27162 -10013 27186
rect -10222 27133 -10208 27140
rect -10436 27092 -10429 27122
rect -10319 27100 -10314 27130
rect -10278 27100 -10271 27130
rect -10250 27100 -10249 27122
rect -10238 27100 -10231 27130
rect -10265 27092 -10243 27100
rect -10217 27092 -10210 27122
rect -10159 27106 -10146 27122
rect -10141 27106 -10137 27136
rect -10059 27110 -10043 27126
rect -10050 27101 -10043 27110
rect -10038 27106 -10036 27128
rect -10021 27106 -10012 27146
rect -9914 27140 -9909 27279
rect -9914 27133 -9907 27140
rect -10067 27098 -10063 27101
rect -10052 27098 -10036 27101
rect -9914 27098 -9909 27133
rect -10436 27070 -10433 27092
rect -10238 27083 -10233 27092
rect -10502 27062 -10450 27070
rect -10443 27062 -10431 27070
rect -10387 27062 -10351 27070
rect -10632 27038 -10618 27046
rect -10688 26996 -10685 27008
rect -10672 26996 -10666 27010
rect -10788 26987 -10786 26996
rect -10668 26987 -10666 26996
rect -10486 26987 -10479 27062
rect -10436 27060 -10433 27062
rect -10450 27052 -10443 27060
rect -10450 27030 -10434 27052
rect -10418 27030 -10411 27060
rect -10360 27052 -10354 27060
rect -10319 27052 -10314 27060
rect -10238 27057 -10231 27083
rect -10238 27052 -10233 27057
rect -10377 27030 -10365 27052
rect -10360 27030 -10359 27052
rect -10354 27030 -10353 27052
rect -10314 27030 -10312 27052
rect -10301 27030 -10286 27052
rect -10353 27027 -10347 27030
rect -10381 27022 -10347 27027
rect -10312 27022 -10307 27030
rect -10250 27022 -10243 27052
rect -10217 27026 -10210 27052
rect -10208 27047 -10200 27082
rect -10129 27027 -10125 27043
rect -10124 27041 -10113 27043
rect -10077 27041 -10071 27098
rect -10058 27071 -10057 27073
rect -10050 27071 -10044 27098
rect -10001 27083 -9998 27091
rect -9991 27081 -9988 27083
rect -10061 27041 -10054 27071
rect -10048 27041 -10043 27063
rect -10038 27041 -10032 27063
rect -10030 27041 -10023 27071
rect -10021 27041 -10012 27081
rect -10011 27041 -10005 27063
rect -10003 27041 -9996 27071
rect -9991 27041 -9985 27081
rect -9968 27049 -9967 27079
rect -9952 27063 -9946 27065
rect -9943 27063 -9937 27079
rect -9914 27073 -9912 27093
rect -9902 27079 -9898 27081
rect -9962 27049 -9952 27063
rect -9950 27049 -9946 27063
rect -9944 27049 -9943 27063
rect -10114 27035 -10113 27041
rect -10050 27033 -10043 27041
rect -10021 27033 -10013 27041
rect -9950 27033 -9944 27049
rect -9923 27043 -9919 27063
rect -9914 27049 -9909 27073
rect -9904 27071 -9898 27079
rect -9903 27049 -9898 27051
rect -9892 27049 -9886 27071
rect -9876 27056 -9874 27317
rect -9828 27312 -9826 27317
rect -9732 27312 -9730 27317
rect -9708 27312 -9706 27317
rect -9612 27312 -9610 27317
rect -9516 27312 -9514 27317
rect -9468 27312 -9466 27317
rect -9862 27304 -9852 27312
rect -9834 27304 -9824 27312
rect -9802 27304 -9794 27312
rect -9774 27304 -9758 27312
rect -9742 27304 -9730 27312
rect -9714 27304 -9702 27312
rect -9682 27304 -9674 27312
rect -9618 27304 -9610 27312
rect -9590 27304 -9582 27312
rect -9558 27304 -9550 27312
rect -9530 27304 -9514 27312
rect -9500 27304 -9488 27312
rect -9472 27304 -9460 27312
rect -9868 27296 -9862 27304
rect -9840 27296 -9834 27304
rect -9871 27083 -9862 27084
rect -9852 27083 -9845 27084
rect -9838 27083 -9837 27279
rect -9828 27083 -9826 27304
rect -9794 27296 -9786 27304
rect -9746 27296 -9742 27304
rect -9871 27082 -9840 27083
rect -9838 27082 -9810 27083
rect -9795 27082 -9785 27104
rect -9878 27046 -9874 27056
rect -9923 27039 -9918 27043
rect -9928 27033 -9919 27039
rect -10226 27022 -10210 27026
rect -10436 26987 -10433 27022
rect -10365 26999 -10361 27015
rect -10360 26987 -10357 26995
rect -10301 26991 -10285 26993
rect -10238 26987 -10233 27022
rect -10050 27018 -10044 27033
rect -10151 27008 -10143 27018
rect -10050 27013 -10035 27018
rect -10141 27008 -10132 27011
rect -10141 26992 -10133 27008
rect -10132 26995 -10125 27008
rect -10050 27003 -10044 27013
rect -10020 26987 -10013 27033
rect -9928 27023 -9927 27033
rect -9958 26991 -9949 27001
rect -9948 26990 -9939 26991
rect -9876 26987 -9874 27046
rect -9868 27041 -9866 27046
rect -9848 27041 -9844 27056
rect -9840 27041 -9838 27071
rect -9828 27041 -9826 27082
rect -9823 27041 -9822 27071
rect -9862 27036 -9826 27041
rect -9792 27038 -9778 27046
rect -9862 27032 -9854 27036
rect -9848 27032 -9844 27036
rect -9862 27031 -9858 27032
rect -9852 27015 -9848 27031
rect -9850 27012 -9848 27015
rect -9842 27012 -9836 27020
rect -9850 27001 -9836 27012
rect -9828 27010 -9826 27036
rect -9742 27025 -9737 27055
rect -9732 27029 -9730 27304
rect -9718 27296 -9714 27304
rect -9708 27034 -9706 27304
rect -9674 27296 -9666 27304
rect -9626 27296 -9618 27304
rect -9732 27027 -9711 27029
rect -9735 27025 -9711 27027
rect -9732 27012 -9730 27025
rect -9832 26996 -9826 27010
rect -9744 27002 -9740 27012
rect -9732 27008 -9716 27012
rect -9710 27008 -9706 27034
rect -9679 27020 -9676 27047
rect -9674 27025 -9663 27047
rect -9661 27025 -9658 27055
rect -9679 27017 -9667 27020
rect -9732 27002 -9730 27008
rect -9828 26987 -9826 26996
rect -9746 26988 -9742 26998
rect -9734 26988 -9730 27002
rect -9733 26987 -9730 26988
rect -9708 26987 -9706 27008
rect -9612 27007 -9610 27304
rect -9598 27296 -9590 27304
rect -9550 27296 -9542 27304
rect -9593 27107 -9582 27111
rect -9581 27107 -9572 27279
rect -9581 27095 -9570 27107
rect -9581 27059 -9572 27095
rect -9516 27059 -9514 27304
rect -9502 27296 -9500 27304
rect -9488 27296 -9486 27304
rect -9474 27296 -9472 27304
rect -9505 27083 -9489 27091
rect -9608 27048 -9590 27059
rect -9583 27048 -9570 27059
rect -9523 27049 -9514 27059
rect -9512 27049 -9506 27079
rect -9505 27077 -9494 27079
rect -9505 27049 -9496 27070
rect -9590 27023 -9583 27047
rect -9598 27017 -9582 27023
rect -9612 26999 -9598 27007
rect -9612 26987 -9610 26999
rect -9590 26991 -9586 27017
rect -9516 27015 -9514 27049
rect -9513 27040 -9506 27049
rect -9494 27040 -9489 27070
rect -9513 27015 -9512 27040
rect -9480 27039 -9476 27049
rect -9468 27039 -9466 27304
rect -9460 27296 -9458 27304
rect -9446 27079 -9442 27081
rect -9448 27071 -9442 27079
rect -9447 27049 -9442 27051
rect -9436 27049 -9430 27071
rect -9420 27055 -9418 27317
rect -9396 27312 -9394 27317
rect -9372 27312 -9370 27317
rect -9406 27304 -9394 27312
rect -9378 27304 -9368 27312
rect -9346 27304 -9338 27312
rect -9318 27304 -9302 27312
rect -9412 27296 -9406 27304
rect -9396 27063 -9394 27304
rect -9384 27296 -9378 27304
rect -9372 27063 -9370 27304
rect -9338 27296 -9330 27304
rect -9401 27055 -9394 27063
rect -9516 26991 -9512 27015
rect -9506 27004 -9504 27014
rect -9494 27004 -9487 27015
rect -9470 27009 -9466 27039
rect -9516 26987 -9514 26991
rect -9513 26987 -9512 26991
rect -9496 26991 -9487 27004
rect -9482 26991 -9478 27004
rect -9496 26990 -9482 26991
rect -9494 26989 -9486 26990
rect -9468 26987 -9466 27009
rect -9420 27025 -9411 27055
rect -9406 27031 -9403 27041
rect -9396 27031 -9394 27055
rect -9391 27031 -9384 27055
rect -9374 27041 -9367 27063
rect -9396 27025 -9380 27031
rect -9372 27025 -9370 27041
rect -9420 27023 -9416 27025
rect -9420 26987 -9417 27023
rect -9396 27015 -9394 27025
rect -9374 27015 -9370 27025
rect -9343 27020 -9340 27047
rect -9338 27025 -9327 27047
rect -9325 27025 -9322 27055
rect -9343 27017 -9331 27020
rect -9408 27002 -9404 27012
rect -9398 27002 -9394 27015
rect -9391 27002 -9384 27015
rect -9398 27001 -9384 27002
rect -9398 26993 -9394 27001
rect -9398 26988 -9392 26993
rect -9391 26988 -9384 27001
rect -9400 26987 -9392 26988
rect -9372 26987 -9370 27015
rect -9300 26987 -9298 27317
rect -9252 27312 -9250 27317
rect -9156 27312 -9154 27317
rect -9132 27312 -9130 27317
rect -9286 27304 -9274 27312
rect -9258 27304 -9246 27312
rect -9226 27304 -9218 27312
rect -9164 27304 -9154 27312
rect -9136 27304 -9126 27312
rect -9290 27296 -9286 27304
rect -9262 27296 -9258 27304
rect -9262 27111 -9261 27279
rect -9252 27111 -9250 27304
rect -9218 27296 -9210 27304
rect -9170 27296 -9164 27304
rect -9262 27095 -9246 27111
rect -9262 27082 -9261 27095
rect -9272 27032 -9268 27056
rect -9264 27022 -9262 27047
rect -9252 27022 -9250 27095
rect -9219 27082 -9209 27104
rect -9168 27079 -9160 27090
rect -9156 27087 -9154 27304
rect -9142 27296 -9136 27304
rect -9176 27074 -9168 27079
rect -9166 27074 -9160 27079
rect -9158 27074 -9151 27087
rect -9136 27079 -9133 27092
rect -9166 27049 -9159 27074
rect -9156 27049 -9154 27074
rect -9247 27022 -9246 27047
rect -9216 27038 -9202 27046
rect -9158 27024 -9151 27049
rect -9144 27039 -9140 27049
rect -9132 27039 -9130 27304
rect -9110 27079 -9106 27081
rect -9112 27071 -9106 27079
rect -9111 27049 -9106 27051
rect -9100 27049 -9094 27071
rect -9084 27059 -9082 27317
rect -9060 27312 -9058 27317
rect -9036 27312 -9034 27317
rect -9068 27304 -9058 27312
rect -9040 27304 -9032 27312
rect -9008 27304 -8992 27312
rect -9076 27296 -9068 27304
rect -9091 27049 -9082 27059
rect -9080 27049 -9074 27079
rect -9060 27049 -9058 27304
rect -9048 27296 -9040 27304
rect -9055 27071 -9048 27079
rect -9036 27071 -9034 27304
rect -9026 27149 -9020 27279
rect -9026 27133 -9018 27149
rect -9036 27049 -9030 27071
rect -9026 27049 -9020 27133
rect -9000 27096 -8996 27106
rect -8988 27096 -8986 27317
rect -8964 27312 -8962 27317
rect -8940 27312 -8938 27317
rect -8976 27304 -8962 27312
rect -8948 27304 -8936 27312
rect -8916 27304 -8908 27312
rect -8980 27296 -8976 27304
rect -8990 27082 -8986 27096
rect -9014 27079 -9010 27081
rect -9016 27071 -9010 27079
rect -9004 27079 -8986 27082
rect -9004 27071 -8979 27079
rect -9015 27049 -9010 27051
rect -9004 27049 -8998 27071
rect -8990 27066 -8979 27071
rect -9264 27020 -9246 27022
rect -9266 27017 -9246 27020
rect -9286 27007 -9282 27017
rect -9276 27007 -9272 27012
rect -9266 27010 -9260 27017
rect -9252 27010 -9250 27017
rect -9276 26996 -9260 27007
rect -9256 26996 -9250 27010
rect -9177 27002 -9170 27014
rect -9156 27008 -9154 27024
rect -9136 27023 -9130 27039
rect -9134 27009 -9130 27023
rect -9276 26991 -9272 26996
rect -9274 26987 -9272 26991
rect -9252 26987 -9250 26996
rect -9158 26987 -9151 27008
rect -9132 26987 -9130 27009
rect -9084 26987 -9082 27049
rect -9081 27041 -9074 27049
rect -9062 27041 -9055 27049
rect -9050 27041 -9030 27049
rect -8988 27041 -8986 27066
rect -9081 27023 -9080 27041
rect -9060 26993 -9058 27041
rect -9050 27039 -9044 27041
rect -9036 27039 -9034 27041
rect -9040 27023 -9034 27039
rect -9038 27009 -9034 27023
rect -9060 26987 -9056 26993
rect -9036 26987 -9034 27009
rect -8991 27023 -8984 27041
rect -8972 27031 -8965 27066
rect -8964 27031 -8962 27304
rect -8952 27296 -8948 27304
rect -8959 27071 -8952 27079
rect -8940 27071 -8938 27304
rect -8908 27296 -8900 27304
rect -8892 27096 -8890 27317
rect -8888 27304 -8880 27312
rect -8880 27296 -8872 27304
rect -8896 27088 -8890 27096
rect -8959 27066 -8955 27071
rect -8945 27051 -8938 27071
rect -8914 27058 -8911 27088
rect -8892 27066 -8889 27088
rect -8869 27066 -8866 27096
rect -8844 27069 -8842 27317
rect -8796 27312 -8794 27317
rect -8700 27312 -8698 27317
rect -8604 27312 -8602 27317
rect -8556 27312 -8554 27317
rect -8826 27304 -8816 27312
rect -8798 27304 -8788 27312
rect -8766 27304 -8758 27312
rect -8738 27304 -8722 27312
rect -8706 27304 -8694 27312
rect -8678 27304 -8666 27312
rect -8646 27304 -8638 27312
rect -8618 27304 -8602 27312
rect -8588 27304 -8576 27312
rect -8560 27304 -8548 27312
rect -8832 27296 -8826 27304
rect -8804 27296 -8798 27304
rect -8816 27132 -8806 27134
rect -8806 27118 -8800 27132
rect -8796 27069 -8794 27304
rect -8758 27296 -8750 27304
rect -8710 27296 -8706 27304
rect -8906 27059 -8898 27066
rect -8892 27059 -8890 27066
rect -8889 27061 -8884 27066
rect -8889 27059 -8875 27061
rect -8906 27058 -8875 27059
rect -8855 27058 -8842 27069
rect -8835 27058 -8815 27069
rect -8808 27058 -8790 27069
rect -8906 27056 -8905 27058
rect -8904 27056 -8900 27058
rect -8892 27056 -8890 27058
rect -8945 27047 -8934 27051
rect -8950 27041 -8934 27047
rect -8959 27031 -8955 27041
rect -8991 26987 -8985 27023
rect -8972 27020 -8969 27031
rect -8976 27010 -8969 27020
rect -8964 27020 -8955 27031
rect -8964 27015 -8954 27020
rect -8972 26990 -8969 27010
rect -8966 27010 -8962 27015
rect -8959 27010 -8954 27015
rect -8945 27015 -8938 27041
rect -8896 27040 -8895 27056
rect -8894 27026 -8890 27056
rect -8966 27001 -8952 27010
rect -8966 26996 -8962 27001
rect -8959 26996 -8954 27001
rect -8980 26987 -8969 26990
rect -8964 26993 -8962 26996
rect -8964 26987 -8960 26993
rect -8945 26987 -8942 27015
rect -8940 26987 -8938 27015
rect -8892 27004 -8890 27026
rect -8905 26994 -8902 26998
rect -8905 26988 -8901 26994
rect -8896 26987 -8890 27004
rect -8844 27057 -8842 27058
rect -8844 27027 -8835 27057
rect -8830 27048 -8827 27057
rect -8815 27048 -8808 27058
rect -8820 27032 -8804 27048
rect -8818 27027 -8817 27032
rect -8816 27027 -8804 27032
rect -8844 26987 -8842 27027
rect -8815 26987 -8808 27027
rect -8796 26987 -8794 27058
rect -8767 27019 -8764 27049
rect -8762 27027 -8751 27049
rect -8749 27027 -8746 27057
rect -8740 27019 -8736 27027
rect -8756 26987 -8747 27019
rect -8700 26987 -8698 27304
rect -8682 27296 -8678 27304
rect -8638 27296 -8630 27304
rect -8695 27048 -8688 27057
rect -8680 27049 -8670 27064
rect -8604 27059 -8602 27304
rect -8590 27296 -8588 27304
rect -8576 27296 -8574 27304
rect -8562 27296 -8560 27304
rect -8593 27083 -8577 27091
rect -8686 27048 -8680 27049
rect -8678 27019 -8671 27049
rect -8669 27048 -8660 27059
rect -8611 27049 -8602 27059
rect -8600 27049 -8594 27079
rect -8593 27077 -8582 27079
rect -8593 27049 -8584 27070
rect -8680 26987 -8676 27019
rect -8604 27015 -8602 27049
rect -8601 27040 -8594 27049
rect -8582 27040 -8577 27070
rect -8601 27015 -8600 27040
rect -8568 27039 -8564 27049
rect -8556 27039 -8554 27304
rect -8548 27296 -8546 27304
rect -8534 27079 -8530 27081
rect -8536 27071 -8530 27079
rect -8535 27049 -8530 27051
rect -8524 27049 -8518 27071
rect -8508 27059 -8506 27317
rect -8484 27312 -8482 27317
rect -8460 27312 -8458 27317
rect -8492 27304 -8482 27312
rect -8464 27304 -8456 27312
rect -8500 27296 -8492 27304
rect -8515 27049 -8506 27059
rect -8504 27049 -8498 27079
rect -8484 27049 -8482 27304
rect -8472 27296 -8464 27304
rect -8479 27071 -8472 27079
rect -8460 27071 -8458 27304
rect -8450 27149 -8444 27279
rect -8450 27133 -8442 27149
rect -8460 27049 -8454 27071
rect -8450 27049 -8444 27133
rect -8438 27079 -8434 27081
rect -8440 27071 -8434 27079
rect -8439 27049 -8434 27051
rect -8428 27049 -8422 27071
rect -8412 27059 -8410 27317
rect -8388 27312 -8386 27317
rect -8364 27312 -8362 27317
rect -8396 27304 -8386 27312
rect -8368 27304 -8360 27312
rect -8404 27296 -8396 27304
rect -8419 27049 -8410 27059
rect -8408 27049 -8402 27079
rect -8388 27049 -8386 27304
rect -8376 27296 -8368 27304
rect -8383 27071 -8376 27079
rect -8364 27071 -8362 27304
rect -8354 27149 -8348 27279
rect -8354 27133 -8346 27149
rect -8364 27049 -8358 27071
rect -8354 27049 -8348 27133
rect -8342 27079 -8338 27081
rect -8344 27071 -8338 27079
rect -8343 27049 -8338 27051
rect -8332 27049 -8326 27071
rect -8316 27059 -8314 27317
rect -8292 27312 -8290 27317
rect -8268 27312 -8266 27317
rect -8196 27312 -8194 27317
rect -8300 27304 -8290 27312
rect -8272 27304 -8264 27312
rect -8202 27304 -8194 27312
rect -8174 27304 -8168 27312
rect -8142 27304 -8134 27312
rect -8114 27304 -8102 27312
rect -8100 27304 -8098 27317
rect -8052 27312 -8050 27317
rect -7932 27312 -7930 27317
rect -7836 27312 -7834 27317
rect -7740 27312 -7738 27317
rect -7692 27312 -7690 27317
rect -7620 27312 -7618 27317
rect -8086 27304 -8074 27312
rect -8058 27304 -8046 27312
rect -8026 27304 -8018 27312
rect -7962 27304 -7954 27312
rect -7934 27304 -7926 27312
rect -7902 27304 -7894 27312
rect -7874 27304 -7858 27312
rect -7842 27304 -7830 27312
rect -7814 27304 -7802 27312
rect -7782 27304 -7774 27312
rect -7754 27304 -7738 27312
rect -7724 27304 -7712 27312
rect -7696 27304 -7684 27312
rect -7626 27304 -7618 27312
rect -7598 27304 -7592 27312
rect -7566 27304 -7558 27312
rect -7538 27304 -7522 27312
rect -7506 27304 -7494 27312
rect -7478 27304 -7466 27312
rect -7446 27304 -7438 27312
rect -7390 27304 -7386 27309
rect -7362 27304 -7358 27309
rect -7356 27304 -7354 27317
rect -7284 27309 -7282 27317
rect -7212 27312 -7210 27317
rect -7188 27312 -7186 27317
rect -8308 27296 -8300 27304
rect -8323 27049 -8314 27059
rect -8312 27049 -8306 27079
rect -8292 27049 -8290 27304
rect -8280 27296 -8272 27304
rect -8287 27071 -8280 27079
rect -8268 27071 -8266 27304
rect -8212 27296 -8202 27304
rect -8258 27149 -8252 27279
rect -8258 27133 -8250 27149
rect -8268 27049 -8262 27071
rect -8258 27049 -8252 27133
rect -8246 27079 -8242 27081
rect -8248 27071 -8242 27079
rect -8247 27049 -8242 27051
rect -8236 27049 -8230 27071
rect -8604 26991 -8600 27015
rect -8594 27004 -8592 27014
rect -8582 27004 -8575 27015
rect -8558 27009 -8554 27039
rect -8604 26987 -8602 26991
rect -8601 26987 -8600 26991
rect -8584 26991 -8575 27004
rect -8570 26991 -8566 27004
rect -8584 26990 -8570 26991
rect -8582 26989 -8574 26990
rect -8556 26987 -8554 27009
rect -8508 26987 -8506 27049
rect -8505 27041 -8498 27049
rect -8486 27041 -8479 27049
rect -8474 27041 -8454 27049
rect -8505 27023 -8504 27041
rect -8484 26993 -8482 27041
rect -8474 27039 -8468 27041
rect -8460 27039 -8458 27041
rect -8464 27023 -8458 27039
rect -8462 27009 -8458 27023
rect -8484 26987 -8480 26993
rect -8460 26987 -8458 27009
rect -8412 26987 -8410 27049
rect -8409 27041 -8402 27049
rect -8390 27041 -8383 27049
rect -8378 27041 -8358 27049
rect -8409 27023 -8408 27041
rect -8388 26993 -8386 27041
rect -8378 27039 -8372 27041
rect -8364 27039 -8362 27041
rect -8368 27023 -8362 27039
rect -8366 27009 -8362 27023
rect -8388 26987 -8384 26993
rect -8364 26987 -8362 27009
rect -8316 26987 -8314 27049
rect -8313 27041 -8306 27049
rect -8294 27041 -8287 27049
rect -8282 27041 -8262 27049
rect -8313 27023 -8312 27041
rect -8292 26993 -8290 27041
rect -8282 27039 -8276 27041
rect -8268 27039 -8266 27041
rect -8272 27023 -8266 27039
rect -8270 27009 -8266 27023
rect -8292 26987 -8288 26993
rect -8268 26987 -8266 27009
rect -8196 27013 -8194 27304
rect -8184 27296 -8174 27304
rect -8134 27296 -8126 27304
rect -8102 27296 -8098 27304
rect -8074 27296 -8070 27304
rect -8191 27048 -8184 27078
rect -8182 27048 -8176 27071
rect -8174 27041 -8167 27071
rect -8165 27048 -8156 27279
rect -8100 27056 -8098 27296
rect -8089 27083 -8073 27099
rect -8095 27082 -8086 27083
rect -8102 27046 -8098 27056
rect -8182 27013 -8180 27023
rect -8174 27015 -8170 27041
rect -8100 27015 -8098 27046
rect -8092 27040 -8090 27046
rect -8089 27040 -8078 27046
rect -8074 27040 -8073 27070
rect -8072 27032 -8068 27040
rect -8196 27001 -8182 27013
rect -8172 27001 -8170 27013
rect -8196 26993 -8194 27001
rect -8196 26987 -8192 26993
rect -8100 26991 -8096 27015
rect -8090 27004 -8088 27014
rect -8072 27006 -8070 27012
rect -8066 27010 -8060 27020
rect -8052 27010 -8050 27304
rect -8046 27296 -8042 27304
rect -8018 27296 -8010 27304
rect -7970 27296 -7962 27304
rect -7942 27296 -7934 27304
rect -7952 27116 -7938 27132
rect -8019 27082 -8009 27104
rect -8016 27038 -8002 27046
rect -7966 27027 -7961 27057
rect -7952 27029 -7940 27038
rect -7932 27034 -7930 27304
rect -7894 27296 -7886 27304
rect -7846 27296 -7842 27304
rect -7954 27027 -7935 27029
rect -8076 27004 -8070 27006
rect -8100 26987 -8098 26991
rect -8080 26990 -8078 27004
rect -8072 26996 -8066 27004
rect -8056 26996 -8050 27010
rect -7979 27002 -7970 27014
rect -7934 27008 -7930 27034
rect -7903 27019 -7900 27049
rect -7898 27027 -7887 27049
rect -7885 27027 -7882 27057
rect -7876 27019 -7872 27027
rect -8052 26987 -8050 26996
rect -7932 26987 -7930 27008
rect -7892 26987 -7883 27019
rect -7836 26987 -7834 27304
rect -7818 27296 -7814 27304
rect -7774 27296 -7766 27304
rect -7831 27048 -7824 27057
rect -7816 27049 -7806 27064
rect -7740 27059 -7738 27304
rect -7726 27296 -7724 27304
rect -7712 27296 -7710 27304
rect -7698 27296 -7696 27304
rect -7729 27083 -7713 27091
rect -7822 27048 -7816 27049
rect -7814 27019 -7807 27049
rect -7805 27048 -7796 27059
rect -7747 27049 -7738 27059
rect -7736 27049 -7730 27079
rect -7729 27077 -7718 27079
rect -7729 27049 -7720 27070
rect -7816 26987 -7812 27019
rect -7740 27015 -7738 27049
rect -7737 27040 -7730 27049
rect -7718 27040 -7713 27070
rect -7737 27015 -7736 27040
rect -7704 27039 -7700 27049
rect -7692 27039 -7690 27304
rect -7684 27296 -7682 27304
rect -7636 27296 -7626 27304
rect -7670 27079 -7666 27081
rect -7672 27071 -7666 27079
rect -7671 27049 -7666 27051
rect -7660 27049 -7654 27071
rect -7740 26991 -7736 27015
rect -7730 27004 -7728 27014
rect -7718 27004 -7711 27015
rect -7694 27009 -7690 27039
rect -7740 26987 -7738 26991
rect -7737 26987 -7736 26991
rect -7720 26991 -7711 27004
rect -7706 26991 -7702 27004
rect -7720 26990 -7706 26991
rect -7718 26989 -7710 26990
rect -7692 26987 -7690 27009
rect -7620 27013 -7618 27304
rect -7608 27296 -7598 27304
rect -7558 27296 -7550 27304
rect -7510 27296 -7506 27304
rect -7482 27296 -7478 27304
rect -7438 27296 -7430 27304
rect -7386 27293 -7374 27304
rect -7358 27294 -7346 27304
rect -7310 27301 -7302 27309
rect -7284 27301 -7274 27309
rect -7254 27301 -7246 27309
rect -7226 27301 -7210 27312
rect -7196 27301 -7184 27312
rect -7168 27301 -7156 27312
rect -7302 27294 -7294 27301
rect -7362 27293 -7346 27294
rect -7310 27293 -7294 27294
rect -7284 27294 -7282 27301
rect -7274 27294 -7266 27301
rect -7246 27294 -7238 27301
rect -7284 27293 -7266 27294
rect -7254 27293 -7238 27294
rect -7226 27293 -7218 27294
rect -7615 27048 -7608 27078
rect -7606 27048 -7600 27071
rect -7598 27041 -7591 27071
rect -7589 27048 -7580 27279
rect -7381 27136 -7377 27146
rect -7398 27106 -7380 27111
rect -7371 27106 -7367 27136
rect -7508 27083 -7497 27090
rect -7380 27083 -7377 27099
rect -7506 27078 -7497 27083
rect -7496 27048 -7485 27078
rect -7606 27013 -7604 27023
rect -7598 27015 -7594 27041
rect -7496 27040 -7487 27048
rect -7396 27040 -7394 27080
rect -7380 27040 -7377 27070
rect -7496 27013 -7494 27015
rect -7620 27001 -7606 27013
rect -7596 27001 -7594 27013
rect -7504 27004 -7494 27013
rect -7380 27004 -7374 27015
rect -7620 26993 -7618 27001
rect -7500 26999 -7490 27004
rect -7380 26995 -7370 27004
rect -7620 26987 -7616 26993
rect -7496 26989 -7494 26990
rect -7380 26989 -7374 26995
rect -7356 26987 -7354 27293
rect -7334 27134 -7324 27140
rect -7332 27128 -7324 27134
rect -7284 27128 -7282 27293
rect -7264 27136 -7257 27146
rect -7264 27131 -7242 27136
rect -7322 27098 -7314 27128
rect -7304 27110 -7288 27126
rect -7295 27101 -7288 27110
rect -7284 27106 -7279 27128
rect -7264 27126 -7248 27131
rect -7284 27101 -7282 27106
rect -7310 27098 -7306 27101
rect -7295 27098 -7264 27101
rect -7320 27041 -7314 27098
rect -7295 27071 -7288 27098
rect -7304 27041 -7297 27071
rect -7284 27063 -7282 27098
rect -7246 27083 -7243 27091
rect -7236 27071 -7233 27083
rect -7273 27063 -7266 27071
rect -7291 27041 -7288 27063
rect -7295 27018 -7288 27041
rect -7284 27041 -7275 27063
rect -7273 27041 -7267 27063
rect -7284 27018 -7282 27041
rect -7295 27013 -7280 27018
rect -7295 27003 -7288 27013
rect -7284 26987 -7282 27013
rect -7265 26987 -7258 27063
rect -7256 27041 -7248 27063
rect -7246 27041 -7240 27071
rect -7212 26987 -7210 27301
rect -7198 27296 -7196 27301
rect -7208 27063 -7207 27079
rect -7192 27063 -7191 27065
rect -7190 27063 -7189 27065
rect -7188 27063 -7186 27301
rect -7184 27296 -7182 27301
rect -7170 27296 -7168 27301
rect -7156 27296 -7154 27301
rect -7154 27133 -7152 27140
rect -7142 27079 -7138 27081
rect -7183 27063 -7182 27079
rect -7144 27071 -7138 27079
rect -7207 27049 -7192 27063
rect -7190 27049 -7183 27063
rect -7163 27049 -7162 27065
rect -7143 27049 -7138 27051
rect -7132 27049 -7126 27071
rect -7116 27055 -7114 27317
rect -7092 27312 -7090 27317
rect -7068 27312 -7066 27317
rect -7102 27304 -7090 27312
rect -7074 27304 -7064 27312
rect -7042 27304 -7034 27312
rect -7108 27296 -7102 27304
rect -7092 27063 -7090 27304
rect -7080 27296 -7074 27304
rect -7068 27063 -7066 27304
rect -7034 27296 -7026 27304
rect -7097 27055 -7090 27063
rect -7190 27033 -7189 27049
rect -7198 26991 -7194 27001
rect -7188 26991 -7186 27049
rect -7168 27043 -7164 27049
rect -7168 27039 -7158 27043
rect -7168 27033 -7164 27039
rect -7116 27025 -7107 27055
rect -7102 27031 -7099 27041
rect -7092 27031 -7090 27055
rect -7087 27031 -7080 27055
rect -7070 27041 -7063 27063
rect -7092 27025 -7076 27031
rect -7068 27025 -7066 27041
rect -7116 27023 -7112 27025
rect -7188 26990 -7184 26991
rect -7188 26987 -7186 26990
rect -7116 26987 -7113 27023
rect -7092 27015 -7090 27025
rect -7070 27015 -7066 27025
rect -7039 27020 -7036 27047
rect -7034 27025 -7023 27047
rect -7021 27025 -7018 27055
rect -7039 27017 -7027 27020
rect -7104 27002 -7100 27012
rect -7094 27002 -7090 27015
rect -7087 27002 -7080 27015
rect -7094 27001 -7080 27002
rect -7094 26993 -7090 27001
rect -7094 26988 -7088 26993
rect -7087 26988 -7080 27001
rect -7096 26987 -7088 26988
rect -7068 26987 -7066 27015
rect -6996 26987 -6994 27317
rect -6972 27312 -6970 27317
rect -6948 27312 -6946 27317
rect -6980 27304 -6970 27312
rect -6952 27304 -6942 27312
rect -6986 27296 -6980 27304
rect -6992 27049 -6974 27059
rect -6972 27047 -6970 27304
rect -6958 27296 -6952 27304
rect -6948 27059 -6946 27304
rect -6967 27049 -6946 27059
rect -6938 27049 -6932 27279
rect -6926 27079 -6922 27081
rect -6928 27071 -6922 27079
rect -6927 27049 -6922 27051
rect -6916 27049 -6910 27071
rect -6900 27059 -6898 27317
rect -6876 27312 -6874 27317
rect -6852 27312 -6850 27317
rect -6884 27304 -6874 27312
rect -6856 27304 -6848 27312
rect -6892 27296 -6884 27304
rect -6907 27049 -6898 27059
rect -6896 27049 -6890 27079
rect -6876 27049 -6874 27304
rect -6864 27296 -6856 27304
rect -6871 27071 -6864 27079
rect -6852 27071 -6850 27304
rect -6842 27149 -6836 27279
rect -6842 27133 -6834 27149
rect -6852 27049 -6846 27071
rect -6842 27049 -6836 27133
rect -6830 27079 -6826 27081
rect -6832 27071 -6826 27079
rect -6831 27049 -6826 27051
rect -6820 27049 -6814 27071
rect -6804 27059 -6802 27317
rect -6780 27312 -6778 27317
rect -6756 27312 -6754 27317
rect -6788 27304 -6778 27312
rect -6760 27304 -6752 27312
rect -6796 27296 -6788 27304
rect -6811 27049 -6802 27059
rect -6800 27049 -6794 27079
rect -6780 27049 -6778 27304
rect -6768 27296 -6760 27304
rect -6775 27071 -6768 27079
rect -6756 27071 -6754 27304
rect -6746 27149 -6740 27279
rect -6746 27133 -6738 27149
rect -6756 27049 -6750 27071
rect -6746 27049 -6740 27133
rect -6734 27079 -6730 27081
rect -6736 27071 -6730 27079
rect -6735 27049 -6730 27051
rect -6724 27049 -6718 27071
rect -6708 27059 -6706 27317
rect -6684 27312 -6682 27317
rect -6660 27312 -6658 27317
rect -6692 27304 -6682 27312
rect -6664 27304 -6656 27312
rect -6700 27296 -6692 27304
rect -6715 27049 -6706 27059
rect -6704 27049 -6698 27079
rect -6684 27049 -6682 27304
rect -6672 27296 -6664 27304
rect -6679 27071 -6672 27079
rect -6660 27071 -6658 27304
rect -6650 27149 -6644 27279
rect -6650 27133 -6642 27149
rect -6660 27049 -6654 27071
rect -6650 27049 -6644 27133
rect -6638 27079 -6634 27081
rect -6640 27071 -6634 27079
rect -6639 27049 -6634 27051
rect -6628 27049 -6622 27071
rect -6612 27059 -6610 27317
rect -6588 27312 -6586 27317
rect -6564 27312 -6562 27317
rect -6596 27304 -6586 27312
rect -6568 27304 -6560 27312
rect -6604 27296 -6596 27304
rect -6619 27049 -6610 27059
rect -6608 27049 -6602 27079
rect -6588 27049 -6586 27304
rect -6576 27296 -6568 27304
rect -6583 27071 -6576 27079
rect -6564 27071 -6562 27304
rect -6554 27149 -6548 27279
rect -6554 27133 -6546 27149
rect -6564 27049 -6558 27071
rect -6554 27049 -6548 27133
rect -6542 27079 -6538 27081
rect -6544 27071 -6538 27079
rect -6543 27049 -6538 27051
rect -6532 27049 -6526 27071
rect -6516 27059 -6514 27317
rect -6492 27312 -6490 27317
rect -6468 27312 -6466 27317
rect -6500 27304 -6490 27312
rect -6472 27304 -6464 27312
rect -6508 27296 -6500 27304
rect -6523 27049 -6514 27059
rect -6512 27049 -6506 27079
rect -6492 27049 -6490 27304
rect -6480 27296 -6472 27304
rect -6487 27071 -6480 27079
rect -6468 27071 -6466 27304
rect -6458 27149 -6452 27279
rect -6458 27133 -6450 27149
rect -6468 27049 -6462 27071
rect -6458 27049 -6452 27133
rect -6446 27079 -6442 27081
rect -6448 27071 -6442 27079
rect -6447 27049 -6442 27051
rect -6436 27049 -6430 27071
rect -6420 27059 -6418 27317
rect -6396 27312 -6394 27317
rect -6372 27312 -6370 27317
rect -6404 27304 -6394 27312
rect -6376 27304 -6368 27312
rect -6412 27296 -6404 27304
rect -6427 27049 -6418 27059
rect -6416 27049 -6410 27079
rect -6396 27049 -6394 27304
rect -6384 27296 -6376 27304
rect -6391 27071 -6384 27079
rect -6372 27071 -6370 27304
rect -6362 27149 -6356 27279
rect -6362 27133 -6354 27149
rect -6372 27049 -6366 27071
rect -6362 27049 -6356 27133
rect -6350 27079 -6346 27081
rect -6352 27071 -6346 27079
rect -6351 27049 -6346 27051
rect -6340 27049 -6334 27071
rect -6324 27059 -6322 27317
rect -6300 27312 -6298 27317
rect -6276 27312 -6274 27317
rect -6308 27304 -6298 27312
rect -6280 27304 -6272 27312
rect -6316 27296 -6308 27304
rect -6331 27049 -6322 27059
rect -6320 27049 -6314 27079
rect -6300 27049 -6298 27304
rect -6288 27296 -6280 27304
rect -6295 27071 -6288 27079
rect -6276 27071 -6274 27304
rect -6266 27149 -6260 27279
rect -6266 27133 -6258 27149
rect -6276 27049 -6270 27071
rect -6266 27049 -6260 27133
rect -6254 27079 -6250 27081
rect -6256 27071 -6250 27079
rect -6255 27049 -6250 27051
rect -6244 27049 -6238 27071
rect -6228 27056 -6226 27317
rect -6180 27312 -6178 27317
rect -6060 27312 -6058 27317
rect -6214 27304 -6204 27312
rect -6186 27304 -6176 27312
rect -6154 27304 -6146 27312
rect -6126 27304 -6110 27312
rect -6094 27304 -6082 27312
rect -6066 27304 -6054 27312
rect -6034 27304 -6026 27312
rect -5978 27304 -5970 27309
rect -5964 27304 -5962 27317
rect -5950 27304 -5942 27309
rect -5940 27304 -5938 27317
rect -5868 27309 -5866 27317
rect -5796 27312 -5794 27317
rect -5652 27312 -5650 27317
rect -5316 27312 -5314 27317
rect -5268 27312 -5266 27317
rect -6220 27296 -6214 27304
rect -6192 27296 -6186 27304
rect -6223 27083 -6214 27084
rect -6204 27083 -6197 27084
rect -6190 27083 -6189 27279
rect -6180 27083 -6178 27304
rect -6146 27296 -6138 27304
rect -6098 27296 -6094 27304
rect -6070 27296 -6066 27304
rect -6082 27116 -6066 27124
rect -6223 27082 -6192 27083
rect -6190 27082 -6162 27083
rect -6147 27082 -6137 27104
rect -6103 27082 -6096 27104
rect -6094 27082 -6087 27112
rect -6082 27110 -6077 27112
rect -6070 27110 -6066 27112
rect -6085 27082 -6079 27104
rect -6974 27017 -6967 27047
rect -6960 27039 -6956 27049
rect -6948 27047 -6946 27049
rect -6948 27039 -6942 27047
rect -6952 27023 -6942 27039
rect -6950 27017 -6942 27023
rect -6972 26991 -6970 27017
rect -6950 27009 -6946 27017
rect -6972 26987 -6958 26991
rect -6948 26987 -6946 27009
rect -6900 26987 -6898 27049
rect -6897 27041 -6890 27049
rect -6878 27041 -6871 27049
rect -6866 27041 -6846 27049
rect -6897 27023 -6896 27041
rect -6876 26993 -6874 27041
rect -6866 27039 -6860 27041
rect -6852 27039 -6850 27041
rect -6856 27023 -6850 27039
rect -6854 27009 -6850 27023
rect -6876 26987 -6872 26993
rect -6852 26987 -6850 27009
rect -6804 26987 -6802 27049
rect -6801 27041 -6794 27049
rect -6782 27041 -6775 27049
rect -6770 27041 -6750 27049
rect -6801 27023 -6800 27041
rect -6780 26993 -6778 27041
rect -6770 27039 -6764 27041
rect -6756 27039 -6754 27041
rect -6760 27023 -6754 27039
rect -6758 27009 -6754 27023
rect -6780 26987 -6776 26993
rect -6756 26987 -6754 27009
rect -6708 26987 -6706 27049
rect -6705 27041 -6698 27049
rect -6686 27041 -6679 27049
rect -6674 27041 -6654 27049
rect -6705 27023 -6704 27041
rect -6684 26993 -6682 27041
rect -6674 27039 -6668 27041
rect -6660 27039 -6658 27041
rect -6664 27023 -6658 27039
rect -6662 27009 -6658 27023
rect -6684 26987 -6680 26993
rect -6660 26987 -6658 27009
rect -6612 26987 -6610 27049
rect -6609 27041 -6602 27049
rect -6590 27041 -6583 27049
rect -6578 27041 -6558 27049
rect -6609 27023 -6608 27041
rect -6588 26993 -6586 27041
rect -6578 27039 -6572 27041
rect -6564 27039 -6562 27041
rect -6568 27023 -6562 27039
rect -6566 27009 -6562 27023
rect -6588 26987 -6584 26993
rect -6564 26987 -6562 27009
rect -6516 26987 -6514 27049
rect -6513 27041 -6506 27049
rect -6494 27041 -6487 27049
rect -6482 27041 -6462 27049
rect -6513 27023 -6512 27041
rect -6492 26993 -6490 27041
rect -6482 27039 -6476 27041
rect -6468 27039 -6466 27041
rect -6472 27023 -6466 27039
rect -6470 27009 -6466 27023
rect -6492 26987 -6488 26993
rect -6468 26987 -6466 27009
rect -6420 26987 -6418 27049
rect -6417 27041 -6410 27049
rect -6398 27041 -6391 27049
rect -6386 27041 -6366 27049
rect -6417 27023 -6416 27041
rect -6396 26993 -6394 27041
rect -6386 27039 -6380 27041
rect -6372 27039 -6370 27041
rect -6376 27023 -6370 27039
rect -6374 27009 -6370 27023
rect -6396 26987 -6392 26993
rect -6372 26987 -6370 27009
rect -6324 26987 -6322 27049
rect -6321 27041 -6314 27049
rect -6302 27041 -6295 27049
rect -6290 27041 -6270 27049
rect -6230 27046 -6226 27056
rect -6321 27023 -6320 27041
rect -6300 26993 -6298 27041
rect -6290 27039 -6284 27041
rect -6276 27039 -6274 27041
rect -6280 27023 -6274 27039
rect -6278 27009 -6274 27023
rect -6300 26987 -6296 26993
rect -6276 26987 -6274 27009
rect -6228 26987 -6226 27046
rect -6220 27041 -6218 27046
rect -6200 27041 -6196 27056
rect -6192 27041 -6190 27071
rect -6180 27041 -6178 27082
rect -6077 27074 -6070 27104
rect -6068 27082 -6061 27104
rect -6175 27041 -6174 27071
rect -6110 27046 -6102 27056
rect -6214 27036 -6178 27041
rect -6144 27038 -6130 27046
rect -6100 27038 -6086 27046
rect -6080 27038 -6076 27056
rect -6214 27032 -6206 27036
rect -6200 27032 -6196 27036
rect -6214 27031 -6210 27032
rect -6204 27015 -6200 27031
rect -6202 27012 -6200 27015
rect -6194 27012 -6188 27020
rect -6202 27001 -6188 27012
rect -6180 27010 -6178 27036
rect -6100 27034 -6092 27038
rect -6100 27032 -6086 27034
rect -6082 27032 -6076 27038
rect -6100 27028 -6090 27032
rect -6094 27024 -6090 27028
rect -6082 27024 -6080 27032
rect -6184 26996 -6178 27010
rect -6100 27002 -6098 27014
rect -6084 27012 -6080 27024
rect -6068 27020 -6064 27024
rect -6074 27012 -6064 27020
rect -6084 27008 -6068 27012
rect -6060 27010 -6058 27304
rect -6026 27296 -6018 27304
rect -5970 27293 -5962 27304
rect -5942 27294 -5934 27304
rect -5894 27301 -5886 27309
rect -5868 27301 -5858 27309
rect -5838 27301 -5830 27309
rect -5810 27301 -5794 27312
rect -5778 27301 -5766 27312
rect -5750 27301 -5738 27312
rect -5718 27304 -5710 27312
rect -5690 27304 -5674 27312
rect -5658 27304 -5646 27312
rect -5630 27304 -5618 27312
rect -5598 27304 -5590 27312
rect -5570 27304 -5554 27312
rect -5538 27304 -5526 27312
rect -5510 27304 -5498 27312
rect -5478 27304 -5470 27312
rect -5450 27304 -5434 27312
rect -5418 27304 -5406 27312
rect -5390 27304 -5378 27312
rect -5358 27304 -5350 27312
rect -5330 27304 -5314 27312
rect -5300 27304 -5288 27312
rect -5272 27304 -5260 27312
rect -5886 27294 -5878 27301
rect -5950 27293 -5934 27294
rect -5894 27293 -5878 27294
rect -5868 27294 -5866 27301
rect -5858 27294 -5850 27301
rect -5830 27294 -5822 27301
rect -5868 27293 -5850 27294
rect -5838 27293 -5822 27294
rect -5810 27293 -5802 27294
rect -5964 27146 -5962 27293
rect -5965 27132 -5956 27146
rect -5965 27116 -5946 27132
rect -5940 27116 -5938 27293
rect -5918 27134 -5908 27140
rect -5916 27128 -5908 27134
rect -5868 27128 -5866 27293
rect -5848 27136 -5841 27146
rect -5848 27131 -5826 27136
rect -5982 27106 -5938 27116
rect -6027 27082 -6017 27104
rect -5965 27083 -5957 27106
rect -5965 27074 -5941 27083
rect -5980 27048 -5972 27074
rect -6024 27038 -6010 27046
rect -5980 27038 -5970 27048
rect -5980 27034 -5972 27038
rect -5980 27028 -5970 27034
rect -5974 27024 -5970 27028
rect -5964 27024 -5957 27074
rect -5951 27041 -5948 27048
rect -6080 26996 -6077 27008
rect -6064 26996 -6058 27010
rect -5980 27002 -5978 27014
rect -5964 27008 -5960 27024
rect -5948 27011 -5943 27024
rect -5959 27008 -5948 27011
rect -6180 26987 -6178 26996
rect -6060 26987 -6058 26996
rect -5964 26987 -5957 27008
rect -5940 26987 -5938 27106
rect -5906 27098 -5898 27128
rect -5888 27110 -5872 27126
rect -5879 27101 -5872 27110
rect -5868 27106 -5863 27128
rect -5848 27126 -5832 27131
rect -5868 27101 -5866 27106
rect -5894 27098 -5890 27101
rect -5879 27098 -5848 27101
rect -5904 27041 -5898 27098
rect -5879 27071 -5872 27098
rect -5888 27041 -5881 27071
rect -5868 27063 -5866 27098
rect -5830 27083 -5827 27091
rect -5820 27071 -5817 27083
rect -5857 27063 -5850 27071
rect -5875 27041 -5872 27063
rect -5879 27018 -5872 27041
rect -5868 27041 -5859 27063
rect -5857 27041 -5851 27063
rect -5868 27018 -5866 27041
rect -5879 27013 -5864 27018
rect -5879 27003 -5872 27013
rect -5868 26987 -5866 27013
rect -5849 26987 -5842 27063
rect -5840 27041 -5832 27063
rect -5830 27041 -5824 27071
rect -5796 27059 -5794 27301
rect -5782 27296 -5778 27301
rect -5754 27296 -5750 27301
rect -5710 27296 -5702 27304
rect -5662 27296 -5658 27304
rect -5768 27128 -5765 27138
rect -5768 27116 -5752 27128
rect -5768 27098 -5765 27116
rect -5797 27057 -5794 27059
rect -5777 27057 -5773 27063
rect -5796 27033 -5794 27057
rect -5791 27033 -5779 27057
rect -5777 27033 -5775 27057
rect -5773 27033 -5770 27057
rect -5768 27033 -5765 27073
rect -5764 27033 -5752 27057
rect -5750 27033 -5748 27063
rect -5796 27027 -5791 27033
rect -5770 27027 -5766 27033
rect -5796 26987 -5794 27027
rect -5719 27019 -5716 27049
rect -5714 27027 -5703 27049
rect -5701 27027 -5698 27057
rect -5692 27019 -5688 27027
rect -5708 26987 -5699 27019
rect -5652 26987 -5650 27304
rect -5634 27296 -5630 27304
rect -5590 27296 -5582 27304
rect -5542 27296 -5538 27304
rect -5514 27296 -5510 27304
rect -5470 27296 -5462 27304
rect -5422 27296 -5418 27304
rect -5394 27296 -5390 27304
rect -5350 27296 -5342 27304
rect -5540 27083 -5529 27090
rect -5420 27083 -5409 27090
rect -5538 27078 -5529 27083
rect -5418 27078 -5409 27083
rect -5647 27048 -5640 27057
rect -5632 27049 -5622 27064
rect -5638 27048 -5632 27049
rect -5630 27019 -5623 27049
rect -5621 27048 -5612 27059
rect -5528 27048 -5517 27078
rect -5408 27048 -5397 27078
rect -5316 27059 -5314 27304
rect -5302 27296 -5300 27304
rect -5288 27296 -5286 27304
rect -5274 27296 -5272 27304
rect -5305 27083 -5289 27091
rect -5323 27049 -5314 27059
rect -5312 27049 -5306 27079
rect -5305 27077 -5294 27079
rect -5305 27049 -5296 27070
rect -5528 27040 -5519 27048
rect -5408 27040 -5399 27048
rect -5632 26987 -5628 27019
rect -5316 27015 -5314 27049
rect -5313 27040 -5306 27049
rect -5294 27040 -5289 27070
rect -5313 27015 -5312 27040
rect -5280 27039 -5276 27049
rect -5268 27039 -5266 27304
rect -5260 27296 -5258 27304
rect -5246 27079 -5242 27081
rect -5248 27071 -5242 27079
rect -5247 27049 -5242 27051
rect -5236 27049 -5230 27071
rect -5220 27059 -5218 27317
rect -5196 27312 -5194 27317
rect -5172 27312 -5170 27317
rect -5204 27304 -5194 27312
rect -5176 27304 -5168 27312
rect -5212 27296 -5204 27304
rect -5227 27049 -5218 27059
rect -5216 27049 -5210 27079
rect -5196 27049 -5194 27304
rect -5184 27296 -5176 27304
rect -5191 27071 -5184 27079
rect -5172 27071 -5170 27304
rect -5162 27149 -5156 27279
rect -5162 27133 -5154 27149
rect -5172 27049 -5166 27071
rect -5162 27049 -5156 27133
rect -5150 27079 -5146 27081
rect -5152 27071 -5146 27079
rect -5151 27049 -5146 27051
rect -5140 27049 -5134 27071
rect -5124 27059 -5122 27317
rect -5100 27312 -5098 27317
rect -5076 27312 -5074 27317
rect -5108 27304 -5098 27312
rect -5080 27304 -5072 27312
rect -5116 27296 -5108 27304
rect -5131 27049 -5122 27059
rect -5120 27049 -5114 27079
rect -5100 27049 -5098 27304
rect -5088 27296 -5080 27304
rect -5095 27071 -5088 27079
rect -5076 27071 -5074 27304
rect -5066 27149 -5060 27279
rect -5066 27133 -5058 27149
rect -5076 27049 -5070 27071
rect -5066 27049 -5060 27133
rect -5054 27079 -5050 27081
rect -5056 27071 -5050 27079
rect -5055 27049 -5050 27051
rect -5044 27049 -5038 27071
rect -5028 27067 -5026 27317
rect -4980 27312 -4978 27317
rect -4884 27312 -4882 27317
rect -4860 27312 -4858 27317
rect -4788 27312 -4786 27317
rect -4692 27312 -4690 27317
rect -4644 27312 -4642 27317
rect -5010 27304 -5004 27312
rect -4982 27304 -4976 27312
rect -4950 27304 -4942 27312
rect -4922 27304 -4908 27312
rect -4892 27304 -4880 27312
rect -4864 27304 -4852 27312
rect -4794 27304 -4786 27312
rect -4766 27304 -4760 27312
rect -4734 27304 -4726 27312
rect -4706 27304 -4690 27312
rect -4676 27304 -4664 27312
rect -4648 27304 -4636 27312
rect -5020 27296 -5010 27304
rect -4992 27296 -4982 27304
rect -5000 27132 -4990 27141
rect -4990 27125 -4984 27132
rect -5037 27057 -5026 27067
rect -4980 27065 -4978 27304
rect -4942 27296 -4934 27304
rect -4908 27296 -4906 27304
rect -4894 27296 -4892 27304
rect -4914 27079 -4908 27089
rect -5009 27057 -5002 27065
rect -5528 27013 -5526 27015
rect -5408 27013 -5406 27015
rect -5536 27004 -5526 27013
rect -5416 27004 -5406 27013
rect -5532 26999 -5522 27004
rect -5412 26999 -5402 27004
rect -5316 26991 -5312 27015
rect -5306 27004 -5304 27014
rect -5294 27004 -5287 27015
rect -5270 27009 -5266 27039
rect -5528 26989 -5526 26990
rect -5408 26989 -5406 26990
rect -5316 26987 -5314 26991
rect -5313 26987 -5312 26991
rect -5296 26991 -5287 27004
rect -5282 26991 -5278 27004
rect -5296 26990 -5282 26991
rect -5294 26989 -5286 26990
rect -5268 26987 -5266 27009
rect -5220 26987 -5218 27049
rect -5217 27041 -5210 27049
rect -5198 27041 -5191 27049
rect -5186 27041 -5166 27049
rect -5217 27023 -5216 27041
rect -5196 26993 -5194 27041
rect -5186 27039 -5180 27041
rect -5172 27039 -5170 27041
rect -5176 27023 -5170 27039
rect -5174 27009 -5170 27023
rect -5196 26987 -5192 26993
rect -5172 26987 -5170 27009
rect -5124 26987 -5122 27049
rect -5121 27041 -5114 27049
rect -5102 27041 -5095 27049
rect -5090 27041 -5070 27049
rect -5028 27041 -5018 27057
rect -5121 27023 -5120 27041
rect -5100 26993 -5098 27041
rect -5090 27039 -5084 27041
rect -5076 27039 -5074 27041
rect -5080 27023 -5074 27039
rect -5078 27009 -5074 27023
rect -5100 26987 -5096 26993
rect -5076 26987 -5074 27009
rect -5028 27027 -5019 27041
rect -5014 27031 -5011 27041
rect -4999 27031 -4992 27057
rect -4990 27041 -4984 27057
rect -4982 27041 -4975 27065
rect -5004 27027 -4988 27031
rect -4980 27027 -4978 27041
rect -5028 27023 -5024 27027
rect -5028 26987 -5025 27023
rect -4982 27015 -4978 27027
rect -4951 27019 -4948 27049
rect -4946 27027 -4935 27049
rect -4933 27027 -4930 27057
rect -4915 27049 -4908 27059
rect -4904 27049 -4898 27079
rect -4884 27049 -4882 27304
rect -4880 27296 -4878 27304
rect -4866 27296 -4864 27304
rect -4879 27049 -4872 27057
rect -4860 27049 -4858 27304
rect -4852 27296 -4850 27304
rect -4804 27296 -4794 27304
rect -4838 27079 -4834 27081
rect -4840 27071 -4834 27079
rect -4850 27049 -4844 27059
rect -4839 27049 -4834 27051
rect -4828 27049 -4822 27071
rect -4924 27019 -4920 27027
rect -4905 27019 -4898 27049
rect -4886 27019 -4879 27049
rect -4872 27039 -4868 27049
rect -4860 27039 -4854 27049
rect -4864 27023 -4854 27039
rect -4862 27019 -4854 27023
rect -4999 26987 -4992 27015
rect -4980 26987 -4978 27015
rect -4940 26987 -4931 27019
rect -4884 26987 -4882 27019
rect -4862 27009 -4858 27019
rect -4860 27001 -4858 27009
rect -4864 26987 -4858 27001
rect -4788 27013 -4786 27304
rect -4776 27296 -4766 27304
rect -4726 27296 -4718 27304
rect -4783 27048 -4776 27078
rect -4774 27048 -4768 27071
rect -4766 27041 -4759 27071
rect -4757 27048 -4748 27279
rect -4692 27059 -4690 27304
rect -4678 27296 -4676 27304
rect -4664 27296 -4662 27304
rect -4650 27296 -4648 27304
rect -4681 27083 -4665 27091
rect -4699 27049 -4690 27059
rect -4688 27049 -4682 27079
rect -4681 27077 -4670 27079
rect -4681 27049 -4672 27070
rect -4774 27013 -4772 27023
rect -4766 27015 -4762 27041
rect -4692 27015 -4690 27049
rect -4689 27040 -4682 27049
rect -4670 27040 -4665 27070
rect -4689 27015 -4688 27040
rect -4656 27039 -4652 27049
rect -4644 27039 -4642 27304
rect -4636 27296 -4634 27304
rect -4622 27079 -4618 27081
rect -4624 27071 -4618 27079
rect -4623 27049 -4618 27051
rect -4612 27049 -4606 27071
rect -4596 27067 -4594 27317
rect -4548 27312 -4546 27317
rect -4428 27312 -4426 27317
rect -4332 27312 -4330 27317
rect -4308 27312 -4306 27317
rect -4578 27304 -4572 27312
rect -4550 27304 -4544 27312
rect -4518 27304 -4510 27312
rect -4490 27304 -4478 27312
rect -4462 27304 -4450 27312
rect -4434 27304 -4422 27312
rect -4402 27304 -4394 27312
rect -4340 27304 -4330 27312
rect -4312 27304 -4302 27312
rect -4588 27296 -4578 27304
rect -4560 27296 -4550 27304
rect -4568 27132 -4558 27141
rect -4558 27125 -4552 27132
rect -4605 27057 -4594 27067
rect -4548 27065 -4546 27304
rect -4510 27296 -4502 27304
rect -4478 27296 -4474 27304
rect -4450 27296 -4446 27304
rect -4483 27112 -4476 27124
rect -4477 27108 -4476 27112
rect -4471 27112 -4466 27279
rect -4471 27108 -4464 27112
rect -4471 27082 -4466 27108
rect -4577 27057 -4570 27065
rect -4788 27001 -4774 27013
rect -4764 27001 -4762 27013
rect -4788 26993 -4786 27001
rect -4788 26987 -4784 26993
rect -4692 26991 -4688 27015
rect -4682 27004 -4680 27014
rect -4670 27004 -4663 27015
rect -4646 27009 -4642 27039
rect -4692 26987 -4690 26991
rect -4689 26987 -4688 26991
rect -4672 26991 -4663 27004
rect -4658 26991 -4654 27004
rect -4672 26990 -4658 26991
rect -4670 26989 -4662 26990
rect -4644 26987 -4642 27009
rect -4596 27041 -4586 27057
rect -4596 27027 -4587 27041
rect -4582 27031 -4579 27041
rect -4567 27031 -4560 27057
rect -4558 27041 -4552 27057
rect -4550 27041 -4543 27065
rect -4572 27027 -4556 27031
rect -4548 27027 -4546 27041
rect -4596 27023 -4592 27027
rect -4596 26987 -4593 27023
rect -4550 27015 -4546 27027
rect -4519 27019 -4516 27049
rect -4514 27027 -4503 27049
rect -4501 27027 -4498 27057
rect -4478 27046 -4476 27056
rect -4492 27019 -4488 27027
rect -4468 27019 -4466 27046
rect -4448 27032 -4444 27056
rect -4440 27022 -4438 27049
rect -4440 27020 -4432 27022
rect -4442 27019 -4432 27020
rect -4567 26987 -4560 27015
rect -4548 26987 -4546 27015
rect -4508 26987 -4499 27019
rect -4442 27010 -4436 27019
rect -4428 27010 -4426 27304
rect -4422 27296 -4418 27304
rect -4394 27296 -4386 27304
rect -4346 27296 -4340 27304
rect -4395 27082 -4385 27104
rect -4344 27079 -4336 27090
rect -4332 27087 -4330 27304
rect -4318 27296 -4312 27304
rect -4352 27074 -4344 27079
rect -4342 27074 -4336 27079
rect -4334 27074 -4327 27087
rect -4312 27079 -4309 27092
rect -4342 27049 -4335 27074
rect -4332 27049 -4330 27074
rect -4423 27019 -4422 27049
rect -4392 27038 -4378 27046
rect -4334 27024 -4327 27049
rect -4320 27039 -4316 27049
rect -4308 27039 -4306 27304
rect -4286 27079 -4282 27081
rect -4288 27071 -4282 27079
rect -4287 27049 -4282 27051
rect -4276 27049 -4270 27071
rect -4260 27067 -4258 27317
rect -4212 27312 -4210 27317
rect -4116 27312 -4114 27317
rect -4092 27312 -4090 27317
rect -4020 27312 -4018 27317
rect -4242 27304 -4236 27312
rect -4214 27304 -4208 27312
rect -4182 27304 -4174 27312
rect -4154 27304 -4140 27312
rect -4124 27304 -4112 27312
rect -4096 27304 -4084 27312
rect -4026 27304 -4018 27312
rect -3998 27304 -3992 27312
rect -3966 27304 -3958 27312
rect -3910 27304 -3906 27309
rect -3882 27304 -3878 27309
rect -3876 27304 -3874 27317
rect -3804 27309 -3802 27317
rect -3732 27312 -3730 27317
rect -3588 27312 -3586 27317
rect -3564 27312 -3562 27317
rect -4252 27296 -4242 27304
rect -4224 27296 -4214 27304
rect -4232 27132 -4222 27141
rect -4222 27125 -4216 27132
rect -4269 27057 -4258 27067
rect -4212 27065 -4210 27304
rect -4174 27296 -4166 27304
rect -4140 27296 -4138 27304
rect -4126 27296 -4124 27304
rect -4146 27079 -4140 27089
rect -4241 27057 -4234 27065
rect -4432 26996 -4426 27010
rect -4353 27002 -4346 27014
rect -4332 27008 -4330 27024
rect -4312 27023 -4306 27039
rect -4310 27009 -4306 27023
rect -4428 26987 -4426 26996
rect -4334 26987 -4327 27008
rect -4308 26987 -4306 27009
rect -4260 27041 -4250 27057
rect -4260 27027 -4251 27041
rect -4246 27031 -4243 27041
rect -4231 27031 -4224 27057
rect -4222 27041 -4216 27057
rect -4214 27041 -4207 27065
rect -4236 27027 -4220 27031
rect -4212 27027 -4210 27041
rect -4260 27023 -4256 27027
rect -4260 26987 -4257 27023
rect -4214 27015 -4210 27027
rect -4183 27019 -4180 27049
rect -4178 27027 -4167 27049
rect -4165 27027 -4162 27057
rect -4147 27049 -4140 27059
rect -4136 27049 -4130 27079
rect -4116 27049 -4114 27304
rect -4112 27296 -4110 27304
rect -4098 27296 -4096 27304
rect -4111 27049 -4104 27057
rect -4092 27049 -4090 27304
rect -4084 27296 -4082 27304
rect -4036 27296 -4026 27304
rect -4070 27079 -4066 27081
rect -4072 27071 -4066 27079
rect -4082 27049 -4076 27059
rect -4071 27049 -4066 27051
rect -4060 27049 -4054 27071
rect -4156 27019 -4152 27027
rect -4137 27019 -4130 27049
rect -4118 27019 -4111 27049
rect -4104 27039 -4100 27049
rect -4092 27039 -4086 27049
rect -4096 27023 -4086 27039
rect -4094 27019 -4086 27023
rect -4231 26987 -4224 27015
rect -4212 26987 -4210 27015
rect -4172 26987 -4163 27019
rect -4116 26987 -4114 27019
rect -4094 27009 -4090 27019
rect -4092 27001 -4090 27009
rect -4096 26987 -4090 27001
rect -4020 27013 -4018 27304
rect -4008 27296 -3998 27304
rect -3958 27296 -3950 27304
rect -3906 27293 -3894 27304
rect -3878 27294 -3866 27304
rect -3830 27301 -3822 27309
rect -3804 27301 -3794 27309
rect -3774 27301 -3766 27309
rect -3746 27301 -3730 27312
rect -3714 27301 -3702 27312
rect -3686 27301 -3674 27312
rect -3654 27304 -3646 27312
rect -3626 27304 -3612 27312
rect -3596 27304 -3584 27312
rect -3568 27304 -3556 27312
rect -3822 27294 -3814 27301
rect -3882 27293 -3866 27294
rect -3830 27293 -3814 27294
rect -3804 27294 -3802 27301
rect -3794 27294 -3786 27301
rect -3766 27294 -3758 27301
rect -3804 27293 -3786 27294
rect -3774 27293 -3758 27294
rect -3746 27293 -3738 27294
rect -4015 27048 -4008 27078
rect -4006 27048 -4000 27071
rect -3998 27041 -3991 27071
rect -3989 27048 -3980 27279
rect -3901 27136 -3897 27146
rect -3918 27106 -3900 27111
rect -3891 27106 -3887 27136
rect -3900 27083 -3897 27099
rect -4006 27013 -4004 27023
rect -3998 27015 -3994 27041
rect -3916 27040 -3914 27080
rect -3900 27040 -3897 27070
rect -4020 27001 -4006 27013
rect -3996 27001 -3994 27013
rect -3900 27004 -3894 27015
rect -4020 26993 -4018 27001
rect -3900 26995 -3890 27004
rect -4020 26987 -4016 26993
rect -3900 26989 -3894 26995
rect -3876 26987 -3874 27293
rect -3854 27134 -3844 27140
rect -3852 27128 -3844 27134
rect -3804 27128 -3802 27293
rect -3784 27136 -3777 27146
rect -3784 27131 -3762 27136
rect -3842 27098 -3834 27128
rect -3824 27110 -3808 27126
rect -3815 27101 -3808 27110
rect -3804 27106 -3799 27128
rect -3784 27126 -3768 27131
rect -3804 27101 -3802 27106
rect -3830 27098 -3826 27101
rect -3815 27098 -3784 27101
rect -3840 27041 -3834 27098
rect -3815 27071 -3808 27098
rect -3824 27041 -3817 27071
rect -3804 27063 -3802 27098
rect -3766 27083 -3763 27091
rect -3756 27071 -3753 27083
rect -3793 27063 -3786 27071
rect -3811 27041 -3808 27063
rect -3815 27018 -3808 27041
rect -3804 27041 -3795 27063
rect -3793 27041 -3787 27063
rect -3804 27018 -3802 27041
rect -3815 27013 -3800 27018
rect -3815 27003 -3808 27013
rect -3804 26987 -3802 27013
rect -3785 26987 -3778 27063
rect -3776 27041 -3768 27063
rect -3766 27041 -3760 27071
rect -3732 27059 -3730 27301
rect -3718 27296 -3714 27301
rect -3690 27296 -3686 27301
rect -3646 27296 -3638 27304
rect -3612 27296 -3610 27304
rect -3598 27296 -3596 27304
rect -3704 27128 -3701 27138
rect -3704 27116 -3688 27128
rect -3704 27098 -3701 27116
rect -3618 27079 -3612 27089
rect -3733 27057 -3730 27059
rect -3713 27057 -3709 27063
rect -3732 27033 -3730 27057
rect -3727 27033 -3715 27057
rect -3713 27033 -3711 27057
rect -3709 27033 -3706 27057
rect -3704 27033 -3701 27073
rect -3700 27033 -3688 27057
rect -3686 27033 -3684 27063
rect -3732 27027 -3727 27033
rect -3706 27027 -3702 27033
rect -3732 26987 -3730 27027
rect -3655 27019 -3652 27049
rect -3650 27027 -3639 27049
rect -3637 27027 -3634 27057
rect -3619 27049 -3612 27059
rect -3608 27049 -3602 27079
rect -3588 27049 -3586 27304
rect -3584 27296 -3582 27304
rect -3570 27296 -3568 27304
rect -3583 27049 -3576 27057
rect -3564 27049 -3562 27304
rect -3556 27296 -3554 27304
rect -3542 27079 -3538 27081
rect -3544 27071 -3538 27079
rect -3554 27049 -3548 27059
rect -3543 27049 -3538 27051
rect -3532 27049 -3526 27071
rect -3516 27059 -3514 27317
rect -3492 27312 -3490 27317
rect -3468 27312 -3466 27317
rect -3500 27304 -3490 27312
rect -3472 27304 -3464 27312
rect -3508 27296 -3500 27304
rect -3523 27049 -3514 27059
rect -3512 27049 -3506 27079
rect -3492 27049 -3490 27304
rect -3480 27296 -3472 27304
rect -3487 27071 -3480 27079
rect -3468 27071 -3466 27304
rect -3458 27149 -3452 27279
rect -3458 27133 -3450 27149
rect -3468 27049 -3462 27071
rect -3458 27049 -3452 27133
rect -3446 27079 -3442 27081
rect -3448 27071 -3442 27079
rect -3447 27049 -3442 27051
rect -3436 27049 -3430 27071
rect -3420 27056 -3418 27317
rect -3372 27312 -3370 27317
rect -3252 27312 -3250 27317
rect -3156 27312 -3154 27317
rect -3132 27312 -3130 27317
rect -3406 27304 -3396 27312
rect -3378 27304 -3368 27312
rect -3346 27304 -3338 27312
rect -3318 27304 -3302 27312
rect -3286 27304 -3274 27312
rect -3258 27304 -3246 27312
rect -3226 27304 -3218 27312
rect -3198 27304 -3182 27312
rect -3166 27304 -3154 27312
rect -3138 27304 -3126 27312
rect -3106 27304 -3098 27312
rect -3412 27296 -3406 27304
rect -3384 27296 -3378 27304
rect -3415 27083 -3406 27084
rect -3396 27083 -3389 27084
rect -3382 27083 -3381 27279
rect -3372 27083 -3370 27304
rect -3338 27296 -3330 27304
rect -3290 27296 -3286 27304
rect -3262 27296 -3258 27304
rect -3274 27116 -3258 27124
rect -3415 27082 -3384 27083
rect -3382 27082 -3354 27083
rect -3339 27082 -3329 27104
rect -3295 27082 -3288 27104
rect -3286 27082 -3279 27112
rect -3274 27110 -3269 27112
rect -3262 27110 -3258 27112
rect -3277 27082 -3271 27104
rect -3628 27019 -3624 27027
rect -3609 27019 -3602 27049
rect -3590 27019 -3583 27049
rect -3576 27039 -3572 27049
rect -3564 27039 -3558 27049
rect -3568 27023 -3558 27039
rect -3566 27019 -3558 27023
rect -3644 26987 -3635 27019
rect -3588 26987 -3586 27019
rect -3566 27009 -3562 27019
rect -3564 27001 -3562 27009
rect -3568 26987 -3562 27001
rect -3516 26987 -3514 27049
rect -3513 27041 -3506 27049
rect -3494 27041 -3487 27049
rect -3482 27041 -3462 27049
rect -3422 27046 -3418 27056
rect -3513 27023 -3512 27041
rect -3492 26993 -3490 27041
rect -3482 27039 -3476 27041
rect -3468 27039 -3466 27041
rect -3472 27023 -3466 27039
rect -3470 27009 -3466 27023
rect -3492 26987 -3488 26993
rect -3468 26987 -3466 27009
rect -3420 26987 -3418 27046
rect -3412 27041 -3410 27046
rect -3392 27041 -3388 27056
rect -3384 27041 -3382 27071
rect -3372 27041 -3370 27082
rect -3269 27074 -3262 27104
rect -3260 27082 -3253 27104
rect -3367 27041 -3366 27071
rect -3302 27046 -3294 27056
rect -3406 27036 -3370 27041
rect -3336 27038 -3322 27046
rect -3292 27038 -3278 27046
rect -3272 27038 -3268 27056
rect -3406 27032 -3398 27036
rect -3392 27032 -3388 27036
rect -3406 27031 -3402 27032
rect -3396 27015 -3392 27031
rect -3394 27012 -3392 27015
rect -3386 27012 -3380 27020
rect -3394 27001 -3380 27012
rect -3372 27010 -3370 27036
rect -3292 27034 -3284 27038
rect -3292 27032 -3278 27034
rect -3274 27032 -3268 27038
rect -3292 27028 -3282 27032
rect -3286 27024 -3282 27028
rect -3274 27024 -3272 27032
rect -3376 26996 -3370 27010
rect -3292 27002 -3290 27014
rect -3276 27012 -3272 27024
rect -3260 27020 -3256 27024
rect -3266 27012 -3256 27020
rect -3276 27008 -3260 27012
rect -3252 27010 -3250 27304
rect -3218 27296 -3210 27304
rect -3170 27296 -3166 27304
rect -3219 27082 -3209 27104
rect -3216 27038 -3202 27046
rect -3166 27025 -3161 27055
rect -3156 27029 -3154 27304
rect -3142 27296 -3138 27304
rect -3132 27034 -3130 27304
rect -3098 27296 -3090 27304
rect -3060 27055 -3058 27317
rect -3012 27312 -3010 27317
rect -2916 27312 -2914 27317
rect -2892 27312 -2890 27317
rect -3042 27304 -3034 27312
rect -3014 27304 -3006 27312
rect -2982 27304 -2974 27312
rect -2954 27304 -2940 27312
rect -2924 27304 -2912 27312
rect -2896 27304 -2884 27312
rect -3050 27296 -3042 27304
rect -3022 27296 -3014 27304
rect -3032 27116 -3016 27123
rect -3156 27027 -3135 27029
rect -3159 27025 -3135 27027
rect -3156 27012 -3154 27025
rect -3272 26996 -3269 27008
rect -3256 26996 -3250 27010
rect -3168 27002 -3164 27012
rect -3156 27008 -3140 27012
rect -3134 27008 -3130 27034
rect -3103 27020 -3100 27047
rect -3098 27025 -3087 27047
rect -3085 27025 -3082 27055
rect -3060 27027 -3051 27055
rect -3031 27027 -3024 27055
rect -3012 27047 -3010 27304
rect -2974 27296 -2966 27304
rect -2940 27296 -2938 27304
rect -2926 27296 -2924 27304
rect -2946 27079 -2940 27089
rect -3022 27027 -3016 27047
rect -3103 27017 -3091 27020
rect -3156 27002 -3154 27008
rect -3372 26987 -3370 26996
rect -3252 26987 -3250 26996
rect -3170 26988 -3166 26998
rect -3158 26988 -3154 27002
rect -3157 26987 -3154 26988
rect -3132 26987 -3130 27008
rect -3060 26987 -3058 27027
rect -3041 27017 -3034 27027
rect -3014 27017 -3007 27047
rect -2983 27019 -2980 27049
rect -2978 27027 -2967 27049
rect -2965 27027 -2962 27057
rect -2947 27049 -2940 27059
rect -2936 27049 -2930 27079
rect -2916 27049 -2914 27304
rect -2912 27296 -2910 27304
rect -2898 27296 -2896 27304
rect -2911 27049 -2904 27057
rect -2892 27049 -2890 27304
rect -2884 27296 -2882 27304
rect -2870 27079 -2866 27081
rect -2872 27071 -2866 27079
rect -2882 27049 -2876 27059
rect -2871 27049 -2866 27051
rect -2860 27049 -2854 27071
rect -2844 27059 -2842 27317
rect -2820 27312 -2818 27317
rect -2796 27312 -2794 27317
rect -2828 27304 -2818 27312
rect -2800 27304 -2792 27312
rect -2836 27296 -2828 27304
rect -2851 27049 -2842 27059
rect -2840 27049 -2834 27079
rect -2820 27049 -2818 27304
rect -2808 27296 -2800 27304
rect -2815 27071 -2808 27079
rect -2796 27071 -2794 27304
rect -2786 27149 -2780 27279
rect -2786 27133 -2778 27149
rect -2796 27049 -2790 27071
rect -2786 27049 -2780 27133
rect -2774 27079 -2770 27081
rect -2776 27071 -2770 27079
rect -2775 27049 -2770 27051
rect -2764 27049 -2758 27071
rect -2748 27067 -2746 27317
rect -2700 27312 -2698 27317
rect -2604 27312 -2602 27317
rect -2580 27312 -2578 27317
rect -2508 27312 -2506 27317
rect -2730 27304 -2724 27312
rect -2702 27304 -2696 27312
rect -2670 27304 -2662 27312
rect -2642 27304 -2628 27312
rect -2612 27304 -2600 27312
rect -2584 27304 -2572 27312
rect -2514 27304 -2506 27312
rect -2486 27304 -2480 27312
rect -2454 27304 -2446 27312
rect -2426 27304 -2414 27312
rect -2412 27304 -2410 27317
rect -2364 27312 -2362 27317
rect -2398 27304 -2386 27312
rect -2370 27304 -2358 27312
rect -2338 27304 -2330 27312
rect -2740 27296 -2730 27304
rect -2712 27296 -2702 27304
rect -2720 27132 -2710 27141
rect -2710 27125 -2704 27132
rect -2757 27057 -2746 27067
rect -2700 27065 -2698 27304
rect -2662 27296 -2654 27304
rect -2628 27296 -2626 27304
rect -2614 27296 -2612 27304
rect -2634 27079 -2628 27089
rect -2729 27057 -2722 27065
rect -2956 27019 -2952 27027
rect -2937 27019 -2930 27049
rect -2918 27019 -2911 27049
rect -2904 27039 -2900 27049
rect -2892 27039 -2886 27049
rect -2896 27023 -2886 27039
rect -2894 27019 -2886 27023
rect -3031 27007 -3024 27017
rect -3014 26991 -3010 27017
rect -3031 26987 -3024 26991
rect -3012 26987 -3010 26991
rect -2972 26987 -2963 27019
rect -2916 26987 -2914 27019
rect -2894 27009 -2890 27019
rect -2892 27001 -2890 27009
rect -2896 26987 -2890 27001
rect -2844 26987 -2842 27049
rect -2841 27041 -2834 27049
rect -2822 27041 -2815 27049
rect -2810 27041 -2790 27049
rect -2748 27041 -2738 27057
rect -2841 27023 -2840 27041
rect -2820 26993 -2818 27041
rect -2810 27039 -2804 27041
rect -2796 27039 -2794 27041
rect -2800 27023 -2794 27039
rect -2798 27009 -2794 27023
rect -2820 26987 -2816 26993
rect -2796 26987 -2794 27009
rect -2748 27027 -2739 27041
rect -2734 27031 -2731 27041
rect -2719 27031 -2712 27057
rect -2710 27041 -2704 27057
rect -2702 27041 -2695 27065
rect -2724 27027 -2708 27031
rect -2700 27027 -2698 27041
rect -2748 27023 -2744 27027
rect -2748 26987 -2745 27023
rect -2702 27015 -2698 27027
rect -2671 27019 -2668 27049
rect -2666 27027 -2655 27049
rect -2653 27027 -2650 27057
rect -2635 27049 -2628 27059
rect -2624 27049 -2618 27079
rect -2604 27049 -2602 27304
rect -2600 27296 -2598 27304
rect -2586 27296 -2584 27304
rect -2599 27049 -2592 27057
rect -2580 27049 -2578 27304
rect -2572 27296 -2570 27304
rect -2524 27296 -2514 27304
rect -2558 27079 -2554 27081
rect -2560 27071 -2554 27079
rect -2570 27049 -2564 27059
rect -2559 27049 -2554 27051
rect -2548 27049 -2542 27071
rect -2644 27019 -2640 27027
rect -2625 27019 -2618 27049
rect -2606 27019 -2599 27049
rect -2592 27039 -2588 27049
rect -2580 27039 -2574 27049
rect -2584 27023 -2574 27039
rect -2582 27019 -2574 27023
rect -2719 26987 -2712 27015
rect -2700 26987 -2698 27015
rect -2660 26987 -2651 27019
rect -2604 26987 -2602 27019
rect -2582 27009 -2578 27019
rect -2580 27001 -2578 27009
rect -2584 26987 -2578 27001
rect -2508 27013 -2506 27304
rect -2496 27296 -2486 27304
rect -2446 27296 -2438 27304
rect -2414 27296 -2410 27304
rect -2386 27296 -2382 27304
rect -2503 27048 -2496 27078
rect -2494 27048 -2488 27071
rect -2486 27041 -2479 27071
rect -2477 27048 -2468 27279
rect -2412 27056 -2410 27296
rect -2412 27055 -2401 27056
rect -2494 27013 -2492 27023
rect -2486 27015 -2482 27041
rect -2412 27025 -2403 27055
rect -2401 27040 -2395 27055
rect -2393 27040 -2386 27063
rect -2508 27001 -2494 27013
rect -2484 27001 -2482 27013
rect -2508 26993 -2506 27001
rect -2508 26987 -2504 26993
rect -2412 26987 -2408 27025
rect -2402 27004 -2400 27014
rect -2392 27002 -2390 27004
rect -2378 27002 -2376 27004
rect -2392 26998 -2378 27002
rect -2402 26990 -2378 26998
rect -2402 26989 -2392 26990
rect -2390 26989 -2382 26990
rect -2364 26987 -2362 27304
rect -2358 27296 -2354 27304
rect -2330 27296 -2322 27304
rect -2335 27020 -2332 27047
rect -2330 27025 -2319 27047
rect -2317 27025 -2314 27055
rect -2335 27017 -2323 27020
rect -2292 26987 -2290 27317
rect -2268 27312 -2266 27317
rect -2244 27312 -2242 27317
rect -2276 27304 -2266 27312
rect -2248 27304 -2238 27312
rect -2282 27296 -2276 27304
rect -2288 27049 -2270 27059
rect -2268 27047 -2266 27304
rect -2254 27296 -2248 27304
rect -2244 27059 -2242 27304
rect -2263 27049 -2242 27059
rect -2234 27049 -2228 27279
rect -2222 27079 -2218 27081
rect -2224 27071 -2218 27079
rect -2223 27049 -2218 27051
rect -2212 27049 -2206 27071
rect -2196 27059 -2194 27317
rect -2172 27312 -2170 27317
rect -2148 27312 -2146 27317
rect -2180 27304 -2170 27312
rect -2152 27304 -2144 27312
rect -2188 27296 -2180 27304
rect -2203 27049 -2194 27059
rect -2192 27049 -2186 27079
rect -2172 27049 -2170 27304
rect -2160 27296 -2152 27304
rect -2167 27071 -2160 27079
rect -2148 27071 -2146 27304
rect -2138 27149 -2132 27279
rect -2138 27133 -2130 27149
rect -2148 27049 -2142 27071
rect -2138 27049 -2132 27133
rect -2126 27079 -2122 27081
rect -2128 27071 -2122 27079
rect -2127 27049 -2122 27051
rect -2116 27049 -2110 27071
rect -2100 27059 -2098 27317
rect -2076 27312 -2074 27317
rect -2052 27312 -2050 27317
rect -1980 27312 -1978 27317
rect -2084 27304 -2074 27312
rect -2056 27304 -2048 27312
rect -1986 27304 -1978 27312
rect -1958 27304 -1952 27312
rect -1926 27304 -1918 27312
rect -1898 27304 -1886 27312
rect -1884 27304 -1882 27317
rect -1836 27312 -1834 27317
rect -1716 27312 -1714 27317
rect -1596 27312 -1594 27317
rect -1476 27312 -1474 27317
rect -1380 27312 -1378 27317
rect -1356 27312 -1354 27317
rect -1870 27304 -1858 27312
rect -1842 27304 -1830 27312
rect -1810 27304 -1802 27312
rect -1782 27304 -1766 27312
rect -1750 27304 -1738 27312
rect -1722 27304 -1710 27312
rect -1690 27304 -1682 27312
rect -1662 27304 -1646 27312
rect -1630 27304 -1618 27312
rect -1602 27304 -1590 27312
rect -1570 27304 -1562 27312
rect -1542 27304 -1526 27312
rect -1510 27304 -1498 27312
rect -1482 27304 -1470 27312
rect -1450 27304 -1442 27312
rect -1388 27304 -1378 27312
rect -1360 27304 -1350 27312
rect -2092 27296 -2084 27304
rect -2107 27049 -2098 27059
rect -2096 27049 -2090 27079
rect -2076 27049 -2074 27304
rect -2064 27296 -2056 27304
rect -2071 27071 -2064 27079
rect -2052 27071 -2050 27304
rect -1996 27296 -1986 27304
rect -2042 27149 -2036 27279
rect -2042 27133 -2034 27149
rect -2052 27049 -2046 27071
rect -2042 27049 -2036 27133
rect -2030 27079 -2026 27081
rect -2032 27071 -2026 27079
rect -2031 27049 -2026 27051
rect -2020 27049 -2014 27071
rect -2270 27017 -2263 27047
rect -2256 27039 -2252 27049
rect -2244 27047 -2242 27049
rect -2244 27039 -2238 27047
rect -2248 27023 -2238 27039
rect -2246 27017 -2238 27023
rect -2268 26991 -2266 27017
rect -2246 27009 -2242 27017
rect -2268 26987 -2254 26991
rect -2244 26987 -2242 27009
rect -2196 26987 -2194 27049
rect -2193 27041 -2186 27049
rect -2174 27041 -2167 27049
rect -2162 27041 -2142 27049
rect -2193 27023 -2192 27041
rect -2172 26993 -2170 27041
rect -2162 27039 -2156 27041
rect -2148 27039 -2146 27041
rect -2152 27023 -2146 27039
rect -2150 27009 -2146 27023
rect -2172 26987 -2168 26993
rect -2148 26987 -2146 27009
rect -2100 26987 -2098 27049
rect -2097 27041 -2090 27049
rect -2078 27041 -2071 27049
rect -2066 27041 -2046 27049
rect -2097 27023 -2096 27041
rect -2076 26993 -2074 27041
rect -2066 27039 -2060 27041
rect -2052 27039 -2050 27041
rect -2056 27023 -2050 27039
rect -2054 27009 -2050 27023
rect -2076 26987 -2072 26993
rect -2052 26987 -2050 27009
rect -1980 27013 -1978 27304
rect -1968 27296 -1958 27304
rect -1918 27296 -1910 27304
rect -1886 27296 -1882 27304
rect -1858 27296 -1854 27304
rect -1975 27048 -1968 27078
rect -1966 27048 -1960 27071
rect -1958 27041 -1951 27071
rect -1949 27048 -1940 27279
rect -1884 27056 -1882 27296
rect -1873 27083 -1857 27099
rect -1879 27082 -1870 27083
rect -1886 27046 -1882 27056
rect -1966 27013 -1964 27023
rect -1958 27015 -1954 27041
rect -1884 27015 -1882 27046
rect -1876 27040 -1874 27046
rect -1873 27040 -1862 27046
rect -1858 27040 -1857 27070
rect -1856 27032 -1852 27040
rect -1980 27001 -1966 27013
rect -1956 27001 -1954 27013
rect -1980 26993 -1978 27001
rect -1980 26987 -1976 26993
rect -1884 26991 -1880 27015
rect -1874 27004 -1872 27014
rect -1856 27006 -1854 27012
rect -1850 27010 -1844 27020
rect -1836 27010 -1834 27304
rect -1830 27296 -1826 27304
rect -1802 27296 -1794 27304
rect -1754 27296 -1750 27304
rect -1726 27296 -1722 27304
rect -1738 27116 -1722 27124
rect -1803 27082 -1793 27104
rect -1759 27082 -1752 27104
rect -1750 27082 -1743 27112
rect -1738 27110 -1733 27112
rect -1726 27110 -1722 27112
rect -1741 27082 -1735 27104
rect -1733 27074 -1726 27104
rect -1724 27082 -1717 27104
rect -1766 27046 -1758 27056
rect -1800 27038 -1786 27046
rect -1756 27038 -1742 27046
rect -1736 27038 -1732 27056
rect -1756 27034 -1748 27038
rect -1756 27032 -1742 27034
rect -1738 27032 -1732 27038
rect -1756 27028 -1746 27032
rect -1750 27024 -1746 27028
rect -1738 27024 -1736 27032
rect -1860 27004 -1854 27006
rect -1884 26987 -1882 26991
rect -1864 26990 -1862 27004
rect -1856 26996 -1850 27004
rect -1840 26996 -1834 27010
rect -1756 27002 -1754 27014
rect -1740 27012 -1736 27024
rect -1724 27020 -1720 27024
rect -1730 27012 -1720 27020
rect -1740 27008 -1724 27012
rect -1716 27010 -1714 27304
rect -1682 27296 -1674 27304
rect -1634 27296 -1630 27304
rect -1606 27296 -1602 27304
rect -1618 27116 -1602 27124
rect -1683 27082 -1673 27104
rect -1639 27082 -1632 27104
rect -1630 27082 -1623 27112
rect -1618 27110 -1613 27112
rect -1606 27110 -1602 27112
rect -1621 27082 -1615 27104
rect -1613 27074 -1606 27104
rect -1604 27082 -1597 27104
rect -1646 27046 -1638 27056
rect -1680 27038 -1666 27046
rect -1636 27038 -1622 27046
rect -1616 27038 -1612 27056
rect -1636 27034 -1628 27038
rect -1636 27032 -1622 27034
rect -1618 27032 -1612 27038
rect -1636 27028 -1626 27032
rect -1630 27024 -1626 27028
rect -1618 27024 -1616 27032
rect -1736 26996 -1733 27008
rect -1720 26996 -1714 27010
rect -1636 27002 -1634 27014
rect -1620 27012 -1616 27024
rect -1604 27020 -1600 27024
rect -1610 27012 -1600 27020
rect -1620 27008 -1604 27012
rect -1596 27010 -1594 27304
rect -1562 27296 -1554 27304
rect -1514 27296 -1510 27304
rect -1486 27296 -1482 27304
rect -1498 27116 -1482 27124
rect -1563 27082 -1553 27104
rect -1519 27082 -1512 27104
rect -1510 27082 -1503 27112
rect -1498 27110 -1493 27112
rect -1486 27110 -1482 27112
rect -1501 27082 -1495 27104
rect -1493 27074 -1486 27104
rect -1484 27082 -1477 27104
rect -1526 27046 -1518 27056
rect -1560 27038 -1546 27046
rect -1516 27038 -1502 27046
rect -1496 27038 -1492 27056
rect -1516 27034 -1508 27038
rect -1516 27032 -1502 27034
rect -1498 27032 -1492 27038
rect -1516 27028 -1506 27032
rect -1510 27024 -1506 27028
rect -1498 27024 -1496 27032
rect -1616 26996 -1613 27008
rect -1600 26996 -1594 27010
rect -1516 27002 -1514 27014
rect -1500 27012 -1496 27024
rect -1484 27020 -1480 27024
rect -1490 27012 -1480 27020
rect -1500 27008 -1484 27012
rect -1476 27010 -1474 27304
rect -1442 27296 -1434 27304
rect -1394 27296 -1388 27304
rect -1443 27082 -1433 27104
rect -1392 27079 -1384 27090
rect -1380 27087 -1378 27304
rect -1366 27296 -1360 27304
rect -1400 27074 -1392 27079
rect -1390 27074 -1384 27079
rect -1382 27074 -1375 27087
rect -1360 27079 -1357 27092
rect -1390 27049 -1383 27074
rect -1380 27049 -1378 27074
rect -1440 27038 -1426 27046
rect -1382 27024 -1375 27049
rect -1368 27039 -1364 27049
rect -1356 27039 -1354 27304
rect -1334 27079 -1330 27081
rect -1336 27071 -1330 27079
rect -1335 27049 -1330 27051
rect -1324 27049 -1318 27071
rect -1308 27056 -1306 27317
rect -1260 27312 -1258 27317
rect -1164 27312 -1162 27317
rect -1140 27312 -1138 27317
rect -1068 27312 -1066 27317
rect -852 27312 -850 27317
rect -804 27312 -802 27317
rect -1294 27304 -1284 27312
rect -1266 27304 -1256 27312
rect -1234 27304 -1226 27312
rect -1172 27304 -1162 27312
rect -1144 27304 -1134 27312
rect -1074 27304 -1066 27312
rect -1046 27304 -1040 27312
rect -1014 27304 -1006 27312
rect -986 27304 -970 27312
rect -954 27304 -942 27312
rect -926 27304 -914 27312
rect -894 27304 -886 27312
rect -866 27304 -850 27312
rect -836 27304 -824 27312
rect -808 27304 -796 27312
rect -1300 27296 -1294 27304
rect -1272 27296 -1266 27304
rect -1303 27083 -1294 27084
rect -1284 27083 -1277 27084
rect -1270 27083 -1269 27279
rect -1260 27083 -1258 27304
rect -1226 27296 -1218 27304
rect -1178 27296 -1172 27304
rect -1303 27082 -1272 27083
rect -1270 27082 -1242 27083
rect -1227 27082 -1217 27104
rect -1310 27046 -1306 27056
rect -1496 26996 -1493 27008
rect -1480 26996 -1474 27010
rect -1401 27002 -1394 27014
rect -1380 27008 -1378 27024
rect -1360 27023 -1354 27039
rect -1358 27009 -1354 27023
rect -1836 26987 -1834 26996
rect -1716 26987 -1714 26996
rect -1596 26987 -1594 26996
rect -1476 26987 -1474 26996
rect -1382 26987 -1375 27008
rect -1356 26987 -1354 27009
rect -1308 26987 -1306 27046
rect -1300 27041 -1298 27046
rect -1280 27041 -1276 27056
rect -1272 27041 -1270 27071
rect -1260 27041 -1258 27082
rect -1176 27079 -1168 27090
rect -1164 27087 -1162 27304
rect -1150 27296 -1144 27304
rect -1184 27074 -1176 27079
rect -1174 27074 -1168 27079
rect -1166 27074 -1159 27087
rect -1144 27079 -1141 27092
rect -1255 27041 -1254 27071
rect -1174 27049 -1167 27074
rect -1164 27049 -1162 27074
rect -1294 27036 -1258 27041
rect -1224 27038 -1210 27046
rect -1294 27032 -1286 27036
rect -1280 27032 -1276 27036
rect -1294 27031 -1290 27032
rect -1284 27015 -1280 27031
rect -1282 27012 -1280 27015
rect -1274 27012 -1268 27020
rect -1282 27001 -1268 27012
rect -1260 27010 -1258 27036
rect -1166 27024 -1159 27049
rect -1152 27039 -1148 27049
rect -1140 27039 -1138 27304
rect -1084 27296 -1074 27304
rect -1118 27079 -1114 27081
rect -1120 27071 -1114 27079
rect -1119 27049 -1114 27051
rect -1108 27049 -1102 27071
rect -1264 26996 -1258 27010
rect -1185 27002 -1178 27014
rect -1164 27008 -1162 27024
rect -1144 27023 -1138 27039
rect -1142 27009 -1138 27023
rect -1260 26987 -1258 26996
rect -1166 26987 -1159 27008
rect -1140 26987 -1138 27009
rect -1068 27013 -1066 27304
rect -1056 27296 -1046 27304
rect -1006 27296 -998 27304
rect -958 27296 -954 27304
rect -930 27296 -926 27304
rect -886 27296 -878 27304
rect -1063 27048 -1056 27078
rect -1054 27048 -1048 27071
rect -1046 27041 -1039 27071
rect -1037 27048 -1028 27279
rect -956 27083 -945 27090
rect -954 27078 -945 27083
rect -944 27048 -933 27078
rect -852 27059 -850 27304
rect -838 27296 -836 27304
rect -824 27296 -822 27304
rect -810 27296 -808 27304
rect -841 27083 -825 27091
rect -859 27049 -850 27059
rect -848 27049 -842 27079
rect -841 27077 -830 27079
rect -841 27049 -832 27070
rect -1054 27013 -1052 27023
rect -1046 27015 -1042 27041
rect -944 27040 -935 27048
rect -852 27015 -850 27049
rect -849 27040 -842 27049
rect -830 27040 -825 27070
rect -849 27015 -848 27040
rect -816 27039 -812 27049
rect -804 27039 -802 27304
rect -796 27296 -794 27304
rect -782 27079 -778 27081
rect -784 27071 -778 27079
rect -783 27049 -778 27051
rect -772 27049 -766 27071
rect -756 27067 -754 27317
rect -708 27312 -706 27317
rect -612 27312 -610 27317
rect -588 27312 -586 27317
rect -738 27304 -732 27312
rect -710 27304 -704 27312
rect -678 27304 -670 27312
rect -650 27304 -636 27312
rect -620 27304 -608 27312
rect -592 27304 -580 27312
rect -748 27296 -738 27304
rect -720 27296 -710 27304
rect -728 27132 -718 27141
rect -718 27125 -712 27132
rect -765 27057 -754 27067
rect -708 27065 -706 27304
rect -670 27296 -662 27304
rect -636 27296 -634 27304
rect -622 27296 -620 27304
rect -642 27079 -636 27089
rect -737 27057 -730 27065
rect -944 27013 -942 27015
rect -1068 27001 -1054 27013
rect -1044 27001 -1042 27013
rect -952 27004 -942 27013
rect -1068 26993 -1066 27001
rect -948 26999 -938 27004
rect -1068 26987 -1064 26993
rect -852 26991 -848 27015
rect -842 27004 -840 27014
rect -830 27004 -823 27015
rect -806 27009 -802 27039
rect -944 26989 -942 26990
rect -852 26987 -850 26991
rect -849 26987 -848 26991
rect -832 26991 -823 27004
rect -818 26991 -814 27004
rect -832 26990 -818 26991
rect -830 26989 -822 26990
rect -804 26987 -802 27009
rect -756 27041 -746 27057
rect -756 27027 -747 27041
rect -742 27031 -739 27041
rect -727 27031 -720 27057
rect -718 27041 -712 27057
rect -710 27041 -703 27065
rect -732 27027 -716 27031
rect -708 27027 -706 27041
rect -756 27023 -752 27027
rect -756 26987 -753 27023
rect -710 27015 -706 27027
rect -679 27019 -676 27049
rect -674 27027 -663 27049
rect -661 27027 -658 27057
rect -643 27049 -636 27059
rect -632 27049 -626 27079
rect -612 27049 -610 27304
rect -608 27296 -606 27304
rect -594 27296 -592 27304
rect -607 27049 -600 27057
rect -588 27049 -586 27304
rect -580 27296 -578 27304
rect -566 27079 -562 27081
rect -568 27071 -562 27079
rect -578 27049 -572 27059
rect -567 27049 -562 27051
rect -556 27049 -550 27071
rect -540 27059 -538 27317
rect -516 27312 -514 27317
rect -492 27312 -490 27317
rect -524 27304 -514 27312
rect -496 27304 -488 27312
rect -532 27296 -524 27304
rect -547 27049 -538 27059
rect -536 27049 -530 27079
rect -516 27049 -514 27304
rect -504 27296 -496 27304
rect -511 27071 -504 27079
rect -492 27071 -490 27304
rect -482 27149 -476 27279
rect -482 27133 -474 27149
rect -492 27049 -486 27071
rect -482 27049 -476 27133
rect -470 27079 -466 27081
rect -472 27071 -466 27079
rect -471 27049 -466 27051
rect -460 27049 -454 27071
rect -444 27067 -442 27317
rect -396 27312 -394 27317
rect -300 27312 -298 27317
rect -276 27312 -274 27317
rect -204 27312 -202 27317
rect -108 27312 -106 27317
rect -60 27312 -58 27317
rect 12 27312 14 27317
rect 108 27312 110 27317
rect 156 27312 158 27317
rect -426 27304 -420 27312
rect -398 27304 -392 27312
rect -366 27304 -358 27312
rect -338 27304 -324 27312
rect -308 27304 -296 27312
rect -280 27304 -268 27312
rect -210 27304 -202 27312
rect -182 27304 -176 27312
rect -150 27304 -142 27312
rect -122 27304 -106 27312
rect -92 27304 -80 27312
rect -64 27304 -52 27312
rect 6 27304 14 27312
rect 34 27304 40 27312
rect 66 27304 74 27312
rect 94 27304 110 27312
rect 124 27304 136 27312
rect 152 27304 164 27312
rect -436 27296 -426 27304
rect -408 27296 -398 27304
rect -416 27132 -406 27141
rect -406 27125 -400 27132
rect -453 27057 -442 27067
rect -396 27065 -394 27304
rect -358 27296 -350 27304
rect -324 27296 -322 27304
rect -310 27296 -308 27304
rect -330 27079 -324 27089
rect -425 27057 -418 27065
rect -652 27019 -648 27027
rect -633 27019 -626 27049
rect -614 27019 -607 27049
rect -600 27039 -596 27049
rect -588 27039 -582 27049
rect -592 27023 -582 27039
rect -590 27019 -582 27023
rect -727 26987 -720 27015
rect -708 26987 -706 27015
rect -668 26987 -659 27019
rect -612 26987 -610 27019
rect -590 27009 -586 27019
rect -588 27001 -586 27009
rect -592 26987 -586 27001
rect -540 26987 -538 27049
rect -537 27041 -530 27049
rect -518 27041 -511 27049
rect -506 27041 -486 27049
rect -444 27041 -434 27057
rect -537 27023 -536 27041
rect -516 26993 -514 27041
rect -506 27039 -500 27041
rect -492 27039 -490 27041
rect -496 27023 -490 27039
rect -494 27009 -490 27023
rect -516 26987 -512 26993
rect -492 26987 -490 27009
rect -444 27027 -435 27041
rect -430 27031 -427 27041
rect -415 27031 -408 27057
rect -406 27041 -400 27057
rect -398 27041 -391 27065
rect -420 27027 -404 27031
rect -396 27027 -394 27041
rect -444 27023 -440 27027
rect -444 26987 -441 27023
rect -398 27015 -394 27027
rect -367 27019 -364 27049
rect -362 27027 -351 27049
rect -349 27027 -346 27057
rect -331 27049 -324 27059
rect -320 27049 -314 27079
rect -300 27049 -298 27304
rect -296 27296 -294 27304
rect -282 27296 -280 27304
rect -295 27049 -288 27057
rect -276 27049 -274 27304
rect -268 27296 -266 27304
rect -220 27296 -210 27304
rect -254 27079 -250 27081
rect -256 27071 -250 27079
rect -266 27049 -260 27059
rect -255 27049 -250 27051
rect -244 27049 -238 27071
rect -340 27019 -336 27027
rect -321 27019 -314 27049
rect -302 27019 -295 27049
rect -288 27039 -284 27049
rect -276 27039 -270 27049
rect -280 27023 -270 27039
rect -278 27019 -270 27023
rect -415 26987 -408 27015
rect -396 26987 -394 27015
rect -356 26987 -347 27019
rect -300 26987 -298 27019
rect -278 27009 -274 27019
rect -276 27001 -274 27009
rect -280 26987 -274 27001
rect -204 27013 -202 27304
rect -192 27296 -182 27304
rect -142 27296 -134 27304
rect -199 27048 -192 27078
rect -190 27048 -184 27071
rect -182 27041 -175 27071
rect -173 27048 -164 27279
rect -108 27059 -106 27304
rect -94 27296 -92 27304
rect -80 27296 -78 27304
rect -66 27296 -64 27304
rect -97 27083 -81 27091
rect -115 27049 -106 27059
rect -104 27049 -98 27079
rect -97 27077 -86 27079
rect -97 27049 -88 27070
rect -190 27013 -188 27023
rect -182 27015 -178 27041
rect -108 27015 -106 27049
rect -105 27040 -98 27049
rect -86 27040 -81 27070
rect -105 27015 -104 27040
rect -72 27039 -68 27049
rect -60 27039 -58 27304
rect -52 27296 -50 27304
rect -4 27296 6 27304
rect -38 27079 -34 27081
rect -40 27071 -34 27079
rect -39 27049 -34 27051
rect -28 27049 -22 27071
rect -204 27001 -190 27013
rect -180 27001 -178 27013
rect -204 26993 -202 27001
rect -204 26987 -200 26993
rect -108 26991 -104 27015
rect -98 27004 -96 27014
rect -86 27004 -79 27015
rect -62 27009 -58 27039
rect -108 26987 -106 26991
rect -105 26987 -104 26991
rect -88 26991 -79 27004
rect -74 26991 -70 27004
rect -88 26990 -74 26991
rect -86 26989 -78 26990
rect -60 26987 -58 27009
rect 12 27013 14 27304
rect 24 27296 34 27304
rect 74 27296 82 27304
rect 17 27048 24 27078
rect 26 27048 32 27071
rect 34 27041 41 27071
rect 43 27048 52 27279
rect 108 27059 110 27304
rect 122 27296 124 27304
rect 136 27296 138 27304
rect 150 27296 152 27304
rect 119 27083 135 27091
rect 101 27049 110 27059
rect 112 27049 118 27079
rect 119 27077 130 27079
rect 119 27049 128 27070
rect 26 27013 28 27023
rect 34 27015 38 27041
rect 108 27015 110 27049
rect 111 27040 118 27049
rect 130 27040 135 27070
rect 111 27015 112 27040
rect 144 27039 148 27049
rect 156 27039 158 27304
rect 164 27296 166 27304
rect 178 27079 182 27081
rect 176 27071 182 27079
rect 177 27049 182 27051
rect 188 27049 194 27071
rect 204 27059 206 27317
rect 228 27312 230 27317
rect 252 27312 254 27317
rect 220 27304 230 27312
rect 248 27304 256 27312
rect 212 27296 220 27304
rect 197 27049 206 27059
rect 208 27049 214 27079
rect 228 27049 230 27304
rect 240 27296 248 27304
rect 233 27071 240 27079
rect 252 27071 254 27304
rect 262 27149 268 27279
rect 262 27133 270 27149
rect 252 27049 258 27071
rect 262 27049 268 27133
rect 274 27079 278 27081
rect 272 27071 278 27079
rect 273 27049 278 27051
rect 284 27049 290 27071
rect 300 27056 302 27317
rect 348 27312 350 27317
rect 468 27312 470 27317
rect 564 27312 566 27317
rect 588 27312 590 27317
rect 314 27304 324 27312
rect 342 27304 352 27312
rect 374 27304 382 27312
rect 402 27304 418 27312
rect 434 27304 446 27312
rect 462 27304 474 27312
rect 494 27304 502 27312
rect 556 27304 566 27312
rect 584 27304 594 27312
rect 308 27296 314 27304
rect 336 27296 342 27304
rect 305 27083 314 27084
rect 324 27083 331 27084
rect 338 27083 339 27279
rect 348 27083 350 27304
rect 382 27296 390 27304
rect 430 27296 434 27304
rect 458 27296 462 27304
rect 446 27116 462 27124
rect 305 27082 336 27083
rect 338 27082 366 27083
rect 381 27082 391 27104
rect 425 27082 432 27104
rect 434 27082 441 27112
rect 446 27110 451 27112
rect 458 27110 462 27112
rect 443 27082 449 27104
rect 12 27001 26 27013
rect 36 27001 38 27013
rect 12 26993 14 27001
rect 12 26987 16 26993
rect 108 26991 112 27015
rect 118 27004 120 27014
rect 130 27004 137 27015
rect 154 27009 158 27039
rect 108 26987 110 26991
rect 111 26987 112 26991
rect 128 26991 137 27004
rect 142 26991 146 27004
rect 128 26990 142 26991
rect 130 26989 138 26990
rect 156 26987 158 27009
rect 204 26987 206 27049
rect 207 27041 214 27049
rect 226 27041 233 27049
rect 238 27041 258 27049
rect 298 27046 302 27056
rect 207 27023 208 27041
rect 228 26993 230 27041
rect 238 27039 244 27041
rect 252 27039 254 27041
rect 248 27023 254 27039
rect 250 27009 254 27023
rect 228 26987 232 26993
rect 252 26987 254 27009
rect 300 26987 302 27046
rect 308 27041 310 27046
rect 328 27041 332 27056
rect 336 27041 338 27071
rect 348 27041 350 27082
rect 451 27074 458 27104
rect 460 27082 467 27104
rect 353 27041 354 27071
rect 418 27046 426 27056
rect 314 27036 350 27041
rect 384 27038 398 27046
rect 428 27038 442 27046
rect 448 27038 452 27056
rect 314 27032 322 27036
rect 328 27032 332 27036
rect 314 27031 318 27032
rect 324 27015 328 27031
rect 326 27012 328 27015
rect 334 27012 340 27020
rect 326 27001 340 27012
rect 348 27010 350 27036
rect 428 27034 436 27038
rect 428 27032 442 27034
rect 446 27032 452 27038
rect 428 27028 438 27032
rect 434 27024 438 27028
rect 446 27024 448 27032
rect 344 26996 350 27010
rect 428 27002 430 27014
rect 444 27012 448 27024
rect 460 27020 464 27024
rect 454 27012 464 27020
rect 444 27008 460 27012
rect 468 27010 470 27304
rect 502 27296 510 27304
rect 550 27296 556 27304
rect 501 27082 511 27104
rect 552 27079 560 27090
rect 564 27087 566 27304
rect 578 27296 584 27304
rect 544 27074 552 27079
rect 554 27074 560 27079
rect 562 27074 569 27087
rect 584 27079 587 27092
rect 554 27049 561 27074
rect 564 27049 566 27074
rect 504 27038 518 27046
rect 562 27024 569 27049
rect 576 27039 580 27049
rect 588 27039 590 27304
rect 610 27079 614 27081
rect 608 27071 614 27079
rect 609 27049 614 27051
rect 620 27049 626 27071
rect 636 27059 638 27317
rect 660 27312 662 27317
rect 684 27312 686 27317
rect 652 27304 662 27312
rect 680 27304 688 27312
rect 644 27296 652 27304
rect 629 27049 638 27059
rect 640 27049 646 27079
rect 660 27049 662 27304
rect 672 27296 680 27304
rect 665 27071 672 27079
rect 684 27071 686 27304
rect 694 27149 700 27279
rect 694 27133 702 27149
rect 684 27049 690 27071
rect 694 27049 700 27133
rect 706 27079 710 27081
rect 704 27071 710 27079
rect 705 27049 710 27051
rect 716 27049 722 27071
rect 732 27055 734 27317
rect 756 27312 758 27317
rect 780 27312 782 27317
rect 876 27312 878 27317
rect 972 27312 974 27317
rect 1020 27312 1022 27317
rect 746 27304 758 27312
rect 774 27304 784 27312
rect 806 27304 814 27312
rect 870 27304 878 27312
rect 898 27304 906 27312
rect 930 27304 938 27312
rect 958 27304 974 27312
rect 988 27304 1000 27312
rect 1016 27304 1028 27312
rect 740 27296 746 27304
rect 756 27063 758 27304
rect 768 27296 774 27304
rect 780 27063 782 27304
rect 814 27296 822 27304
rect 862 27296 870 27304
rect 751 27055 758 27063
rect 448 26996 451 27008
rect 464 26996 470 27010
rect 543 27002 550 27014
rect 564 27008 566 27024
rect 584 27023 590 27039
rect 586 27009 590 27023
rect 348 26987 350 26996
rect 468 26987 470 26996
rect 562 26987 569 27008
rect 588 26987 590 27009
rect 636 26987 638 27049
rect 639 27041 646 27049
rect 658 27041 665 27049
rect 670 27041 690 27049
rect 639 27023 640 27041
rect 660 26993 662 27041
rect 670 27039 676 27041
rect 684 27039 686 27041
rect 680 27023 686 27039
rect 682 27009 686 27023
rect 660 26987 664 26993
rect 684 26987 686 27009
rect 732 27025 741 27055
rect 746 27031 749 27041
rect 756 27031 758 27055
rect 761 27031 768 27055
rect 778 27041 785 27063
rect 756 27025 772 27031
rect 780 27025 782 27041
rect 732 27023 736 27025
rect 732 26987 735 27023
rect 756 27015 758 27025
rect 778 27015 782 27025
rect 809 27020 812 27047
rect 814 27025 825 27047
rect 827 27025 830 27055
rect 809 27017 821 27020
rect 744 27002 748 27012
rect 754 27002 758 27015
rect 761 27002 768 27015
rect 754 27001 768 27002
rect 754 26993 758 27001
rect 754 26988 760 26993
rect 761 26988 768 27001
rect 752 26987 760 26988
rect 780 26987 782 27015
rect 876 27007 878 27304
rect 890 27296 898 27304
rect 938 27296 946 27304
rect 895 27107 906 27111
rect 907 27107 916 27279
rect 907 27095 918 27107
rect 907 27059 916 27095
rect 972 27059 974 27304
rect 986 27296 988 27304
rect 1000 27296 1002 27304
rect 1014 27296 1016 27304
rect 983 27083 999 27091
rect 880 27048 898 27059
rect 905 27048 918 27059
rect 965 27049 974 27059
rect 976 27049 982 27079
rect 983 27077 994 27079
rect 983 27049 992 27070
rect 898 27023 905 27047
rect 890 27017 906 27023
rect 876 26999 890 27007
rect 876 26987 878 26999
rect 898 26991 902 27017
rect 972 27015 974 27049
rect 975 27040 982 27049
rect 994 27040 999 27070
rect 975 27015 976 27040
rect 1008 27039 1012 27049
rect 1020 27039 1022 27304
rect 1028 27296 1030 27304
rect 1042 27079 1046 27081
rect 1040 27071 1046 27079
rect 1041 27049 1046 27051
rect 1052 27049 1058 27071
rect 1068 27059 1070 27317
rect 1092 27312 1094 27317
rect 1116 27312 1118 27317
rect 1084 27304 1094 27312
rect 1112 27304 1120 27312
rect 1076 27296 1084 27304
rect 1061 27049 1070 27059
rect 1072 27049 1078 27079
rect 1092 27049 1094 27304
rect 1104 27296 1112 27304
rect 1097 27071 1104 27079
rect 1116 27071 1118 27304
rect 1126 27149 1132 27279
rect 1126 27133 1134 27149
rect 1116 27049 1122 27071
rect 1126 27049 1132 27133
rect 1138 27079 1142 27081
rect 1136 27071 1142 27079
rect 1137 27049 1142 27051
rect 1148 27049 1154 27071
rect 1164 27067 1166 27317
rect 1212 27312 1214 27317
rect 1308 27312 1310 27317
rect 1332 27312 1334 27317
rect 1182 27304 1188 27312
rect 1210 27304 1216 27312
rect 1242 27304 1250 27312
rect 1270 27304 1284 27312
rect 1300 27304 1312 27312
rect 1328 27304 1340 27312
rect 1172 27296 1182 27304
rect 1200 27296 1210 27304
rect 1192 27132 1202 27141
rect 1202 27125 1208 27132
rect 1155 27057 1166 27067
rect 1212 27065 1214 27304
rect 1250 27296 1258 27304
rect 1284 27296 1286 27304
rect 1298 27296 1300 27304
rect 1278 27079 1284 27089
rect 1183 27057 1190 27065
rect 972 26991 976 27015
rect 982 27004 984 27014
rect 994 27004 1001 27015
rect 1018 27009 1022 27039
rect 972 26987 974 26991
rect 975 26987 976 26991
rect 992 26991 1001 27004
rect 1006 26991 1010 27004
rect 992 26990 1006 26991
rect 994 26989 1002 26990
rect 1020 26987 1022 27009
rect 1068 26987 1070 27049
rect 1071 27041 1078 27049
rect 1090 27041 1097 27049
rect 1102 27041 1122 27049
rect 1164 27041 1174 27057
rect 1071 27023 1072 27041
rect 1092 26993 1094 27041
rect 1102 27039 1108 27041
rect 1116 27039 1118 27041
rect 1112 27023 1118 27039
rect 1114 27009 1118 27023
rect 1092 26987 1096 26993
rect 1116 26987 1118 27009
rect 1164 27027 1173 27041
rect 1178 27031 1181 27041
rect 1193 27031 1200 27057
rect 1202 27041 1208 27057
rect 1210 27041 1217 27065
rect 1188 27027 1204 27031
rect 1212 27027 1214 27041
rect 1164 27023 1168 27027
rect 1164 26987 1167 27023
rect 1210 27015 1214 27027
rect 1241 27019 1244 27049
rect 1246 27027 1257 27049
rect 1259 27027 1262 27057
rect 1277 27049 1284 27059
rect 1288 27049 1294 27079
rect 1308 27049 1310 27304
rect 1312 27296 1314 27304
rect 1326 27296 1328 27304
rect 1313 27049 1320 27057
rect 1332 27049 1334 27304
rect 1340 27296 1342 27304
rect 1354 27079 1358 27081
rect 1352 27071 1358 27079
rect 1342 27049 1348 27059
rect 1353 27049 1358 27051
rect 1364 27049 1370 27071
rect 1380 27056 1382 27317
rect 1428 27312 1430 27317
rect 1524 27312 1526 27317
rect 1548 27312 1550 27317
rect 1394 27304 1404 27312
rect 1422 27304 1432 27312
rect 1454 27304 1462 27312
rect 1516 27304 1526 27312
rect 1544 27304 1554 27312
rect 1388 27296 1394 27304
rect 1416 27296 1422 27304
rect 1385 27083 1394 27084
rect 1404 27083 1411 27084
rect 1418 27083 1419 27279
rect 1428 27083 1430 27304
rect 1462 27296 1470 27304
rect 1510 27296 1516 27304
rect 1385 27082 1416 27083
rect 1418 27082 1446 27083
rect 1461 27082 1471 27104
rect 1268 27019 1272 27027
rect 1287 27019 1294 27049
rect 1306 27019 1313 27049
rect 1320 27039 1324 27049
rect 1332 27039 1338 27049
rect 1378 27046 1382 27056
rect 1328 27023 1338 27039
rect 1330 27019 1338 27023
rect 1193 26987 1200 27015
rect 1212 26987 1214 27015
rect 1252 26987 1261 27019
rect 1308 26987 1310 27019
rect 1330 27009 1334 27019
rect 1332 27001 1334 27009
rect 1328 26987 1334 27001
rect 1380 26987 1382 27046
rect 1388 27041 1390 27046
rect 1408 27041 1412 27056
rect 1416 27041 1418 27071
rect 1428 27041 1430 27082
rect 1512 27079 1520 27090
rect 1524 27087 1526 27304
rect 1538 27296 1544 27304
rect 1504 27074 1512 27079
rect 1514 27074 1520 27079
rect 1522 27074 1529 27087
rect 1544 27079 1547 27092
rect 1433 27041 1434 27071
rect 1514 27049 1521 27074
rect 1524 27049 1526 27074
rect 1394 27036 1430 27041
rect 1464 27038 1478 27046
rect 1394 27032 1402 27036
rect 1408 27032 1412 27036
rect 1394 27031 1398 27032
rect 1404 27015 1408 27031
rect 1406 27012 1408 27015
rect 1414 27012 1420 27020
rect 1406 27001 1420 27012
rect 1428 27010 1430 27036
rect 1522 27024 1529 27049
rect 1536 27039 1540 27049
rect 1548 27039 1550 27304
rect 1570 27079 1574 27081
rect 1568 27071 1574 27079
rect 1569 27049 1574 27051
rect 1580 27049 1586 27071
rect 1596 27059 1598 27317
rect 1620 27312 1622 27317
rect 1644 27312 1646 27317
rect 1612 27304 1622 27312
rect 1640 27304 1648 27312
rect 1604 27296 1612 27304
rect 1589 27049 1598 27059
rect 1600 27049 1606 27079
rect 1620 27049 1622 27304
rect 1632 27296 1640 27304
rect 1625 27071 1632 27079
rect 1644 27071 1646 27304
rect 1654 27149 1660 27279
rect 1654 27133 1662 27149
rect 1644 27049 1650 27071
rect 1654 27049 1660 27133
rect 1666 27079 1670 27081
rect 1664 27071 1670 27079
rect 1665 27049 1670 27051
rect 1676 27049 1682 27071
rect 1692 27059 1694 27317
rect 1716 27312 1718 27317
rect 1740 27312 1742 27317
rect 1708 27304 1718 27312
rect 1736 27304 1744 27312
rect 1700 27296 1708 27304
rect 1685 27049 1694 27059
rect 1696 27049 1702 27079
rect 1716 27049 1718 27304
rect 1728 27296 1736 27304
rect 1721 27071 1728 27079
rect 1740 27071 1742 27304
rect 1750 27149 1756 27279
rect 1750 27133 1758 27149
rect 1740 27049 1746 27071
rect 1750 27049 1756 27133
rect 1762 27079 1766 27081
rect 1760 27071 1766 27079
rect 1761 27049 1766 27051
rect 1772 27049 1778 27071
rect 1788 27059 1790 27317
rect 1812 27312 1814 27317
rect 1836 27312 1838 27317
rect 1804 27304 1814 27312
rect 1832 27304 1840 27312
rect 1796 27296 1804 27304
rect 1781 27049 1790 27059
rect 1792 27049 1798 27079
rect 1812 27049 1814 27304
rect 1824 27296 1832 27304
rect 1817 27071 1824 27079
rect 1836 27071 1838 27304
rect 1846 27149 1852 27279
rect 1846 27133 1854 27149
rect 1836 27049 1842 27071
rect 1846 27049 1852 27133
rect 1858 27079 1862 27081
rect 1856 27071 1862 27079
rect 1857 27049 1862 27051
rect 1868 27049 1874 27071
rect 1884 27059 1886 27317
rect 1908 27312 1910 27317
rect 1932 27312 1934 27317
rect 1900 27304 1910 27312
rect 1928 27304 1936 27312
rect 1892 27296 1900 27304
rect 1877 27049 1886 27059
rect 1888 27049 1894 27079
rect 1908 27049 1910 27304
rect 1920 27296 1928 27304
rect 1913 27071 1920 27079
rect 1932 27071 1934 27304
rect 1942 27149 1948 27279
rect 1942 27133 1950 27149
rect 1932 27049 1938 27071
rect 1942 27049 1948 27133
rect 1954 27079 1958 27081
rect 1952 27071 1958 27079
rect 1953 27049 1958 27051
rect 1964 27049 1970 27071
rect 1980 27059 1982 27317
rect 2004 27312 2006 27317
rect 2028 27312 2030 27317
rect 1996 27304 2006 27312
rect 2024 27304 2032 27312
rect 1988 27296 1996 27304
rect 1973 27049 1982 27059
rect 1984 27049 1990 27079
rect 2004 27049 2006 27304
rect 2016 27296 2024 27304
rect 2009 27071 2016 27079
rect 2028 27071 2030 27304
rect 2038 27149 2044 27279
rect 2038 27133 2046 27149
rect 2028 27049 2034 27071
rect 2038 27049 2044 27133
rect 2050 27079 2054 27081
rect 2048 27071 2054 27079
rect 2049 27049 2054 27051
rect 2060 27049 2066 27071
rect 2076 27059 2078 27317
rect 2100 27312 2102 27317
rect 2124 27312 2126 27317
rect 2092 27304 2102 27312
rect 2120 27304 2128 27312
rect 2084 27296 2092 27304
rect 2069 27049 2078 27059
rect 2080 27049 2086 27079
rect 2100 27049 2102 27304
rect 2112 27296 2120 27304
rect 2105 27071 2112 27079
rect 2124 27071 2126 27304
rect 2134 27149 2140 27279
rect 2134 27133 2142 27149
rect 2124 27049 2130 27071
rect 2134 27049 2140 27133
rect 2146 27079 2150 27081
rect 2144 27071 2150 27079
rect 2145 27049 2150 27051
rect 2156 27049 2162 27071
rect 2172 27059 2174 27317
rect 2196 27312 2198 27317
rect 2220 27312 2222 27317
rect 2188 27304 2198 27312
rect 2216 27304 2224 27312
rect 2180 27296 2188 27304
rect 2165 27049 2174 27059
rect 2176 27049 2182 27079
rect 2196 27049 2198 27304
rect 2208 27296 2216 27304
rect 2201 27071 2208 27079
rect 2220 27071 2222 27304
rect 2230 27149 2236 27279
rect 2230 27133 2238 27149
rect 2220 27049 2226 27071
rect 2230 27049 2236 27133
rect 2242 27079 2246 27081
rect 2240 27071 2246 27079
rect 2241 27049 2246 27051
rect 2252 27049 2258 27071
rect 2268 27059 2270 27317
rect 2292 27312 2294 27317
rect 2316 27312 2318 27317
rect 2284 27304 2294 27312
rect 2312 27304 2320 27312
rect 2276 27296 2284 27304
rect 2261 27049 2270 27059
rect 2272 27049 2278 27079
rect 2292 27049 2294 27304
rect 2304 27296 2312 27304
rect 2297 27071 2304 27079
rect 2316 27071 2318 27304
rect 2326 27149 2332 27279
rect 2326 27133 2334 27149
rect 2316 27049 2322 27071
rect 2326 27049 2332 27133
rect 2338 27079 2342 27081
rect 2336 27071 2342 27079
rect 2337 27049 2342 27051
rect 2348 27049 2354 27071
rect 2364 27059 2366 27317
rect 2388 27312 2390 27317
rect 2412 27312 2414 27317
rect 2380 27304 2390 27312
rect 2408 27304 2416 27312
rect 2372 27296 2380 27304
rect 2357 27049 2366 27059
rect 2368 27049 2374 27079
rect 2388 27049 2390 27304
rect 2400 27296 2408 27304
rect 2393 27071 2400 27079
rect 2412 27071 2414 27304
rect 2422 27149 2428 27279
rect 2422 27133 2430 27149
rect 2412 27049 2418 27071
rect 2422 27049 2428 27133
rect 2434 27079 2438 27081
rect 2432 27071 2438 27079
rect 2433 27049 2438 27051
rect 2444 27049 2450 27071
rect 2460 27059 2462 27317
rect 2484 27312 2486 27317
rect 2508 27312 2510 27317
rect 2476 27304 2486 27312
rect 2504 27304 2512 27312
rect 2468 27296 2476 27304
rect 2453 27049 2462 27059
rect 2464 27049 2470 27079
rect 2484 27049 2486 27304
rect 2496 27296 2504 27304
rect 2489 27071 2496 27079
rect 2508 27071 2510 27304
rect 2518 27149 2524 27279
rect 2518 27133 2526 27149
rect 2508 27049 2514 27071
rect 2518 27049 2524 27133
rect 2530 27079 2534 27081
rect 2528 27071 2534 27079
rect 2529 27049 2534 27051
rect 2540 27049 2546 27071
rect 2556 27059 2558 27317
rect 2580 27312 2582 27317
rect 2604 27312 2606 27317
rect 2572 27304 2582 27312
rect 2600 27304 2608 27312
rect 2564 27296 2572 27304
rect 2549 27049 2558 27059
rect 2560 27049 2566 27079
rect 2580 27049 2582 27304
rect 2592 27296 2600 27304
rect 2585 27071 2592 27079
rect 2604 27071 2606 27304
rect 2614 27149 2620 27279
rect 2614 27133 2622 27149
rect 2604 27049 2610 27071
rect 2614 27049 2620 27133
rect 2626 27079 2630 27081
rect 2624 27071 2630 27079
rect 2625 27049 2630 27051
rect 2636 27049 2642 27071
rect 2652 27059 2654 27317
rect 2676 27312 2678 27317
rect 2700 27312 2702 27317
rect 2668 27304 2678 27312
rect 2696 27304 2704 27312
rect 2660 27296 2668 27304
rect 2645 27049 2654 27059
rect 2656 27049 2662 27079
rect 2676 27049 2678 27304
rect 2688 27296 2696 27304
rect 2681 27071 2688 27079
rect 2700 27071 2702 27304
rect 2710 27149 2716 27279
rect 2710 27133 2718 27149
rect 2700 27049 2706 27071
rect 2710 27049 2716 27133
rect 2722 27079 2726 27081
rect 2720 27071 2726 27079
rect 2721 27049 2726 27051
rect 2732 27049 2738 27071
rect 2748 27059 2750 27317
rect 2772 27312 2774 27317
rect 2796 27312 2798 27317
rect 2764 27304 2774 27312
rect 2792 27304 2800 27312
rect 2824 27304 2840 27312
rect 2756 27296 2764 27304
rect 2741 27049 2750 27059
rect 2752 27049 2758 27079
rect 2772 27049 2774 27304
rect 2784 27296 2792 27304
rect 2777 27071 2784 27079
rect 2796 27071 2798 27304
rect 2806 27149 2812 27279
rect 2806 27133 2814 27149
rect 2796 27049 2802 27071
rect 2806 27049 2812 27133
rect 2832 27096 2836 27106
rect 2844 27096 2846 27317
rect 2868 27312 2870 27317
rect 2892 27312 2894 27317
rect 2856 27304 2870 27312
rect 2884 27304 2896 27312
rect 2916 27304 2924 27312
rect 2852 27296 2856 27304
rect 2842 27082 2846 27096
rect 2818 27079 2822 27081
rect 2816 27071 2822 27079
rect 2828 27079 2846 27082
rect 2828 27071 2853 27079
rect 2817 27049 2822 27051
rect 2828 27049 2834 27071
rect 2842 27066 2853 27071
rect 1424 26996 1430 27010
rect 1503 27002 1510 27014
rect 1524 27008 1526 27024
rect 1544 27023 1550 27039
rect 1546 27009 1550 27023
rect 1428 26987 1430 26996
rect 1522 26987 1529 27008
rect 1548 26987 1550 27009
rect 1596 26987 1598 27049
rect 1599 27041 1606 27049
rect 1618 27041 1625 27049
rect 1630 27041 1650 27049
rect 1599 27023 1600 27041
rect 1620 26993 1622 27041
rect 1630 27039 1636 27041
rect 1644 27039 1646 27041
rect 1640 27023 1646 27039
rect 1642 27009 1646 27023
rect 1620 26987 1624 26993
rect 1644 26987 1646 27009
rect 1692 26987 1694 27049
rect 1695 27041 1702 27049
rect 1714 27041 1721 27049
rect 1726 27041 1746 27049
rect 1695 27023 1696 27041
rect 1716 26993 1718 27041
rect 1726 27039 1732 27041
rect 1740 27039 1742 27041
rect 1736 27023 1742 27039
rect 1738 27009 1742 27023
rect 1716 26987 1720 26993
rect 1740 26987 1742 27009
rect 1788 26987 1790 27049
rect 1791 27041 1798 27049
rect 1810 27041 1817 27049
rect 1822 27041 1842 27049
rect 1791 27023 1792 27041
rect 1812 26993 1814 27041
rect 1822 27039 1828 27041
rect 1836 27039 1838 27041
rect 1832 27023 1838 27039
rect 1834 27009 1838 27023
rect 1812 26987 1816 26993
rect 1836 26987 1838 27009
rect 1884 26987 1886 27049
rect 1887 27041 1894 27049
rect 1906 27041 1913 27049
rect 1918 27041 1938 27049
rect 1887 27023 1888 27041
rect 1908 26993 1910 27041
rect 1918 27039 1924 27041
rect 1932 27039 1934 27041
rect 1928 27023 1934 27039
rect 1930 27009 1934 27023
rect 1908 26987 1912 26993
rect 1932 26987 1934 27009
rect 1980 26987 1982 27049
rect 1983 27041 1990 27049
rect 2002 27041 2009 27049
rect 2014 27041 2034 27049
rect 1983 27023 1984 27041
rect 2004 26993 2006 27041
rect 2014 27039 2020 27041
rect 2028 27039 2030 27041
rect 2024 27023 2030 27039
rect 2026 27009 2030 27023
rect 2004 26987 2008 26993
rect 2028 26987 2030 27009
rect 2076 26987 2078 27049
rect 2079 27041 2086 27049
rect 2098 27041 2105 27049
rect 2110 27041 2130 27049
rect 2079 27023 2080 27041
rect 2100 26993 2102 27041
rect 2110 27039 2116 27041
rect 2124 27039 2126 27041
rect 2120 27023 2126 27039
rect 2122 27009 2126 27023
rect 2100 26987 2104 26993
rect 2124 26987 2126 27009
rect 2172 26987 2174 27049
rect 2175 27041 2182 27049
rect 2194 27041 2201 27049
rect 2206 27041 2226 27049
rect 2175 27023 2176 27041
rect 2196 26993 2198 27041
rect 2206 27039 2212 27041
rect 2220 27039 2222 27041
rect 2216 27023 2222 27039
rect 2218 27009 2222 27023
rect 2196 26987 2200 26993
rect 2220 26987 2222 27009
rect 2268 26987 2270 27049
rect 2271 27041 2278 27049
rect 2290 27041 2297 27049
rect 2302 27041 2322 27049
rect 2271 27023 2272 27041
rect 2292 26993 2294 27041
rect 2302 27039 2308 27041
rect 2316 27039 2318 27041
rect 2312 27023 2318 27039
rect 2314 27009 2318 27023
rect 2292 26987 2296 26993
rect 2316 26987 2318 27009
rect 2364 26987 2366 27049
rect 2367 27041 2374 27049
rect 2386 27041 2393 27049
rect 2398 27041 2418 27049
rect 2367 27023 2368 27041
rect 2388 26993 2390 27041
rect 2398 27039 2404 27041
rect 2412 27039 2414 27041
rect 2408 27023 2414 27039
rect 2410 27009 2414 27023
rect 2388 26987 2392 26993
rect 2412 26987 2414 27009
rect 2460 26987 2462 27049
rect 2463 27041 2470 27049
rect 2482 27041 2489 27049
rect 2494 27041 2514 27049
rect 2463 27023 2464 27041
rect 2484 26993 2486 27041
rect 2494 27039 2500 27041
rect 2508 27039 2510 27041
rect 2504 27023 2510 27039
rect 2506 27009 2510 27023
rect 2484 26987 2488 26993
rect 2508 26987 2510 27009
rect 2556 26987 2558 27049
rect 2559 27041 2566 27049
rect 2578 27041 2585 27049
rect 2590 27041 2610 27049
rect 2559 27023 2560 27041
rect 2580 26993 2582 27041
rect 2590 27039 2596 27041
rect 2604 27039 2606 27041
rect 2600 27023 2606 27039
rect 2602 27009 2606 27023
rect 2580 26987 2584 26993
rect 2604 26987 2606 27009
rect 2652 26987 2654 27049
rect 2655 27041 2662 27049
rect 2674 27041 2681 27049
rect 2686 27041 2706 27049
rect 2655 27023 2656 27041
rect 2676 26993 2678 27041
rect 2686 27039 2692 27041
rect 2700 27039 2702 27041
rect 2696 27023 2702 27039
rect 2698 27009 2702 27023
rect 2676 26987 2680 26993
rect 2700 26987 2702 27009
rect 2748 26987 2750 27049
rect 2751 27041 2758 27049
rect 2770 27041 2777 27049
rect 2782 27041 2802 27049
rect 2844 27041 2846 27066
rect 2751 27023 2752 27041
rect 2772 26993 2774 27041
rect 2782 27039 2788 27041
rect 2796 27039 2798 27041
rect 2792 27023 2798 27039
rect 2794 27009 2798 27023
rect 2772 26987 2776 26993
rect 2796 26987 2798 27009
rect 2841 27023 2848 27041
rect 2860 27031 2867 27066
rect 2868 27031 2870 27304
rect 2880 27296 2884 27304
rect 2873 27071 2880 27079
rect 2892 27071 2894 27304
rect 2924 27296 2932 27304
rect 2940 27096 2942 27317
rect 3012 27312 3014 27317
rect 2944 27304 2952 27312
rect 3006 27304 3016 27312
rect 3034 27304 3044 27312
rect 3066 27304 3074 27312
rect 3094 27304 3106 27312
rect 3108 27304 3110 27317
rect 3156 27312 3158 27317
rect 3252 27312 3254 27317
rect 3122 27304 3134 27312
rect 3150 27304 3162 27312
rect 3182 27304 3190 27312
rect 3246 27304 3254 27312
rect 3274 27304 3282 27312
rect 3306 27304 3314 27312
rect 3334 27304 3346 27312
rect 3348 27304 3350 27317
rect 3396 27312 3398 27317
rect 3362 27304 3374 27312
rect 3390 27304 3402 27312
rect 3422 27304 3430 27312
rect 3450 27304 3466 27312
rect 2952 27296 2960 27304
rect 3000 27296 3006 27304
rect 2936 27088 2942 27096
rect 2873 27066 2877 27071
rect 2887 27051 2894 27071
rect 2918 27058 2921 27088
rect 2940 27066 2943 27088
rect 2963 27066 2966 27096
rect 2926 27059 2934 27066
rect 2940 27059 2942 27066
rect 2943 27061 2948 27066
rect 2943 27059 2957 27061
rect 2926 27058 2957 27059
rect 2926 27056 2927 27058
rect 2928 27056 2932 27058
rect 2940 27056 2942 27058
rect 2887 27047 2898 27051
rect 2882 27041 2898 27047
rect 2873 27031 2877 27041
rect 2841 26987 2847 27023
rect 2860 27020 2863 27031
rect 2856 27010 2863 27020
rect 2868 27020 2877 27031
rect 2868 27015 2878 27020
rect 2860 26990 2863 27010
rect 2866 27010 2870 27015
rect 2873 27010 2878 27015
rect 2887 27015 2894 27041
rect 2936 27040 2937 27056
rect 2938 27026 2942 27056
rect 2866 27001 2880 27010
rect 2866 26996 2870 27001
rect 2873 26996 2878 27001
rect 2852 26987 2863 26990
rect 2868 26993 2870 26996
rect 2868 26987 2872 26993
rect 2887 26987 2890 27015
rect 2892 26987 2894 27015
rect 2940 27004 2942 27026
rect 2927 26994 2930 26998
rect 2927 26988 2931 26994
rect 2936 26987 2942 27004
rect 3012 27023 3014 27304
rect 3028 27296 3034 27304
rect 3074 27296 3082 27304
rect 3106 27296 3110 27304
rect 3134 27296 3138 27304
rect 3031 27118 3042 27119
rect 3043 27100 3052 27279
rect 3043 27091 3054 27100
rect 3017 27049 3024 27078
rect 3026 27058 3032 27078
rect 3034 27058 3041 27086
rect 3043 27058 3052 27091
rect 3028 27049 3031 27051
rect 3016 27048 3031 27049
rect 3034 27032 3038 27058
rect 3108 27056 3110 27296
rect 3108 27055 3119 27056
rect 3108 27025 3117 27055
rect 3119 27040 3125 27055
rect 3127 27040 3134 27063
rect 3012 27018 3016 27023
rect 3026 27018 3028 27023
rect 3012 27010 3014 27018
rect 3012 26996 3016 27010
rect 3012 26987 3017 26996
rect 3108 26987 3112 27025
rect 3118 27004 3120 27014
rect 3128 27002 3130 27004
rect 3142 27002 3144 27004
rect 3128 26998 3142 27002
rect 3118 26990 3142 26998
rect 3118 26989 3128 26990
rect 3130 26989 3138 26990
rect 3156 26987 3158 27304
rect 3162 27296 3166 27304
rect 3190 27296 3198 27304
rect 3238 27296 3246 27304
rect 3185 27020 3188 27047
rect 3190 27025 3201 27047
rect 3203 27025 3206 27055
rect 3185 27017 3197 27020
rect 3252 27007 3254 27304
rect 3266 27296 3274 27304
rect 3314 27296 3322 27304
rect 3346 27296 3350 27304
rect 3374 27296 3378 27304
rect 3271 27107 3282 27111
rect 3283 27107 3292 27279
rect 3283 27095 3294 27107
rect 3283 27059 3292 27095
rect 3256 27048 3274 27059
rect 3281 27048 3294 27059
rect 3348 27056 3350 27296
rect 3348 27055 3359 27056
rect 3274 27023 3281 27047
rect 3348 27025 3357 27055
rect 3359 27040 3365 27055
rect 3367 27040 3374 27063
rect 3266 27017 3282 27023
rect 3252 26999 3266 27007
rect 3252 26987 3254 26999
rect 3274 26991 3278 27017
rect 3348 26987 3352 27025
rect 3358 27004 3360 27014
rect 3368 27002 3370 27004
rect 3382 27002 3384 27004
rect 3368 26998 3382 27002
rect 3358 26990 3382 26998
rect 3358 26989 3368 26990
rect 3370 26989 3378 26990
rect 3396 26987 3398 27304
rect 3402 27296 3406 27304
rect 3430 27296 3438 27304
rect 3468 27055 3470 27317
rect 3492 27312 3494 27317
rect 3516 27312 3518 27317
rect 3482 27304 3494 27312
rect 3510 27304 3522 27312
rect 3542 27304 3550 27312
rect 3570 27304 3586 27312
rect 3478 27296 3482 27304
rect 3425 27020 3428 27047
rect 3430 27025 3441 27047
rect 3443 27025 3446 27055
rect 3468 27025 3477 27055
rect 3492 27025 3494 27304
rect 3506 27296 3510 27304
rect 3497 27025 3504 27055
rect 3516 27047 3518 27304
rect 3550 27296 3558 27304
rect 3588 27055 3590 27317
rect 3612 27312 3614 27317
rect 3636 27312 3638 27317
rect 3602 27304 3614 27312
rect 3630 27304 3642 27312
rect 3662 27304 3670 27312
rect 3598 27296 3602 27304
rect 3425 27017 3437 27020
rect 3468 26987 3470 27025
rect 3487 27017 3494 27025
rect 3514 27017 3521 27047
rect 3545 27020 3548 27047
rect 3550 27025 3561 27047
rect 3563 27025 3566 27055
rect 3588 27025 3597 27055
rect 3612 27025 3614 27304
rect 3626 27296 3630 27304
rect 3617 27025 3624 27055
rect 3636 27047 3638 27304
rect 3670 27296 3678 27304
rect 3545 27017 3557 27020
rect 3480 27002 3484 27012
rect 3492 27002 3494 27017
rect 3497 27007 3504 27017
rect 3490 26988 3504 27002
rect 3514 26991 3518 27017
rect 3491 26987 3504 26988
rect 3516 26987 3518 26991
rect 3588 26987 3590 27025
rect 3607 27017 3614 27025
rect 3634 27017 3641 27047
rect 3665 27020 3668 27047
rect 3670 27025 3681 27047
rect 3683 27025 3686 27055
rect 3665 27017 3677 27020
rect 3600 27002 3604 27012
rect 3612 27002 3614 27017
rect 3617 27007 3624 27017
rect 3610 26988 3624 27002
rect 3634 26991 3638 27017
rect 3611 26987 3624 26988
rect 3636 26987 3638 26991
rect 3708 26987 3710 27317
rect 3732 27312 3734 27317
rect 3756 27312 3758 27317
rect 3724 27304 3734 27312
rect 3752 27304 3762 27312
rect 3718 27296 3724 27304
rect 3712 27049 3730 27059
rect 3732 27047 3734 27304
rect 3746 27296 3752 27304
rect 3756 27059 3758 27304
rect 3737 27049 3758 27059
rect 3766 27049 3772 27279
rect 3778 27079 3782 27081
rect 3776 27071 3782 27079
rect 3777 27049 3782 27051
rect 3788 27049 3794 27071
rect 3804 27059 3806 27317
rect 3828 27312 3830 27317
rect 3852 27312 3854 27317
rect 3820 27304 3830 27312
rect 3848 27304 3856 27312
rect 3812 27296 3820 27304
rect 3797 27049 3806 27059
rect 3808 27049 3814 27079
rect 3828 27049 3830 27304
rect 3840 27296 3848 27304
rect 3833 27071 3840 27079
rect 3852 27071 3854 27304
rect 3862 27149 3868 27279
rect 3862 27133 3870 27149
rect 3852 27049 3858 27071
rect 3862 27049 3868 27133
rect 3874 27079 3878 27081
rect 3872 27071 3878 27079
rect 3873 27049 3878 27051
rect 3884 27049 3890 27071
rect 3900 27059 3902 27317
rect 3924 27312 3926 27317
rect 3948 27312 3950 27317
rect 3916 27304 3926 27312
rect 3944 27304 3952 27312
rect 3908 27296 3916 27304
rect 3893 27049 3902 27059
rect 3904 27049 3910 27079
rect 3924 27049 3926 27304
rect 3936 27296 3944 27304
rect 3929 27071 3936 27079
rect 3948 27071 3950 27304
rect 3958 27149 3964 27279
rect 3958 27133 3966 27149
rect 3948 27049 3954 27071
rect 3958 27049 3964 27133
rect 3970 27079 3974 27081
rect 3968 27071 3974 27079
rect 3969 27049 3974 27051
rect 3980 27049 3986 27071
rect 3996 27059 3998 27317
rect 4020 27312 4022 27317
rect 4044 27312 4046 27317
rect 4012 27304 4022 27312
rect 4040 27304 4048 27312
rect 4004 27296 4012 27304
rect 3989 27049 3998 27059
rect 4000 27049 4006 27079
rect 4020 27049 4022 27304
rect 4032 27296 4040 27304
rect 4025 27071 4032 27079
rect 4044 27071 4046 27304
rect 4054 27149 4060 27279
rect 4054 27133 4062 27149
rect 4044 27049 4050 27071
rect 4054 27049 4060 27133
rect 4066 27079 4070 27081
rect 4064 27071 4070 27079
rect 4065 27049 4070 27051
rect 4076 27049 4082 27071
rect 4092 27059 4094 27317
rect 4116 27312 4118 27317
rect 4140 27312 4142 27317
rect 4108 27304 4118 27312
rect 4136 27304 4144 27312
rect 4100 27296 4108 27304
rect 4085 27049 4094 27059
rect 4096 27049 4102 27079
rect 4116 27049 4118 27304
rect 4128 27296 4136 27304
rect 4121 27071 4128 27079
rect 4140 27071 4142 27304
rect 4150 27149 4156 27279
rect 4150 27133 4158 27149
rect 4140 27049 4146 27071
rect 4150 27049 4156 27133
rect 4162 27079 4166 27081
rect 4160 27071 4166 27079
rect 4161 27049 4166 27051
rect 4172 27049 4178 27071
rect 4188 27059 4190 27317
rect 4212 27312 4214 27317
rect 4236 27312 4238 27317
rect 4204 27304 4214 27312
rect 4232 27304 4240 27312
rect 4196 27296 4204 27304
rect 4181 27049 4190 27059
rect 4192 27049 4198 27079
rect 4212 27049 4214 27304
rect 4224 27296 4232 27304
rect 4217 27071 4224 27079
rect 4236 27071 4238 27304
rect 4246 27149 4252 27279
rect 4246 27133 4254 27149
rect 4236 27049 4242 27071
rect 4246 27049 4252 27133
rect 4258 27079 4262 27081
rect 4256 27071 4262 27079
rect 4257 27049 4262 27051
rect 4268 27049 4274 27071
rect 4284 27059 4286 27317
rect 4308 27312 4310 27317
rect 4332 27312 4334 27317
rect 4300 27304 4310 27312
rect 4328 27304 4336 27312
rect 4292 27296 4300 27304
rect 4277 27049 4286 27059
rect 4288 27049 4294 27079
rect 4308 27049 4310 27304
rect 4320 27296 4328 27304
rect 4313 27071 4320 27079
rect 4332 27071 4334 27304
rect 4342 27149 4348 27279
rect 4342 27133 4350 27149
rect 4332 27049 4338 27071
rect 4342 27049 4348 27133
rect 4354 27079 4358 27081
rect 4352 27071 4358 27079
rect 4353 27049 4358 27051
rect 4364 27049 4370 27071
rect 4380 27059 4382 27317
rect 4404 27312 4406 27317
rect 4428 27312 4430 27317
rect 4396 27304 4406 27312
rect 4424 27304 4432 27312
rect 4388 27296 4396 27304
rect 4373 27049 4382 27059
rect 4384 27049 4390 27079
rect 4404 27049 4406 27304
rect 4416 27296 4424 27304
rect 4409 27071 4416 27079
rect 4428 27071 4430 27304
rect 4438 27149 4444 27279
rect 4438 27133 4446 27149
rect 4428 27049 4434 27071
rect 4438 27049 4444 27133
rect 4450 27079 4454 27081
rect 4448 27071 4454 27079
rect 4449 27049 4454 27051
rect 4460 27049 4466 27071
rect 4476 27059 4478 27317
rect 4500 27312 4502 27317
rect 4524 27312 4526 27317
rect 4596 27312 4598 27317
rect 4492 27304 4502 27312
rect 4520 27304 4528 27312
rect 4590 27304 4598 27312
rect 4618 27304 4624 27312
rect 4650 27304 4658 27312
rect 4678 27304 4694 27312
rect 4710 27304 4722 27312
rect 4738 27304 4750 27312
rect 4770 27304 4778 27312
rect 4798 27304 4808 27312
rect 4812 27304 4814 27317
rect 4860 27312 4862 27317
rect 4826 27304 4836 27312
rect 4854 27304 4864 27312
rect 4884 27304 4892 27312
rect 4484 27296 4492 27304
rect 4469 27049 4478 27059
rect 4480 27049 4486 27079
rect 4500 27049 4502 27304
rect 4512 27296 4520 27304
rect 4505 27071 4512 27079
rect 4524 27071 4526 27304
rect 4580 27296 4590 27304
rect 4534 27149 4540 27279
rect 4534 27133 4542 27149
rect 4524 27049 4530 27071
rect 4534 27049 4540 27133
rect 4546 27079 4550 27081
rect 4544 27071 4550 27079
rect 4545 27049 4550 27051
rect 4556 27049 4562 27071
rect 3730 27017 3737 27047
rect 3744 27039 3748 27049
rect 3756 27047 3758 27049
rect 3756 27039 3762 27047
rect 3752 27023 3762 27039
rect 3754 27017 3762 27023
rect 3732 26991 3734 27017
rect 3754 27009 3758 27017
rect 3732 26987 3746 26991
rect 3756 26987 3758 27009
rect 3804 26987 3806 27049
rect 3807 27041 3814 27049
rect 3826 27041 3833 27049
rect 3838 27041 3858 27049
rect 3807 27023 3808 27041
rect 3828 26993 3830 27041
rect 3838 27039 3844 27041
rect 3852 27039 3854 27041
rect 3848 27023 3854 27039
rect 3850 27009 3854 27023
rect 3828 26987 3832 26993
rect 3852 26987 3854 27009
rect 3900 26987 3902 27049
rect 3903 27041 3910 27049
rect 3922 27041 3929 27049
rect 3934 27041 3954 27049
rect 3903 27023 3904 27041
rect 3924 26993 3926 27041
rect 3934 27039 3940 27041
rect 3948 27039 3950 27041
rect 3944 27023 3950 27039
rect 3946 27009 3950 27023
rect 3924 26987 3928 26993
rect 3948 26987 3950 27009
rect 3996 26987 3998 27049
rect 3999 27041 4006 27049
rect 4018 27041 4025 27049
rect 4030 27041 4050 27049
rect 3999 27023 4000 27041
rect 4020 26993 4022 27041
rect 4030 27039 4036 27041
rect 4044 27039 4046 27041
rect 4040 27023 4046 27039
rect 4042 27009 4046 27023
rect 4020 26987 4024 26993
rect 4044 26987 4046 27009
rect 4092 26987 4094 27049
rect 4095 27041 4102 27049
rect 4114 27041 4121 27049
rect 4126 27041 4146 27049
rect 4095 27023 4096 27041
rect 4116 26993 4118 27041
rect 4126 27039 4132 27041
rect 4140 27039 4142 27041
rect 4136 27023 4142 27039
rect 4138 27009 4142 27023
rect 4116 26987 4120 26993
rect 4140 26987 4142 27009
rect 4188 26987 4190 27049
rect 4191 27041 4198 27049
rect 4210 27041 4217 27049
rect 4222 27041 4242 27049
rect 4191 27023 4192 27041
rect 4212 26993 4214 27041
rect 4222 27039 4228 27041
rect 4236 27039 4238 27041
rect 4232 27023 4238 27039
rect 4234 27009 4238 27023
rect 4212 26987 4216 26993
rect 4236 26987 4238 27009
rect 4284 26987 4286 27049
rect 4287 27041 4294 27049
rect 4306 27041 4313 27049
rect 4318 27041 4338 27049
rect 4287 27023 4288 27041
rect 4308 26993 4310 27041
rect 4318 27039 4324 27041
rect 4332 27039 4334 27041
rect 4328 27023 4334 27039
rect 4330 27009 4334 27023
rect 4308 26987 4312 26993
rect 4332 26987 4334 27009
rect 4380 26987 4382 27049
rect 4383 27041 4390 27049
rect 4402 27041 4409 27049
rect 4414 27041 4434 27049
rect 4383 27023 4384 27041
rect 4404 26993 4406 27041
rect 4414 27039 4420 27041
rect 4428 27039 4430 27041
rect 4424 27023 4430 27039
rect 4426 27009 4430 27023
rect 4404 26987 4408 26993
rect 4428 26987 4430 27009
rect 4476 26987 4478 27049
rect 4479 27041 4486 27049
rect 4498 27041 4505 27049
rect 4510 27041 4530 27049
rect 4479 27023 4480 27041
rect 4500 26993 4502 27041
rect 4510 27039 4516 27041
rect 4524 27039 4526 27041
rect 4520 27023 4526 27039
rect 4522 27009 4526 27023
rect 4500 26987 4504 26993
rect 4524 26987 4526 27009
rect 4596 27013 4598 27304
rect 4608 27296 4618 27304
rect 4658 27296 4666 27304
rect 4706 27296 4710 27304
rect 4734 27296 4738 27304
rect 4778 27296 4786 27304
rect 4808 27296 4814 27304
rect 4836 27296 4842 27304
rect 4601 27048 4608 27078
rect 4610 27048 4616 27071
rect 4618 27041 4625 27071
rect 4627 27048 4636 27279
rect 4800 27096 4804 27106
rect 4812 27096 4814 27296
rect 4828 27096 4835 27099
rect 4708 27083 4719 27090
rect 4710 27078 4719 27083
rect 4810 27082 4814 27096
rect 4823 27083 4839 27096
rect 4796 27078 4814 27082
rect 4720 27048 4731 27078
rect 4796 27070 4821 27078
rect 4826 27070 4839 27082
rect 4810 27066 4821 27070
rect 4823 27066 4826 27070
rect 4828 27066 4835 27070
rect 4610 27013 4612 27023
rect 4618 27015 4622 27041
rect 4720 27040 4729 27048
rect 4812 27040 4814 27066
rect 4823 27040 4835 27066
rect 4848 27051 4852 27061
rect 4860 27051 4862 27304
rect 4864 27296 4870 27304
rect 4892 27296 4900 27304
rect 4908 27096 4910 27317
rect 4912 27304 4920 27312
rect 4940 27304 4954 27312
rect 4956 27304 4958 27317
rect 4980 27312 4982 27317
rect 5004 27312 5006 27317
rect 4970 27304 4982 27312
rect 4998 27304 5010 27312
rect 5030 27304 5038 27312
rect 4920 27296 4928 27304
rect 4954 27296 4958 27304
rect 4968 27296 4970 27304
rect 4980 27296 4984 27304
rect 4996 27296 4998 27304
rect 4904 27088 4910 27096
rect 4886 27058 4889 27088
rect 4908 27066 4911 27088
rect 4931 27066 4934 27096
rect 4956 27067 4958 27296
rect 4980 27067 4982 27296
rect 5004 27067 5006 27304
rect 5010 27296 5012 27304
rect 5038 27296 5046 27304
rect 4894 27059 4902 27066
rect 4908 27059 4910 27066
rect 4911 27061 4916 27066
rect 4911 27059 4925 27061
rect 4894 27058 4925 27059
rect 4945 27058 4958 27067
rect 4965 27058 4985 27067
rect 4992 27058 5010 27067
rect 4894 27056 4895 27058
rect 4896 27056 4900 27058
rect 4908 27056 4910 27058
rect 4720 27013 4722 27015
rect 4596 27001 4610 27013
rect 4620 27001 4622 27013
rect 4712 27004 4722 27013
rect 4596 26993 4598 27001
rect 4716 26999 4726 27004
rect 4596 26987 4600 26993
rect 4720 26989 4722 26990
rect 4809 26987 4816 27040
rect 4822 27004 4824 27014
rect 4828 27005 4831 27040
rect 4858 27037 4862 27051
rect 4904 27040 4905 27056
rect 4832 27005 4842 27010
rect 4832 27004 4845 27005
rect 4832 26996 4846 27004
rect 4829 26990 4845 26996
rect 4829 26989 4832 26990
rect 4828 26987 4831 26989
rect 4860 26987 4862 27037
rect 4906 27026 4910 27056
rect 4908 27004 4910 27026
rect 4895 26994 4898 26998
rect 4895 26988 4899 26994
rect 4904 26987 4910 27004
rect 4956 27055 4958 27058
rect 4956 27025 4965 27055
rect 4970 27048 4973 27055
rect 4980 27048 4982 27058
rect 4985 27048 4992 27058
rect 4980 27032 4996 27048
rect 4980 27025 4983 27032
rect 4956 26987 4958 27025
rect 4968 27002 4972 27012
rect 4980 27010 4982 27025
rect 4980 27002 4984 27010
rect 4966 26988 4974 26998
rect 4978 26996 4984 27002
rect 4985 26996 4992 27032
rect 4978 26988 4992 26996
rect 4976 26987 4985 26988
rect 5004 26987 5006 27058
rect 5033 27020 5036 27047
rect 5038 27025 5049 27047
rect 5051 27025 5054 27055
rect 5033 27017 5045 27020
rect 5076 26987 5078 27317
rect 5100 27312 5102 27317
rect 5124 27312 5126 27317
rect 5092 27304 5102 27312
rect 5120 27304 5130 27312
rect 5086 27296 5092 27304
rect 5080 27049 5098 27059
rect 5100 27047 5102 27304
rect 5114 27296 5120 27304
rect 5124 27059 5126 27304
rect 5105 27049 5126 27059
rect 5134 27049 5140 27279
rect 5146 27079 5150 27081
rect 5144 27071 5150 27079
rect 5145 27049 5150 27051
rect 5156 27049 5162 27071
rect 5172 27059 5174 27317
rect 5196 27312 5198 27317
rect 5220 27312 5222 27317
rect 5188 27304 5198 27312
rect 5216 27304 5224 27312
rect 5180 27296 5188 27304
rect 5165 27049 5174 27059
rect 5176 27049 5182 27079
rect 5196 27049 5198 27304
rect 5208 27296 5216 27304
rect 5201 27071 5208 27079
rect 5220 27071 5222 27304
rect 5230 27149 5236 27279
rect 5230 27133 5238 27149
rect 5220 27049 5226 27071
rect 5230 27049 5236 27133
rect 5242 27079 5246 27081
rect 5240 27071 5246 27079
rect 5241 27049 5246 27051
rect 5252 27049 5258 27071
rect 5268 27055 5270 27317
rect 5292 27312 5294 27317
rect 5316 27312 5318 27317
rect 5282 27304 5294 27312
rect 5310 27304 5320 27312
rect 5342 27304 5350 27312
rect 5276 27296 5282 27304
rect 5292 27063 5294 27304
rect 5304 27296 5310 27304
rect 5316 27063 5318 27304
rect 5350 27296 5358 27304
rect 5287 27055 5294 27063
rect 5098 27017 5105 27047
rect 5112 27039 5116 27049
rect 5124 27047 5126 27049
rect 5124 27039 5130 27047
rect 5120 27023 5130 27039
rect 5122 27017 5130 27023
rect 5100 26991 5102 27017
rect 5122 27009 5126 27017
rect 5100 26987 5114 26991
rect 5124 26987 5126 27009
rect 5172 26987 5174 27049
rect 5175 27041 5182 27049
rect 5194 27041 5201 27049
rect 5206 27041 5226 27049
rect 5175 27023 5176 27041
rect 5196 26993 5198 27041
rect 5206 27039 5212 27041
rect 5220 27039 5222 27041
rect 5216 27023 5222 27039
rect 5218 27009 5222 27023
rect 5196 26987 5200 26993
rect 5220 26987 5222 27009
rect 5268 27025 5277 27055
rect 5282 27031 5285 27041
rect 5292 27031 5294 27055
rect 5297 27031 5304 27055
rect 5314 27041 5321 27063
rect 5292 27025 5308 27031
rect 5316 27025 5318 27041
rect 5268 27023 5272 27025
rect 5268 26987 5271 27023
rect 5292 27015 5294 27025
rect 5314 27015 5318 27025
rect 5345 27020 5348 27047
rect 5350 27025 5361 27047
rect 5363 27025 5366 27055
rect 5345 27017 5357 27020
rect 5280 27002 5284 27012
rect 5290 27002 5294 27015
rect 5297 27002 5304 27015
rect 5290 27001 5304 27002
rect 5290 26993 5294 27001
rect 5290 26988 5296 26993
rect 5297 26988 5304 27001
rect 5288 26987 5296 26988
rect 5316 26987 5318 27015
rect 5388 26987 5390 27317
rect 5412 27312 5414 27317
rect 5436 27312 5438 27317
rect 5404 27304 5414 27312
rect 5432 27304 5442 27312
rect 5398 27296 5404 27304
rect 5392 27049 5410 27059
rect 5412 27047 5414 27304
rect 5426 27296 5432 27304
rect 5436 27059 5438 27304
rect 5417 27049 5438 27059
rect 5446 27049 5452 27279
rect 5458 27079 5462 27081
rect 5456 27071 5462 27079
rect 5457 27049 5462 27051
rect 5468 27049 5474 27071
rect 5484 27059 5486 27317
rect 5508 27312 5510 27317
rect 5532 27312 5534 27317
rect 5500 27304 5510 27312
rect 5528 27304 5536 27312
rect 5492 27296 5500 27304
rect 5477 27049 5486 27059
rect 5488 27049 5494 27079
rect 5508 27049 5510 27304
rect 5520 27296 5528 27304
rect 5513 27071 5520 27079
rect 5532 27071 5534 27304
rect 5542 27149 5548 27279
rect 5542 27133 5550 27149
rect 5532 27049 5538 27071
rect 5542 27049 5548 27133
rect 5554 27079 5558 27081
rect 5552 27071 5558 27079
rect 5553 27049 5558 27051
rect 5564 27049 5570 27071
rect 5580 27056 5582 27317
rect 5628 27312 5630 27317
rect 5724 27312 5726 27317
rect 5748 27312 5750 27317
rect 5594 27304 5604 27312
rect 5622 27304 5632 27312
rect 5654 27304 5662 27312
rect 5716 27304 5726 27312
rect 5744 27304 5754 27312
rect 5588 27296 5594 27304
rect 5616 27296 5622 27304
rect 5585 27083 5594 27084
rect 5604 27083 5611 27084
rect 5618 27083 5619 27279
rect 5628 27083 5630 27304
rect 5662 27296 5670 27304
rect 5710 27296 5716 27304
rect 5585 27082 5616 27083
rect 5618 27082 5646 27083
rect 5661 27082 5671 27104
rect 5410 27017 5417 27047
rect 5424 27039 5428 27049
rect 5436 27047 5438 27049
rect 5436 27039 5442 27047
rect 5432 27023 5442 27039
rect 5434 27017 5442 27023
rect 5412 26991 5414 27017
rect 5434 27009 5438 27017
rect 5412 26987 5426 26991
rect 5436 26987 5438 27009
rect 5484 26987 5486 27049
rect 5487 27041 5494 27049
rect 5506 27041 5513 27049
rect 5518 27041 5538 27049
rect 5578 27046 5582 27056
rect 5487 27023 5488 27041
rect 5508 26993 5510 27041
rect 5518 27039 5524 27041
rect 5532 27039 5534 27041
rect 5528 27023 5534 27039
rect 5530 27009 5534 27023
rect 5508 26987 5512 26993
rect 5532 26987 5534 27009
rect 5580 26987 5582 27046
rect 5588 27041 5590 27046
rect 5608 27041 5612 27056
rect 5616 27041 5618 27071
rect 5628 27041 5630 27082
rect 5712 27079 5720 27090
rect 5724 27087 5726 27304
rect 5738 27296 5744 27304
rect 5704 27074 5712 27079
rect 5714 27074 5720 27079
rect 5722 27074 5729 27087
rect 5744 27079 5747 27092
rect 5633 27041 5634 27071
rect 5714 27049 5721 27074
rect 5724 27049 5726 27074
rect 5594 27036 5630 27041
rect 5664 27038 5678 27046
rect 5594 27032 5602 27036
rect 5608 27032 5612 27036
rect 5594 27031 5598 27032
rect 5604 27015 5608 27031
rect 5606 27012 5608 27015
rect 5614 27012 5620 27020
rect 5606 27001 5620 27012
rect 5628 27010 5630 27036
rect 5722 27024 5729 27049
rect 5736 27039 5740 27049
rect 5748 27039 5750 27304
rect 5770 27079 5774 27081
rect 5768 27071 5774 27079
rect 5769 27049 5774 27051
rect 5780 27049 5786 27071
rect 5796 27059 5798 27317
rect 5820 27312 5822 27317
rect 5844 27312 5846 27317
rect 5916 27312 5918 27317
rect 6132 27312 6134 27317
rect 6180 27312 6182 27317
rect 5812 27304 5822 27312
rect 5840 27304 5848 27312
rect 5910 27304 5918 27312
rect 5938 27304 5944 27312
rect 5970 27304 5978 27312
rect 5998 27304 6014 27312
rect 6030 27304 6042 27312
rect 6058 27304 6070 27312
rect 6090 27304 6098 27312
rect 6118 27304 6134 27312
rect 6148 27304 6160 27312
rect 6176 27304 6188 27312
rect 5804 27296 5812 27304
rect 5789 27049 5798 27059
rect 5800 27049 5806 27079
rect 5820 27049 5822 27304
rect 5832 27296 5840 27304
rect 5825 27071 5832 27079
rect 5844 27071 5846 27304
rect 5900 27296 5910 27304
rect 5854 27149 5860 27279
rect 5854 27133 5862 27149
rect 5844 27049 5850 27071
rect 5854 27049 5860 27133
rect 5866 27079 5870 27081
rect 5864 27071 5870 27079
rect 5865 27049 5870 27051
rect 5876 27049 5882 27071
rect 5624 26996 5630 27010
rect 5703 27002 5710 27014
rect 5724 27008 5726 27024
rect 5744 27023 5750 27039
rect 5746 27009 5750 27023
rect 5628 26987 5630 26996
rect 5722 26987 5729 27008
rect 5748 26987 5750 27009
rect 5796 26987 5798 27049
rect 5799 27041 5806 27049
rect 5818 27041 5825 27049
rect 5830 27041 5850 27049
rect 5799 27023 5800 27041
rect 5820 26993 5822 27041
rect 5830 27039 5836 27041
rect 5844 27039 5846 27041
rect 5840 27023 5846 27039
rect 5842 27009 5846 27023
rect 5820 26987 5824 26993
rect 5844 26987 5846 27009
rect 5916 27013 5918 27304
rect 5928 27296 5938 27304
rect 5978 27296 5986 27304
rect 6026 27296 6030 27304
rect 6054 27296 6058 27304
rect 6098 27296 6106 27304
rect 5921 27048 5928 27078
rect 5930 27048 5936 27071
rect 5938 27041 5945 27071
rect 5947 27048 5956 27279
rect 6028 27083 6039 27090
rect 6030 27078 6039 27083
rect 6040 27048 6051 27078
rect 6132 27059 6134 27304
rect 6146 27296 6148 27304
rect 6160 27296 6162 27304
rect 6174 27296 6176 27304
rect 6143 27083 6159 27091
rect 6125 27049 6134 27059
rect 6136 27049 6142 27079
rect 6143 27077 6154 27079
rect 6143 27049 6152 27070
rect 5930 27013 5932 27023
rect 5938 27015 5942 27041
rect 6040 27040 6049 27048
rect 6132 27015 6134 27049
rect 6135 27040 6142 27049
rect 6154 27040 6159 27070
rect 6135 27015 6136 27040
rect 6168 27039 6172 27049
rect 6180 27039 6182 27304
rect 6188 27296 6190 27304
rect 6202 27079 6206 27081
rect 6200 27071 6206 27079
rect 6201 27049 6206 27051
rect 6212 27049 6218 27071
rect 6228 27059 6230 27317
rect 6252 27312 6254 27317
rect 6276 27312 6278 27317
rect 6244 27304 6254 27312
rect 6272 27304 6280 27312
rect 6236 27296 6244 27304
rect 6221 27049 6230 27059
rect 6232 27049 6238 27079
rect 6252 27049 6254 27304
rect 6264 27296 6272 27304
rect 6257 27071 6264 27079
rect 6276 27071 6278 27304
rect 6286 27149 6292 27279
rect 6286 27133 6294 27149
rect 6276 27049 6282 27071
rect 6286 27049 6292 27133
rect 6298 27079 6302 27081
rect 6296 27071 6302 27079
rect 6297 27049 6302 27051
rect 6308 27049 6314 27071
rect 6324 27056 6326 27317
rect 6372 27312 6374 27317
rect 6468 27312 6470 27317
rect 6492 27312 6494 27317
rect 6338 27304 6348 27312
rect 6366 27304 6376 27312
rect 6398 27304 6406 27312
rect 6426 27304 6442 27312
rect 6458 27304 6470 27312
rect 6486 27304 6498 27312
rect 6518 27304 6526 27312
rect 6332 27296 6338 27304
rect 6360 27296 6366 27304
rect 6329 27083 6338 27084
rect 6348 27083 6355 27084
rect 6362 27083 6363 27279
rect 6372 27083 6374 27304
rect 6406 27296 6414 27304
rect 6454 27296 6458 27304
rect 6329 27082 6360 27083
rect 6362 27082 6390 27083
rect 6405 27082 6415 27104
rect 6040 27013 6042 27015
rect 5916 27001 5930 27013
rect 5940 27001 5942 27013
rect 6032 27004 6042 27013
rect 5916 26993 5918 27001
rect 6036 26999 6046 27004
rect 5916 26987 5920 26993
rect 6132 26991 6136 27015
rect 6142 27004 6144 27014
rect 6154 27004 6161 27015
rect 6178 27009 6182 27039
rect 6040 26989 6042 26990
rect 6132 26987 6134 26991
rect 6135 26987 6136 26991
rect 6152 26991 6161 27004
rect 6166 26991 6170 27004
rect 6152 26990 6166 26991
rect 6154 26989 6162 26990
rect 6180 26987 6182 27009
rect 6228 26987 6230 27049
rect 6231 27041 6238 27049
rect 6250 27041 6257 27049
rect 6262 27041 6282 27049
rect 6322 27046 6326 27056
rect 6231 27023 6232 27041
rect 6252 26993 6254 27041
rect 6262 27039 6268 27041
rect 6276 27039 6278 27041
rect 6272 27023 6278 27039
rect 6274 27009 6278 27023
rect 6252 26987 6256 26993
rect 6276 26987 6278 27009
rect 6324 26987 6326 27046
rect 6332 27041 6334 27046
rect 6352 27041 6356 27056
rect 6360 27041 6362 27071
rect 6372 27041 6374 27082
rect 6377 27041 6378 27071
rect 6338 27036 6374 27041
rect 6408 27038 6422 27046
rect 6338 27032 6346 27036
rect 6352 27032 6356 27036
rect 6338 27031 6342 27032
rect 6348 27015 6352 27031
rect 6350 27012 6352 27015
rect 6358 27012 6364 27020
rect 6350 27001 6364 27012
rect 6372 27010 6374 27036
rect 6458 27025 6463 27055
rect 6468 27029 6470 27304
rect 6482 27296 6486 27304
rect 6492 27034 6494 27304
rect 6526 27296 6534 27304
rect 6468 27027 6489 27029
rect 6465 27025 6489 27027
rect 6468 27012 6470 27025
rect 6368 26996 6374 27010
rect 6456 27002 6460 27012
rect 6468 27008 6484 27012
rect 6490 27008 6494 27034
rect 6521 27020 6524 27047
rect 6526 27025 6537 27047
rect 6539 27025 6542 27055
rect 6521 27017 6533 27020
rect 6468 27002 6470 27008
rect 6372 26987 6374 26996
rect 6454 26988 6458 26998
rect 6466 26988 6470 27002
rect 6467 26987 6470 26988
rect 6492 26987 6494 27008
rect 6564 26987 6566 27317
rect 6588 27312 6590 27317
rect 6612 27312 6614 27317
rect 6580 27304 6590 27312
rect 6608 27304 6618 27312
rect 6574 27296 6580 27304
rect 6568 27049 6586 27059
rect 6588 27047 6590 27304
rect 6602 27296 6608 27304
rect 6612 27059 6614 27304
rect 6593 27049 6614 27059
rect 6622 27049 6628 27279
rect 6634 27079 6638 27081
rect 6632 27071 6638 27079
rect 6633 27049 6638 27051
rect 6644 27049 6650 27071
rect 6660 27055 6662 27317
rect 6684 27312 6686 27317
rect 6708 27312 6710 27317
rect 6674 27304 6686 27312
rect 6702 27304 6712 27312
rect 6734 27304 6742 27312
rect 6668 27296 6674 27304
rect 6684 27063 6686 27304
rect 6696 27296 6702 27304
rect 6708 27063 6710 27304
rect 6742 27296 6750 27304
rect 6679 27055 6686 27063
rect 6586 27017 6593 27047
rect 6600 27039 6604 27049
rect 6612 27047 6614 27049
rect 6612 27039 6618 27047
rect 6608 27023 6618 27039
rect 6610 27017 6618 27023
rect 6660 27025 6669 27055
rect 6674 27031 6677 27041
rect 6684 27031 6686 27055
rect 6689 27031 6696 27055
rect 6706 27041 6713 27063
rect 6684 27025 6700 27031
rect 6708 27025 6710 27041
rect 6660 27023 6664 27025
rect 6588 26991 6590 27017
rect 6610 27009 6614 27017
rect 6588 26987 6602 26991
rect 6612 26987 6614 27009
rect 6660 26987 6663 27023
rect 6684 27015 6686 27025
rect 6706 27015 6710 27025
rect 6737 27020 6740 27047
rect 6742 27025 6753 27047
rect 6755 27025 6758 27055
rect 6737 27017 6749 27020
rect 6672 27002 6676 27012
rect 6682 27002 6686 27015
rect 6689 27002 6696 27015
rect 6682 27001 6696 27002
rect 6682 26993 6686 27001
rect 6682 26988 6688 26993
rect 6689 26988 6696 27001
rect 6680 26987 6688 26988
rect 6708 26987 6710 27015
rect 6780 26987 6782 27317
rect 6804 27312 6806 27317
rect 6828 27312 6830 27317
rect 6796 27304 6806 27312
rect 6824 27304 6834 27312
rect 6790 27296 6796 27304
rect 6784 27049 6802 27059
rect 6804 27047 6806 27304
rect 6818 27296 6824 27304
rect 6828 27059 6830 27304
rect 6809 27049 6830 27059
rect 6838 27049 6844 27279
rect 6850 27079 6854 27081
rect 6848 27071 6854 27079
rect 6849 27049 6854 27051
rect 6860 27049 6866 27071
rect 6876 27059 6878 27317
rect 6900 27312 6902 27317
rect 6924 27312 6926 27317
rect 6892 27304 6902 27312
rect 6920 27304 6928 27312
rect 6884 27296 6892 27304
rect 6869 27049 6878 27059
rect 6880 27049 6886 27079
rect 6900 27049 6902 27304
rect 6912 27296 6920 27304
rect 6905 27071 6912 27079
rect 6924 27071 6926 27304
rect 6934 27149 6940 27279
rect 6934 27133 6942 27149
rect 6924 27049 6930 27071
rect 6934 27049 6940 27133
rect 6946 27079 6950 27081
rect 6944 27071 6950 27079
rect 6945 27049 6950 27051
rect 6956 27049 6962 27071
rect 6972 27056 6974 27317
rect 7020 27312 7022 27317
rect 7140 27312 7142 27317
rect 7236 27312 7238 27317
rect 7260 27312 7262 27317
rect 6986 27304 6996 27312
rect 7014 27304 7024 27312
rect 7046 27304 7054 27312
rect 7074 27304 7090 27312
rect 7106 27304 7118 27312
rect 7134 27304 7146 27312
rect 7166 27304 7174 27312
rect 7194 27304 7210 27312
rect 7226 27304 7238 27312
rect 7254 27304 7266 27312
rect 7286 27304 7294 27312
rect 6980 27296 6986 27304
rect 7008 27296 7014 27304
rect 6977 27083 6986 27084
rect 6996 27083 7003 27084
rect 7010 27083 7011 27279
rect 7020 27083 7022 27304
rect 7054 27296 7062 27304
rect 7102 27296 7106 27304
rect 7130 27296 7134 27304
rect 7118 27116 7134 27124
rect 6977 27082 7008 27083
rect 7010 27082 7038 27083
rect 7053 27082 7063 27104
rect 7097 27082 7104 27104
rect 7106 27082 7113 27112
rect 7118 27110 7123 27112
rect 7130 27110 7134 27112
rect 7115 27082 7121 27104
rect 6802 27017 6809 27047
rect 6816 27039 6820 27049
rect 6828 27047 6830 27049
rect 6828 27039 6834 27047
rect 6824 27023 6834 27039
rect 6826 27017 6834 27023
rect 6804 26991 6806 27017
rect 6826 27009 6830 27017
rect 6804 26987 6818 26991
rect 6828 26987 6830 27009
rect 6876 26987 6878 27049
rect 6879 27041 6886 27049
rect 6898 27041 6905 27049
rect 6910 27041 6930 27049
rect 6970 27046 6974 27056
rect 6879 27023 6880 27041
rect 6900 26993 6902 27041
rect 6910 27039 6916 27041
rect 6924 27039 6926 27041
rect 6920 27023 6926 27039
rect 6922 27009 6926 27023
rect 6900 26987 6904 26993
rect 6924 26987 6926 27009
rect 6972 26987 6974 27046
rect 6980 27041 6982 27046
rect 7000 27041 7004 27056
rect 7008 27041 7010 27071
rect 7020 27041 7022 27082
rect 7123 27074 7130 27104
rect 7132 27082 7139 27104
rect 7025 27041 7026 27071
rect 7090 27046 7098 27056
rect 6986 27036 7022 27041
rect 7056 27038 7070 27046
rect 7100 27038 7114 27046
rect 7120 27038 7124 27056
rect 6986 27032 6994 27036
rect 7000 27032 7004 27036
rect 6986 27031 6990 27032
rect 6996 27015 7000 27031
rect 6998 27012 7000 27015
rect 7006 27012 7012 27020
rect 6998 27001 7012 27012
rect 7020 27010 7022 27036
rect 7100 27034 7108 27038
rect 7100 27032 7114 27034
rect 7118 27032 7124 27038
rect 7100 27028 7110 27032
rect 7106 27024 7110 27028
rect 7118 27024 7120 27032
rect 7016 26996 7022 27010
rect 7100 27002 7102 27014
rect 7116 27012 7120 27024
rect 7132 27020 7136 27024
rect 7126 27012 7136 27020
rect 7116 27008 7132 27012
rect 7140 27010 7142 27304
rect 7174 27296 7182 27304
rect 7222 27296 7226 27304
rect 7173 27082 7183 27104
rect 7176 27038 7190 27046
rect 7226 27025 7231 27055
rect 7236 27029 7238 27304
rect 7250 27296 7254 27304
rect 7260 27034 7262 27304
rect 7294 27296 7302 27304
rect 7236 27027 7257 27029
rect 7233 27025 7257 27027
rect 7236 27012 7238 27025
rect 7120 26996 7123 27008
rect 7136 26996 7142 27010
rect 7224 27002 7228 27012
rect 7236 27008 7252 27012
rect 7258 27008 7262 27034
rect 7289 27020 7292 27047
rect 7294 27025 7305 27047
rect 7307 27025 7310 27055
rect 7289 27017 7301 27020
rect 7236 27002 7238 27008
rect 7020 26987 7022 26996
rect 7140 26987 7142 26996
rect 7222 26988 7226 26998
rect 7234 26988 7238 27002
rect 7235 26987 7238 26988
rect 7260 26987 7262 27008
rect 7332 26987 7334 27317
rect 7356 27312 7358 27317
rect 7380 27312 7382 27317
rect 7348 27304 7358 27312
rect 7376 27304 7386 27312
rect 7342 27296 7348 27304
rect 7336 27049 7354 27059
rect 7356 27047 7358 27304
rect 7370 27296 7376 27304
rect 7380 27059 7382 27304
rect 7361 27049 7382 27059
rect 7390 27049 7396 27279
rect 7402 27079 7406 27081
rect 7400 27071 7406 27079
rect 7401 27049 7406 27051
rect 7412 27049 7418 27071
rect 7428 27059 7430 27317
rect 7452 27312 7454 27317
rect 7476 27312 7478 27317
rect 7444 27304 7454 27312
rect 7472 27304 7480 27312
rect 7436 27296 7444 27304
rect 7421 27049 7430 27059
rect 7432 27049 7438 27079
rect 7452 27049 7454 27304
rect 7464 27296 7472 27304
rect 7457 27071 7464 27079
rect 7476 27071 7478 27304
rect 7486 27149 7492 27279
rect 7486 27133 7494 27149
rect 7476 27049 7482 27071
rect 7486 27049 7492 27133
rect 7498 27079 7502 27081
rect 7496 27071 7502 27079
rect 7497 27049 7502 27051
rect 7508 27049 7514 27071
rect 7524 27059 7526 27317
rect 7548 27312 7550 27317
rect 7572 27312 7574 27317
rect 7540 27304 7550 27312
rect 7568 27304 7576 27312
rect 7532 27296 7540 27304
rect 7517 27049 7526 27059
rect 7528 27049 7534 27079
rect 7548 27049 7550 27304
rect 7560 27296 7568 27304
rect 7553 27071 7560 27079
rect 7572 27071 7574 27304
rect 7582 27149 7588 27279
rect 7582 27133 7590 27149
rect 7572 27049 7578 27071
rect 7582 27049 7588 27133
rect 7594 27079 7598 27081
rect 7592 27071 7598 27079
rect 7593 27049 7598 27051
rect 7604 27049 7610 27071
rect 7620 27059 7622 27317
rect 7644 27312 7646 27317
rect 7668 27312 7670 27317
rect 7636 27304 7646 27312
rect 7664 27304 7672 27312
rect 7628 27296 7636 27304
rect 7613 27049 7622 27059
rect 7624 27049 7630 27079
rect 7644 27049 7646 27304
rect 7656 27296 7664 27304
rect 7649 27071 7656 27079
rect 7668 27071 7670 27304
rect 7678 27149 7684 27279
rect 7678 27133 7686 27149
rect 7668 27049 7674 27071
rect 7678 27049 7684 27133
rect 7690 27079 7694 27081
rect 7688 27071 7694 27079
rect 7689 27049 7694 27051
rect 7700 27049 7706 27071
rect 7716 27055 7718 27317
rect 7740 27312 7742 27317
rect 7764 27312 7766 27317
rect 7730 27304 7742 27312
rect 7758 27304 7768 27312
rect 7790 27304 7798 27312
rect 7724 27296 7730 27304
rect 7740 27063 7742 27304
rect 7752 27296 7758 27304
rect 7764 27063 7766 27304
rect 7798 27296 7806 27304
rect 7735 27055 7742 27063
rect 7354 27017 7361 27047
rect 7368 27039 7372 27049
rect 7380 27047 7382 27049
rect 7380 27039 7386 27047
rect 7376 27023 7386 27039
rect 7378 27017 7386 27023
rect 7356 26991 7358 27017
rect 7378 27009 7382 27017
rect 7356 26987 7370 26991
rect 7380 26987 7382 27009
rect 7428 26987 7430 27049
rect 7431 27041 7438 27049
rect 7450 27041 7457 27049
rect 7462 27041 7482 27049
rect 7431 27023 7432 27041
rect 7452 26993 7454 27041
rect 7462 27039 7468 27041
rect 7476 27039 7478 27041
rect 7472 27023 7478 27039
rect 7474 27009 7478 27023
rect 7452 26987 7456 26993
rect 7476 26987 7478 27009
rect 7524 26987 7526 27049
rect 7527 27041 7534 27049
rect 7546 27041 7553 27049
rect 7558 27041 7578 27049
rect 7527 27023 7528 27041
rect 7548 26993 7550 27041
rect 7558 27039 7564 27041
rect 7572 27039 7574 27041
rect 7568 27023 7574 27039
rect 7570 27009 7574 27023
rect 7548 26987 7552 26993
rect 7572 26987 7574 27009
rect 7620 26987 7622 27049
rect 7623 27041 7630 27049
rect 7642 27041 7649 27049
rect 7654 27041 7674 27049
rect 7623 27023 7624 27041
rect 7644 26993 7646 27041
rect 7654 27039 7660 27041
rect 7668 27039 7670 27041
rect 7664 27023 7670 27039
rect 7666 27009 7670 27023
rect 7644 26987 7648 26993
rect 7668 26987 7670 27009
rect 7716 27025 7725 27055
rect 7730 27031 7733 27041
rect 7740 27031 7742 27055
rect 7745 27031 7752 27055
rect 7762 27041 7769 27063
rect 7740 27025 7756 27031
rect 7764 27025 7766 27041
rect 7716 27023 7720 27025
rect 7716 26987 7719 27023
rect 7740 27015 7742 27025
rect 7762 27015 7766 27025
rect 7793 27020 7796 27047
rect 7798 27025 7809 27047
rect 7811 27025 7814 27055
rect 7793 27017 7805 27020
rect 7728 27002 7732 27012
rect 7738 27002 7742 27015
rect 7745 27002 7752 27015
rect 7738 27001 7752 27002
rect 7738 26993 7742 27001
rect 7738 26988 7744 26993
rect 7745 26988 7752 27001
rect 7736 26987 7744 26988
rect 7764 26987 7766 27015
rect 7836 26987 7838 27317
rect 7860 27312 7862 27317
rect 7884 27312 7886 27317
rect 7852 27304 7862 27312
rect 7880 27304 7890 27312
rect 7846 27296 7852 27304
rect 7840 27049 7858 27059
rect 7860 27047 7862 27304
rect 7874 27296 7880 27304
rect 7884 27059 7886 27304
rect 7865 27049 7886 27059
rect 7894 27049 7900 27279
rect 7906 27079 7910 27081
rect 7904 27071 7910 27079
rect 7905 27049 7910 27051
rect 7916 27049 7922 27071
rect 7932 27059 7934 27317
rect 7956 27312 7958 27317
rect 7980 27312 7982 27317
rect 8052 27312 8054 27317
rect 8148 27312 8150 27317
rect 8196 27312 8198 27317
rect 7948 27304 7958 27312
rect 7976 27304 7984 27312
rect 8046 27304 8054 27312
rect 8074 27304 8080 27312
rect 8106 27304 8114 27312
rect 8134 27304 8150 27312
rect 8164 27304 8176 27312
rect 8192 27304 8204 27312
rect 7940 27296 7948 27304
rect 7925 27049 7934 27059
rect 7936 27049 7942 27079
rect 7956 27049 7958 27304
rect 7968 27296 7976 27304
rect 7961 27071 7968 27079
rect 7980 27071 7982 27304
rect 8036 27296 8046 27304
rect 7990 27149 7996 27279
rect 7990 27133 7998 27149
rect 7980 27049 7986 27071
rect 7990 27049 7996 27133
rect 8002 27079 8006 27081
rect 8000 27071 8006 27079
rect 8001 27049 8006 27051
rect 8012 27049 8018 27071
rect 7858 27017 7865 27047
rect 7872 27039 7876 27049
rect 7884 27047 7886 27049
rect 7884 27039 7890 27047
rect 7880 27023 7890 27039
rect 7882 27017 7890 27023
rect 7860 26991 7862 27017
rect 7882 27009 7886 27017
rect 7860 26987 7874 26991
rect 7884 26987 7886 27009
rect 7932 26987 7934 27049
rect 7935 27041 7942 27049
rect 7954 27041 7961 27049
rect 7966 27041 7986 27049
rect 7935 27023 7936 27041
rect 7956 26993 7958 27041
rect 7966 27039 7972 27041
rect 7980 27039 7982 27041
rect 7976 27023 7982 27039
rect 7978 27009 7982 27023
rect 7956 26987 7960 26993
rect 7980 26987 7982 27009
rect 8052 27013 8054 27304
rect 8064 27296 8074 27304
rect 8114 27296 8122 27304
rect 8057 27048 8064 27078
rect 8066 27048 8072 27071
rect 8074 27041 8081 27071
rect 8083 27048 8092 27279
rect 8148 27059 8150 27304
rect 8162 27296 8164 27304
rect 8176 27296 8178 27304
rect 8190 27296 8192 27304
rect 8159 27083 8175 27091
rect 8141 27049 8150 27059
rect 8152 27049 8158 27079
rect 8159 27077 8170 27079
rect 8159 27049 8168 27070
rect 8066 27013 8068 27023
rect 8074 27015 8078 27041
rect 8148 27015 8150 27049
rect 8151 27040 8158 27049
rect 8170 27040 8175 27070
rect 8151 27015 8152 27040
rect 8184 27039 8188 27049
rect 8196 27039 8198 27304
rect 8204 27296 8206 27304
rect 8218 27079 8222 27081
rect 8216 27071 8222 27079
rect 8217 27049 8222 27051
rect 8228 27049 8234 27071
rect 8244 27059 8246 27317
rect 8268 27312 8270 27317
rect 8292 27312 8294 27317
rect 8260 27304 8270 27312
rect 8288 27304 8296 27312
rect 8252 27296 8260 27304
rect 8237 27049 8246 27059
rect 8248 27049 8254 27079
rect 8268 27049 8270 27304
rect 8280 27296 8288 27304
rect 8273 27071 8280 27079
rect 8292 27071 8294 27304
rect 8302 27149 8308 27279
rect 8302 27133 8310 27149
rect 8292 27049 8298 27071
rect 8302 27049 8308 27133
rect 8314 27079 8318 27081
rect 8312 27071 8318 27079
rect 8313 27049 8318 27051
rect 8324 27049 8330 27071
rect 8340 27059 8342 27317
rect 8364 27312 8366 27317
rect 8388 27312 8390 27317
rect 8356 27304 8366 27312
rect 8384 27304 8392 27312
rect 8348 27296 8356 27304
rect 8333 27049 8342 27059
rect 8344 27049 8350 27079
rect 8364 27049 8366 27304
rect 8376 27296 8384 27304
rect 8369 27071 8376 27079
rect 8388 27071 8390 27304
rect 8398 27149 8404 27279
rect 8398 27133 8406 27149
rect 8388 27049 8394 27071
rect 8398 27049 8404 27133
rect 8410 27079 8414 27081
rect 8408 27071 8414 27079
rect 8409 27049 8414 27051
rect 8420 27049 8426 27071
rect 8436 27055 8438 27317
rect 8460 27312 8462 27317
rect 8484 27312 8486 27317
rect 8450 27304 8462 27312
rect 8478 27304 8488 27312
rect 8510 27304 8518 27312
rect 8538 27304 8554 27312
rect 8444 27296 8450 27304
rect 8460 27063 8462 27304
rect 8472 27296 8478 27304
rect 8484 27063 8486 27304
rect 8518 27296 8526 27304
rect 8455 27055 8462 27063
rect 8052 27001 8066 27013
rect 8076 27001 8078 27013
rect 8052 26993 8054 27001
rect 8052 26987 8056 26993
rect 8148 26991 8152 27015
rect 8158 27004 8160 27014
rect 8170 27004 8177 27015
rect 8194 27009 8198 27039
rect 8148 26987 8150 26991
rect 8151 26987 8152 26991
rect 8168 26991 8177 27004
rect 8182 26991 8186 27004
rect 8168 26990 8182 26991
rect 8170 26989 8178 26990
rect 8196 26987 8198 27009
rect 8244 26987 8246 27049
rect 8247 27041 8254 27049
rect 8266 27041 8273 27049
rect 8278 27041 8298 27049
rect 8247 27023 8248 27041
rect 8268 26993 8270 27041
rect 8278 27039 8284 27041
rect 8292 27039 8294 27041
rect 8288 27023 8294 27039
rect 8290 27009 8294 27023
rect 8268 26987 8272 26993
rect 8292 26987 8294 27009
rect 8340 26987 8342 27049
rect 8343 27041 8350 27049
rect 8362 27041 8369 27049
rect 8374 27041 8394 27049
rect 8343 27023 8344 27041
rect 8364 26993 8366 27041
rect 8374 27039 8380 27041
rect 8388 27039 8390 27041
rect 8384 27023 8390 27039
rect 8386 27009 8390 27023
rect 8364 26987 8368 26993
rect 8388 26987 8390 27009
rect 8436 27025 8445 27055
rect 8450 27031 8453 27041
rect 8460 27031 8462 27055
rect 8465 27031 8472 27055
rect 8482 27041 8489 27063
rect 8556 27055 8558 27317
rect 8580 27312 8582 27317
rect 8604 27312 8606 27317
rect 8570 27304 8582 27312
rect 8598 27304 8610 27312
rect 8630 27304 8638 27312
rect 8658 27304 8672 27312
rect 8566 27296 8570 27304
rect 8460 27025 8476 27031
rect 8484 27025 8486 27041
rect 8436 27023 8440 27025
rect 8436 26987 8439 27023
rect 8460 27015 8462 27025
rect 8482 27015 8486 27025
rect 8513 27020 8516 27047
rect 8518 27025 8529 27047
rect 8531 27025 8534 27055
rect 8556 27025 8565 27055
rect 8580 27025 8582 27304
rect 8594 27296 8598 27304
rect 8585 27025 8592 27055
rect 8604 27047 8606 27304
rect 8638 27296 8646 27304
rect 8672 27296 8674 27304
rect 8664 27096 8668 27106
rect 8676 27096 8678 27317
rect 8700 27312 8702 27317
rect 8724 27312 8726 27317
rect 8688 27304 8702 27312
rect 8716 27304 8728 27312
rect 8748 27304 8756 27312
rect 8686 27296 8688 27304
rect 8674 27066 8678 27096
rect 8513 27017 8525 27020
rect 8448 27002 8452 27012
rect 8458 27002 8462 27015
rect 8465 27002 8472 27015
rect 8458 27001 8472 27002
rect 8458 26993 8462 27001
rect 8458 26988 8464 26993
rect 8465 26988 8472 27001
rect 8456 26987 8464 26988
rect 8484 26987 8486 27015
rect 8556 26987 8558 27025
rect 8575 27017 8582 27025
rect 8602 27017 8609 27047
rect 8633 27020 8636 27047
rect 8638 27025 8649 27047
rect 8651 27025 8654 27055
rect 8633 27017 8645 27020
rect 8568 27002 8572 27012
rect 8580 27002 8582 27017
rect 8585 27007 8592 27017
rect 8578 26988 8592 27002
rect 8602 26991 8606 27017
rect 8676 27004 8678 27066
rect 8692 27055 8699 27065
rect 8692 27047 8695 27055
rect 8692 27020 8699 27047
rect 8688 27017 8699 27020
rect 8688 27010 8695 27017
rect 8700 27010 8702 27304
rect 8714 27296 8716 27304
rect 8724 27104 8726 27304
rect 8728 27296 8730 27304
rect 8756 27296 8764 27304
rect 8719 27096 8726 27104
rect 8772 27096 8774 27317
rect 8820 27312 8822 27317
rect 8844 27312 8846 27317
rect 8868 27312 8870 27317
rect 9333 27314 9349 27317
rect 8776 27304 8784 27312
rect 8804 27304 8822 27312
rect 8836 27304 8848 27312
rect 8864 27304 8876 27312
rect 8931 27304 8940 27312
rect 8960 27304 8968 27312
rect 8991 27304 9001 27312
rect 9020 27304 9029 27312
rect 9049 27304 9057 27312
rect 9077 27304 9085 27312
rect 9105 27304 9114 27312
rect 9133 27304 9142 27312
rect 9162 27304 9170 27312
rect 9190 27304 9198 27312
rect 9218 27304 9226 27312
rect 9246 27304 9254 27312
rect 9274 27304 9282 27312
rect 9302 27304 9310 27312
rect 9496 27309 9498 27317
rect 9358 27304 9366 27309
rect 9386 27304 9394 27309
rect 8784 27296 8792 27304
rect 8714 27095 8730 27096
rect 8705 27047 8709 27055
rect 8712 27051 8716 27061
rect 8719 27051 8722 27065
rect 8724 27051 8726 27095
rect 8768 27088 8774 27096
rect 8750 27058 8753 27088
rect 8772 27066 8775 27088
rect 8795 27066 8798 27096
rect 8758 27059 8766 27066
rect 8772 27059 8774 27066
rect 8775 27061 8780 27066
rect 8775 27059 8789 27061
rect 8758 27058 8789 27059
rect 8758 27056 8759 27058
rect 8760 27056 8764 27058
rect 8772 27056 8774 27058
rect 8719 27047 8726 27051
rect 8719 27021 8730 27047
rect 8768 27040 8769 27056
rect 8770 27026 8774 27056
rect 8719 27020 8726 27021
rect 8579 26987 8592 26988
rect 8604 26987 8606 26991
rect 8673 26987 8678 27004
rect 8692 26987 8695 27010
rect 8698 27007 8702 27010
rect 8705 27007 8710 27020
rect 8714 27017 8726 27020
rect 8698 26996 8712 27007
rect 8700 26987 8709 26996
rect 8719 26991 8726 27017
rect 8772 27004 8774 27026
rect 8719 26987 8722 26991
rect 8724 26987 8726 26991
rect 8759 26994 8762 26998
rect 8759 26988 8763 26994
rect 8768 26987 8774 27004
rect 8820 26987 8822 27304
rect 8832 27296 8836 27304
rect 8844 27087 8846 27304
rect 8860 27296 8864 27304
rect 8868 27087 8870 27304
rect 8924 27296 8931 27304
rect 8952 27296 8960 27304
rect 9001 27296 9007 27304
rect 9029 27296 9036 27304
rect 9057 27296 9065 27304
rect 9085 27296 9093 27304
rect 9114 27296 9121 27304
rect 9142 27296 9149 27304
rect 9170 27296 9178 27304
rect 9198 27296 9206 27304
rect 9226 27296 9234 27304
rect 9254 27296 9262 27304
rect 9282 27296 9290 27304
rect 9310 27296 9318 27304
rect 9366 27293 9374 27304
rect 9394 27294 9402 27304
rect 9442 27301 9450 27309
rect 9470 27301 9478 27309
rect 9496 27301 9506 27309
rect 9526 27301 9538 27312
rect 9554 27301 9566 27312
rect 9582 27301 9594 27312
rect 9614 27304 9622 27312
rect 9450 27294 9458 27301
rect 9478 27294 9486 27301
rect 9386 27293 9402 27294
rect 9442 27293 9458 27294
rect 9470 27293 9486 27294
rect 9496 27294 9498 27301
rect 9506 27294 9514 27301
rect 9538 27296 9542 27301
rect 9566 27296 9570 27301
rect 9594 27296 9598 27301
rect 9622 27296 9630 27304
rect 9496 27293 9514 27294
rect 9526 27293 9534 27294
rect 9046 27279 9179 27287
rect 9184 27279 9237 27287
rect 8878 27146 8884 27279
rect 9194 27261 9198 27270
rect 9262 27269 9269 27278
rect 9245 27257 9251 27262
rect 9270 27257 9279 27269
rect 9241 27252 9245 27257
rect 9270 27253 9286 27257
rect 9287 27253 9290 27257
rect 8878 27133 8886 27146
rect 8842 27079 8849 27087
rect 8824 27049 8829 27079
rect 8834 27049 8840 27058
rect 8844 27051 8846 27079
rect 8868 27058 8874 27087
rect 8878 27058 8884 27133
rect 8890 27079 8894 27081
rect 8954 27080 8960 27248
rect 9019 27238 9025 27246
rect 9056 27238 9067 27242
rect 9029 27230 9035 27238
rect 9010 27210 9025 27230
rect 9056 27227 9069 27238
rect 9094 27230 9101 27238
rect 9085 27227 9101 27230
rect 9132 27227 9142 27249
rect 9010 27200 9029 27210
rect 9036 27200 9055 27210
rect 9029 27198 9035 27200
rect 9076 27198 9079 27227
rect 9085 27208 9093 27227
rect 9159 27219 9165 27249
rect 9200 27219 9205 27249
rect 9241 27227 9242 27252
rect 9274 27227 9281 27253
rect 9081 27200 9094 27208
rect 9029 27192 9036 27198
rect 9029 27190 9043 27192
rect 9029 27185 9052 27190
rect 9018 27160 9025 27170
rect 9036 27168 9052 27185
rect 9062 27168 9069 27198
rect 9083 27195 9101 27198
rect 9076 27166 9083 27190
rect 9091 27168 9101 27195
rect 9274 27193 9279 27227
rect 9311 27221 9320 27222
rect 9317 27219 9320 27221
rect 9152 27190 9158 27193
rect 9036 27160 9090 27166
rect 9091 27160 9100 27168
rect 9117 27163 9133 27190
rect 9152 27163 9155 27190
rect 9158 27163 9159 27190
rect 9193 27185 9198 27193
rect 9193 27163 9209 27185
rect 9215 27163 9223 27185
rect 9117 27160 9124 27163
rect 9159 27160 9165 27163
rect 9026 27153 9035 27160
rect 9193 27155 9231 27163
rect 9262 27155 9269 27185
rect 9274 27163 9281 27193
rect 9496 27186 9498 27293
rect 9283 27163 9290 27185
rect 9295 27163 9299 27185
rect 9283 27155 9300 27163
rect 9384 27156 9396 27172
rect 8964 27125 8970 27130
rect 8888 27071 8894 27079
rect 8849 27053 8856 27058
rect 8849 27051 8865 27053
rect 8841 27049 8865 27051
rect 8844 27010 8846 27049
rect 8854 27039 8860 27049
rect 8868 27039 8870 27058
rect 8889 27049 8894 27051
rect 8900 27049 8906 27071
rect 8952 27041 8957 27071
rect 9026 27070 9033 27153
rect 9076 27122 9079 27133
rect 9158 27132 9165 27148
rect 9167 27133 9197 27140
rect 9274 27130 9279 27155
rect 9475 27148 9476 27164
rect 9491 27162 9499 27186
rect 9290 27133 9304 27140
rect 9076 27092 9083 27122
rect 9193 27100 9198 27130
rect 9234 27100 9241 27130
rect 9262 27100 9263 27122
rect 9274 27100 9281 27130
rect 9247 27092 9269 27100
rect 9295 27092 9302 27122
rect 9353 27106 9366 27122
rect 9371 27106 9375 27136
rect 9453 27110 9469 27126
rect 9462 27101 9469 27110
rect 9474 27106 9476 27128
rect 9491 27106 9500 27146
rect 9445 27098 9449 27101
rect 9460 27098 9476 27101
rect 9076 27070 9079 27092
rect 9274 27083 9279 27092
rect 9010 27062 9062 27070
rect 9069 27062 9081 27070
rect 9125 27062 9161 27070
rect 8864 27023 8870 27039
rect 8834 26991 8838 27000
rect 8844 26996 8848 27010
rect 8866 27009 8870 27023
rect 8842 26987 8849 26996
rect 8868 26987 8870 27009
rect 9026 26987 9033 27062
rect 9076 27060 9079 27062
rect 9062 27052 9069 27060
rect 9062 27030 9078 27052
rect 9094 27030 9101 27060
rect 9152 27052 9158 27060
rect 9193 27052 9198 27060
rect 9274 27057 9281 27083
rect 9274 27052 9279 27057
rect 9135 27030 9147 27052
rect 9152 27030 9153 27052
rect 9158 27030 9159 27052
rect 9198 27030 9200 27052
rect 9211 27030 9226 27052
rect 9159 27027 9165 27030
rect 9131 27022 9165 27027
rect 9200 27022 9205 27030
rect 9262 27022 9269 27052
rect 9295 27026 9302 27052
rect 9304 27047 9312 27082
rect 9383 27027 9387 27043
rect 9388 27041 9399 27043
rect 9435 27041 9441 27098
rect 9454 27071 9455 27073
rect 9462 27071 9468 27098
rect 9511 27083 9514 27091
rect 9521 27081 9524 27083
rect 9451 27041 9458 27071
rect 9464 27041 9469 27063
rect 9474 27041 9480 27063
rect 9482 27041 9489 27071
rect 9491 27041 9500 27081
rect 9501 27041 9507 27063
rect 9509 27041 9516 27071
rect 9521 27041 9527 27081
rect 9530 27055 9531 27065
rect 9398 27035 9399 27041
rect 9462 27033 9469 27041
rect 9491 27033 9499 27041
rect 9286 27022 9302 27026
rect 9076 26987 9079 27022
rect 9147 26999 9151 27015
rect 9152 26987 9155 26995
rect 9211 26991 9227 26993
rect 9274 26987 9279 27022
rect 9462 27018 9468 27033
rect 9361 27008 9369 27018
rect 9462 27013 9477 27018
rect 9371 27008 9380 27011
rect 9371 26992 9379 27008
rect 9380 26995 9387 27008
rect 9462 27003 9468 27013
rect 9492 26987 9499 27033
rect 9540 27025 9545 27055
rect 9550 27033 9557 27055
rect 9559 27033 9566 27063
rect 9586 27033 9593 27063
rect 9540 27013 9541 27025
rect 9553 27000 9560 27025
rect 9550 26990 9562 26998
rect 9568 26988 9575 27033
rect 9617 27020 9620 27047
rect 9622 27025 9633 27047
rect 9635 27025 9638 27055
rect 9617 27017 9629 27020
rect 9660 26987 9662 27317
rect 9684 27312 9686 27317
rect 9708 27312 9710 27317
rect 9676 27304 9686 27312
rect 9704 27304 9714 27312
rect 9670 27296 9676 27304
rect 9664 27049 9682 27059
rect 9684 27047 9686 27304
rect 9698 27296 9704 27304
rect 9708 27059 9710 27304
rect 9689 27049 9710 27059
rect 9718 27049 9724 27279
rect 9730 27079 9734 27081
rect 9728 27071 9734 27079
rect 9729 27049 9734 27051
rect 9740 27049 9746 27071
rect 9756 27059 9758 27317
rect 9780 27312 9782 27317
rect 9804 27312 9806 27317
rect 9772 27304 9782 27312
rect 9800 27304 9808 27312
rect 9764 27296 9772 27304
rect 9749 27049 9758 27059
rect 9760 27049 9766 27079
rect 9780 27049 9782 27304
rect 9792 27296 9800 27304
rect 9785 27071 9792 27079
rect 9804 27071 9806 27304
rect 9814 27149 9820 27279
rect 9814 27133 9822 27149
rect 9804 27049 9810 27071
rect 9814 27049 9820 27133
rect 9826 27079 9830 27081
rect 9824 27071 9830 27079
rect 9825 27049 9830 27051
rect 9836 27049 9842 27071
rect 9852 27059 9854 27317
rect 9876 27312 9878 27317
rect 9900 27312 9902 27317
rect 9868 27304 9878 27312
rect 9896 27304 9904 27312
rect 9860 27296 9868 27304
rect 9845 27049 9854 27059
rect 9856 27049 9862 27079
rect 9876 27049 9878 27304
rect 9888 27296 9896 27304
rect 9881 27071 9888 27079
rect 9900 27071 9902 27304
rect 9910 27149 9916 27279
rect 9910 27133 9918 27149
rect 9900 27049 9906 27071
rect 9910 27049 9916 27133
rect 9922 27079 9926 27081
rect 9920 27071 9926 27079
rect 9921 27049 9926 27051
rect 9932 27049 9938 27071
rect 9948 27055 9950 27317
rect 9972 27312 9974 27317
rect 9996 27312 9998 27317
rect 9962 27304 9974 27312
rect 9990 27304 10000 27312
rect 10022 27304 10030 27312
rect 9956 27296 9962 27304
rect 9972 27063 9974 27304
rect 9984 27296 9990 27304
rect 9996 27063 9998 27304
rect 10030 27296 10038 27304
rect 9967 27055 9974 27063
rect 9682 27017 9689 27047
rect 9696 27039 9700 27049
rect 9708 27047 9710 27049
rect 9708 27039 9714 27047
rect 9704 27023 9714 27039
rect 9706 27017 9714 27023
rect 9684 26991 9686 27017
rect 9706 27009 9710 27017
rect 9684 26987 9698 26991
rect 9708 26987 9710 27009
rect 9756 26987 9758 27049
rect 9759 27041 9766 27049
rect 9778 27041 9785 27049
rect 9790 27041 9810 27049
rect 9759 27023 9760 27041
rect 9780 26993 9782 27041
rect 9790 27039 9796 27041
rect 9804 27039 9806 27041
rect 9800 27023 9806 27039
rect 9802 27009 9806 27023
rect 9780 26987 9784 26993
rect 9804 26987 9806 27009
rect 9852 26987 9854 27049
rect 9855 27041 9862 27049
rect 9874 27041 9881 27049
rect 9886 27041 9906 27049
rect 9855 27023 9856 27041
rect 9876 26993 9878 27041
rect 9886 27039 9892 27041
rect 9900 27039 9902 27041
rect 9896 27023 9902 27039
rect 9898 27009 9902 27023
rect 9876 26987 9880 26993
rect 9900 26987 9902 27009
rect 9948 27025 9957 27055
rect 9962 27031 9965 27041
rect 9972 27031 9974 27055
rect 9977 27031 9984 27055
rect 9994 27041 10001 27063
rect 9972 27025 9988 27031
rect 9996 27025 9998 27041
rect 9948 27023 9952 27025
rect 9948 26987 9951 27023
rect 9972 27015 9974 27025
rect 9994 27015 9998 27025
rect 10025 27020 10028 27047
rect 10030 27025 10041 27047
rect 10043 27025 10046 27055
rect 10025 27017 10037 27020
rect 9960 27002 9964 27012
rect 9970 27002 9974 27015
rect 9977 27002 9984 27015
rect 9970 27001 9984 27002
rect 9970 26993 9974 27001
rect 9970 26988 9976 26993
rect 9977 26988 9984 27001
rect 9968 26987 9976 26988
rect 9996 26987 9998 27015
rect 10068 26987 10070 27317
rect 10092 27312 10094 27317
rect 10116 27312 10118 27317
rect 10084 27304 10094 27312
rect 10112 27304 10122 27312
rect 10078 27296 10084 27304
rect 10072 27049 10090 27059
rect 10092 27047 10094 27304
rect 10106 27296 10112 27304
rect 10116 27059 10118 27304
rect 10097 27049 10118 27059
rect 10126 27049 10132 27279
rect 10138 27079 10142 27081
rect 10136 27071 10142 27079
rect 10137 27049 10142 27051
rect 10148 27049 10154 27071
rect 10164 27059 10166 27317
rect 10188 27312 10190 27317
rect 10212 27312 10214 27317
rect 10180 27304 10190 27312
rect 10208 27304 10216 27312
rect 10172 27296 10180 27304
rect 10157 27049 10166 27059
rect 10168 27049 10174 27079
rect 10188 27049 10190 27304
rect 10200 27296 10208 27304
rect 10193 27071 10200 27079
rect 10212 27071 10214 27304
rect 10222 27149 10228 27279
rect 10222 27133 10230 27149
rect 10212 27049 10218 27071
rect 10222 27049 10228 27133
rect 10234 27079 10238 27081
rect 10232 27071 10238 27079
rect 10233 27049 10238 27051
rect 10244 27049 10250 27071
rect 10260 27055 10262 27317
rect 10284 27312 10286 27317
rect 10308 27312 10310 27317
rect 10274 27304 10286 27312
rect 10302 27304 10312 27312
rect 10334 27304 10342 27312
rect 10268 27296 10274 27304
rect 10284 27063 10286 27304
rect 10296 27296 10302 27304
rect 10308 27063 10310 27304
rect 10342 27296 10350 27304
rect 10279 27055 10286 27063
rect 10090 27017 10097 27047
rect 10104 27039 10108 27049
rect 10116 27047 10118 27049
rect 10116 27039 10122 27047
rect 10112 27023 10122 27039
rect 10114 27017 10122 27023
rect 10092 26991 10094 27017
rect 10114 27009 10118 27017
rect 10092 26987 10106 26991
rect 10116 26987 10118 27009
rect 10164 26987 10166 27049
rect 10167 27041 10174 27049
rect 10186 27041 10193 27049
rect 10198 27041 10218 27049
rect 10167 27023 10168 27041
rect 10188 26993 10190 27041
rect 10198 27039 10204 27041
rect 10212 27039 10214 27041
rect 10208 27023 10214 27039
rect 10210 27009 10214 27023
rect 10188 26987 10192 26993
rect 10212 26987 10214 27009
rect 10260 27025 10269 27055
rect 10274 27031 10277 27041
rect 10284 27031 10286 27055
rect 10289 27031 10296 27055
rect 10306 27041 10313 27063
rect 10284 27025 10300 27031
rect 10308 27025 10310 27041
rect 10260 27023 10264 27025
rect 10260 26987 10263 27023
rect 10284 27015 10286 27025
rect 10306 27015 10310 27025
rect 10337 27020 10340 27047
rect 10342 27025 10353 27047
rect 10355 27025 10358 27055
rect 10337 27017 10349 27020
rect 10272 27002 10276 27012
rect 10282 27002 10286 27015
rect 10289 27002 10296 27015
rect 10282 27001 10296 27002
rect 10282 26993 10286 27001
rect 10282 26988 10288 26993
rect 10289 26988 10296 27001
rect 10280 26987 10288 26988
rect 10308 26987 10310 27015
rect 10380 26987 10382 27317
rect 10404 27312 10406 27317
rect 10428 27312 10430 27317
rect 10396 27304 10406 27312
rect 10424 27304 10434 27312
rect 10390 27296 10396 27304
rect 10384 27049 10402 27059
rect 10404 27047 10406 27304
rect 10418 27296 10424 27304
rect 10428 27059 10430 27304
rect 10409 27049 10430 27059
rect 10438 27049 10444 27279
rect 10450 27079 10454 27081
rect 10448 27071 10454 27079
rect 10449 27049 10454 27051
rect 10460 27049 10466 27071
rect 10476 27059 10478 27317
rect 10500 27312 10502 27317
rect 10524 27312 10526 27317
rect 10492 27304 10502 27312
rect 10520 27304 10528 27312
rect 10484 27296 10492 27304
rect 10469 27049 10478 27059
rect 10480 27049 10486 27079
rect 10500 27049 10502 27304
rect 10512 27296 10520 27304
rect 10505 27071 10512 27079
rect 10524 27071 10526 27304
rect 10534 27149 10540 27279
rect 10534 27133 10542 27149
rect 10524 27049 10530 27071
rect 10534 27049 10540 27133
rect 10546 27079 10550 27081
rect 10544 27071 10550 27079
rect 10545 27049 10550 27051
rect 10556 27049 10562 27071
rect 10572 27059 10574 27317
rect 10596 27312 10598 27317
rect 10620 27312 10622 27317
rect 10588 27304 10598 27312
rect 10616 27304 10624 27312
rect 10580 27296 10588 27304
rect 10565 27049 10574 27059
rect 10576 27049 10582 27079
rect 10596 27049 10598 27304
rect 10608 27296 10616 27304
rect 10601 27071 10608 27079
rect 10620 27071 10622 27304
rect 10630 27149 10636 27279
rect 10630 27133 10638 27149
rect 10620 27049 10626 27071
rect 10630 27049 10636 27133
rect 10642 27079 10646 27081
rect 10640 27071 10646 27079
rect 10641 27049 10646 27051
rect 10652 27049 10658 27071
rect 10668 27055 10670 27317
rect 10692 27312 10694 27317
rect 10716 27312 10718 27317
rect 10682 27304 10694 27312
rect 10710 27304 10720 27312
rect 10742 27304 10750 27312
rect 10770 27304 10786 27312
rect 10676 27296 10682 27304
rect 10692 27063 10694 27304
rect 10704 27296 10710 27304
rect 10716 27063 10718 27304
rect 10750 27296 10758 27304
rect 10687 27055 10694 27063
rect 10402 27017 10409 27047
rect 10416 27039 10420 27049
rect 10428 27047 10430 27049
rect 10428 27039 10434 27047
rect 10424 27023 10434 27039
rect 10426 27017 10434 27023
rect 10404 26991 10406 27017
rect 10426 27009 10430 27017
rect 10404 26987 10418 26991
rect 10428 26987 10430 27009
rect 10476 26987 10478 27049
rect 10479 27041 10486 27049
rect 10498 27041 10505 27049
rect 10510 27041 10530 27049
rect 10479 27023 10480 27041
rect 10500 26993 10502 27041
rect 10510 27039 10516 27041
rect 10524 27039 10526 27041
rect 10520 27023 10526 27039
rect 10522 27009 10526 27023
rect 10500 26987 10504 26993
rect 10524 26987 10526 27009
rect 10572 26987 10574 27049
rect 10575 27041 10582 27049
rect 10594 27041 10601 27049
rect 10606 27041 10626 27049
rect 10575 27023 10576 27041
rect 10596 26993 10598 27041
rect 10606 27039 10612 27041
rect 10620 27039 10622 27041
rect 10616 27023 10622 27039
rect 10618 27009 10622 27023
rect 10596 26987 10600 26993
rect 10620 26987 10622 27009
rect 10668 27025 10677 27055
rect 10682 27031 10685 27041
rect 10692 27031 10694 27055
rect 10697 27031 10704 27055
rect 10714 27041 10721 27063
rect 10692 27025 10708 27031
rect 10716 27025 10718 27041
rect 10668 27023 10672 27025
rect 10668 26987 10671 27023
rect 10692 27015 10694 27025
rect 10714 27015 10718 27025
rect 10745 27020 10748 27047
rect 10750 27025 10761 27047
rect 10763 27025 10766 27055
rect 10745 27017 10757 27020
rect 10680 27002 10684 27012
rect 10690 27002 10694 27015
rect 10697 27002 10704 27015
rect 10690 27001 10704 27002
rect 10690 26993 10694 27001
rect 10690 26988 10696 26993
rect 10697 26988 10704 27001
rect 10688 26987 10696 26988
rect 10716 26987 10718 27015
rect 10788 26987 10790 27317
rect 10836 27312 10838 27317
rect 10956 27312 10958 27317
rect 11052 27312 11054 27317
rect 11076 27312 11078 27317
rect 10802 27304 10814 27312
rect 10830 27304 10842 27312
rect 10862 27304 10870 27312
rect 10926 27304 10934 27312
rect 10954 27304 10962 27312
rect 10986 27304 10994 27312
rect 11014 27304 11024 27312
rect 11042 27304 11054 27312
rect 11070 27304 11080 27312
rect 11100 27304 11108 27312
rect 10798 27296 10802 27304
rect 10826 27296 10830 27304
rect 10826 27111 10827 27279
rect 10836 27111 10838 27304
rect 10870 27296 10878 27304
rect 10918 27296 10926 27304
rect 10946 27296 10954 27304
rect 10936 27116 10950 27132
rect 10826 27095 10842 27111
rect 10826 27082 10827 27095
rect 10816 27032 10820 27056
rect 10824 27022 10826 27047
rect 10836 27022 10838 27095
rect 10869 27082 10879 27104
rect 10841 27022 10842 27047
rect 10872 27038 10886 27046
rect 10922 27027 10927 27057
rect 10936 27029 10948 27038
rect 10956 27034 10958 27304
rect 10994 27296 11002 27304
rect 11024 27296 11030 27304
rect 11052 27296 11058 27304
rect 11044 27057 11051 27067
rect 10934 27027 10953 27029
rect 10824 27020 10842 27022
rect 10822 27017 10842 27020
rect 10802 27007 10806 27017
rect 10812 27007 10816 27012
rect 10822 27010 10828 27017
rect 10836 27010 10838 27017
rect 10812 26996 10828 27007
rect 10832 26996 10838 27010
rect 10909 27002 10918 27014
rect 10954 27008 10958 27034
rect 10985 27019 10988 27049
rect 10990 27027 11001 27049
rect 11003 27027 11006 27057
rect 11044 27049 11047 27057
rect 11012 27019 11016 27027
rect 11044 27020 11051 27049
rect 11040 27019 11051 27020
rect 10812 26991 10816 26996
rect 10814 26987 10816 26991
rect 10836 26987 10838 26996
rect 10956 26987 10958 27008
rect 10996 26987 11005 27019
rect 11040 27010 11047 27019
rect 11052 27010 11054 27296
rect 11057 27049 11061 27057
rect 11064 27051 11068 27061
rect 11071 27051 11074 27067
rect 11076 27051 11078 27304
rect 11080 27296 11086 27304
rect 11108 27296 11116 27304
rect 11124 27096 11126 27317
rect 11128 27304 11136 27312
rect 11136 27296 11144 27304
rect 11120 27088 11126 27096
rect 11102 27058 11105 27088
rect 11124 27066 11127 27088
rect 11147 27066 11150 27096
rect 11172 27069 11174 27317
rect 11220 27312 11222 27317
rect 11340 27312 11342 27317
rect 11436 27312 11438 27317
rect 11532 27312 11534 27317
rect 11580 27312 11582 27317
rect 11190 27304 11200 27312
rect 11218 27304 11228 27312
rect 11250 27304 11258 27312
rect 11278 27304 11294 27312
rect 11310 27304 11322 27312
rect 11338 27304 11350 27312
rect 11370 27304 11378 27312
rect 11398 27304 11414 27312
rect 11430 27304 11442 27312
rect 11458 27304 11470 27312
rect 11490 27304 11498 27312
rect 11518 27304 11534 27312
rect 11548 27304 11560 27312
rect 11576 27304 11588 27312
rect 11184 27296 11190 27304
rect 11212 27296 11218 27304
rect 11200 27132 11210 27134
rect 11210 27118 11216 27132
rect 11220 27069 11222 27304
rect 11258 27296 11266 27304
rect 11306 27296 11310 27304
rect 11334 27296 11338 27304
rect 11110 27059 11118 27066
rect 11124 27059 11126 27066
rect 11127 27061 11132 27066
rect 11127 27059 11141 27061
rect 11110 27058 11141 27059
rect 11161 27058 11174 27069
rect 11181 27058 11201 27069
rect 11208 27058 11226 27069
rect 11110 27056 11111 27058
rect 11112 27056 11116 27058
rect 11124 27056 11126 27058
rect 11071 27049 11078 27051
rect 11071 27021 11082 27049
rect 11120 27040 11121 27056
rect 11122 27026 11126 27056
rect 11071 27020 11078 27021
rect 11044 26987 11047 27010
rect 11050 26996 11054 27010
rect 11057 26996 11062 27020
rect 11066 27019 11078 27020
rect 11052 26987 11054 26996
rect 11071 26987 11074 27019
rect 11076 26987 11078 27019
rect 11124 27004 11126 27026
rect 11111 26994 11114 26998
rect 11111 26988 11115 26994
rect 11120 26987 11126 27004
rect 11172 27057 11174 27058
rect 11172 27027 11181 27057
rect 11186 27048 11189 27057
rect 11201 27048 11208 27058
rect 11196 27032 11212 27048
rect 11198 27027 11199 27032
rect 11200 27027 11212 27032
rect 11172 26987 11174 27027
rect 11201 26987 11208 27027
rect 11220 26987 11222 27058
rect 11283 27057 11292 27067
rect 11249 27019 11252 27049
rect 11254 27027 11265 27049
rect 11267 27027 11270 27057
rect 11276 27019 11280 27027
rect 11293 27019 11302 27057
rect 11321 27027 11328 27057
rect 11340 27049 11342 27304
rect 11378 27296 11386 27304
rect 11426 27296 11430 27304
rect 11330 27027 11336 27049
rect 11311 27019 11318 27027
rect 11338 27019 11345 27049
rect 11369 27019 11372 27049
rect 11374 27027 11385 27049
rect 11387 27027 11390 27057
rect 11396 27019 11400 27027
rect 11260 26987 11269 27019
rect 11321 26987 11328 27019
rect 11340 26987 11342 27019
rect 11380 26987 11389 27019
rect 11436 26987 11438 27304
rect 11454 27296 11458 27304
rect 11498 27296 11506 27304
rect 11441 27048 11448 27057
rect 11456 27049 11466 27064
rect 11532 27059 11534 27304
rect 11546 27296 11548 27304
rect 11560 27296 11562 27304
rect 11574 27296 11576 27304
rect 11543 27083 11559 27091
rect 11450 27048 11456 27049
rect 11458 27019 11465 27049
rect 11467 27048 11476 27059
rect 11525 27049 11534 27059
rect 11536 27049 11542 27079
rect 11543 27077 11554 27079
rect 11543 27049 11552 27070
rect 11456 26987 11460 27019
rect 11532 27015 11534 27049
rect 11535 27040 11542 27049
rect 11554 27040 11559 27070
rect 11535 27015 11536 27040
rect 11568 27039 11572 27049
rect 11580 27039 11582 27304
rect 11588 27296 11590 27304
rect 11602 27079 11606 27081
rect 11600 27071 11606 27079
rect 11601 27049 11606 27051
rect 11612 27049 11618 27071
rect 11628 27055 11630 27317
rect 11652 27312 11654 27317
rect 11676 27312 11678 27317
rect 11642 27304 11654 27312
rect 11670 27304 11680 27312
rect 11702 27304 11710 27312
rect 11636 27296 11642 27304
rect 11652 27063 11654 27304
rect 11664 27296 11670 27304
rect 11676 27063 11678 27304
rect 11710 27296 11718 27304
rect 11647 27055 11654 27063
rect 11532 26991 11536 27015
rect 11542 27004 11544 27014
rect 11554 27004 11561 27015
rect 11578 27009 11582 27039
rect 11532 26987 11534 26991
rect 11535 26987 11536 26991
rect 11552 26991 11561 27004
rect 11566 26991 11570 27004
rect 11552 26990 11566 26991
rect 11554 26989 11562 26990
rect 11580 26987 11582 27009
rect 11628 27025 11637 27055
rect 11642 27031 11645 27041
rect 11652 27031 11654 27055
rect 11657 27031 11664 27055
rect 11674 27041 11681 27063
rect 11652 27025 11668 27031
rect 11676 27025 11678 27041
rect 11628 27023 11632 27025
rect 11628 26987 11631 27023
rect 11652 27015 11654 27025
rect 11674 27015 11678 27025
rect 11705 27020 11708 27047
rect 11710 27025 11721 27047
rect 11723 27025 11726 27055
rect 11705 27017 11717 27020
rect 11640 27002 11644 27012
rect 11650 27002 11654 27015
rect 11657 27002 11664 27015
rect 11650 27001 11664 27002
rect 11650 26993 11654 27001
rect 11650 26988 11656 26993
rect 11657 26988 11664 27001
rect 11648 26987 11656 26988
rect 11676 26987 11678 27015
rect 11748 26987 11750 27317
rect 11772 27312 11774 27317
rect 11796 27312 11798 27317
rect 11764 27304 11774 27312
rect 11792 27304 11802 27312
rect 11758 27296 11764 27304
rect 11752 27049 11770 27059
rect 11772 27047 11774 27304
rect 11786 27296 11792 27304
rect 11796 27059 11798 27304
rect 11777 27049 11798 27059
rect 11806 27049 11812 27279
rect 11818 27079 11822 27081
rect 11816 27071 11822 27079
rect 11817 27049 11822 27051
rect 11828 27049 11834 27071
rect 11844 27067 11846 27317
rect 11892 27312 11894 27317
rect 11988 27312 11990 27317
rect 12012 27312 12014 27317
rect 11862 27304 11868 27312
rect 11890 27304 11896 27312
rect 11922 27304 11930 27312
rect 11950 27304 11962 27312
rect 11978 27304 11990 27312
rect 12006 27304 12018 27312
rect 12038 27304 12046 27312
rect 11852 27296 11862 27304
rect 11880 27296 11890 27304
rect 11872 27132 11882 27141
rect 11882 27125 11888 27132
rect 11835 27057 11846 27067
rect 11892 27065 11894 27304
rect 11930 27296 11938 27304
rect 11962 27296 11966 27304
rect 11988 27296 11994 27304
rect 11863 27057 11870 27065
rect 11770 27017 11777 27047
rect 11784 27039 11788 27049
rect 11796 27047 11798 27049
rect 11796 27039 11802 27047
rect 11792 27023 11802 27039
rect 11794 27017 11802 27023
rect 11844 27041 11854 27057
rect 11844 27027 11853 27041
rect 11858 27031 11861 27041
rect 11873 27031 11880 27057
rect 11882 27041 11888 27057
rect 11890 27041 11897 27065
rect 11988 27063 11990 27296
rect 11983 27057 11990 27063
rect 11868 27027 11884 27031
rect 11892 27027 11894 27041
rect 11844 27023 11848 27027
rect 11772 26991 11774 27017
rect 11794 27009 11798 27017
rect 11772 26987 11786 26991
rect 11796 26987 11798 27009
rect 11844 26987 11847 27023
rect 11890 27015 11894 27027
rect 11921 27019 11924 27049
rect 11926 27027 11937 27049
rect 11939 27027 11942 27057
rect 11948 27019 11952 27027
rect 11966 27025 11973 27055
rect 11988 27025 11990 27057
rect 11993 27025 12000 27057
rect 12012 27049 12014 27304
rect 12018 27296 12022 27304
rect 12046 27296 12054 27304
rect 12084 27055 12086 27317
rect 12132 27312 12134 27317
rect 12228 27312 12230 27317
rect 12252 27312 12254 27317
rect 12102 27304 12110 27312
rect 12130 27304 12138 27312
rect 12162 27304 12170 27312
rect 12190 27304 12204 27312
rect 12220 27304 12232 27312
rect 12248 27304 12260 27312
rect 12094 27296 12102 27304
rect 12122 27296 12130 27304
rect 12112 27116 12128 27123
rect 11983 27019 11990 27025
rect 12010 27019 12017 27049
rect 12041 27020 12044 27047
rect 12046 27025 12057 27047
rect 12059 27025 12062 27055
rect 12084 27027 12093 27055
rect 12113 27027 12120 27055
rect 12132 27047 12134 27304
rect 12170 27296 12178 27304
rect 12204 27296 12206 27304
rect 12218 27296 12220 27304
rect 12198 27079 12204 27089
rect 12122 27027 12128 27047
rect 11873 26987 11880 27015
rect 11892 26987 11894 27015
rect 11932 26987 11941 27019
rect 11976 27002 11980 27012
rect 11988 27002 11990 27019
rect 11986 26988 11990 27002
rect 11993 26988 12000 27019
rect 11987 26987 11990 26988
rect 12008 26987 12010 27012
rect 12012 26987 12014 27019
rect 12041 27017 12053 27020
rect 12084 26987 12086 27027
rect 12103 27017 12110 27027
rect 12130 27017 12137 27047
rect 12161 27019 12164 27049
rect 12166 27027 12177 27049
rect 12179 27027 12182 27057
rect 12197 27049 12204 27059
rect 12208 27049 12214 27079
rect 12228 27049 12230 27304
rect 12232 27296 12234 27304
rect 12246 27296 12248 27304
rect 12233 27049 12240 27057
rect 12252 27049 12254 27304
rect 12260 27296 12262 27304
rect 12274 27079 12278 27081
rect 12272 27071 12278 27079
rect 12262 27049 12268 27059
rect 12273 27049 12278 27051
rect 12284 27049 12290 27071
rect 12300 27059 12302 27317
rect 12324 27312 12326 27317
rect 12348 27312 12350 27317
rect 12316 27304 12326 27312
rect 12344 27304 12352 27312
rect 12308 27296 12316 27304
rect 12293 27049 12302 27059
rect 12304 27049 12310 27079
rect 12324 27049 12326 27304
rect 12336 27296 12344 27304
rect 12329 27071 12336 27079
rect 12348 27071 12350 27304
rect 12358 27149 12364 27279
rect 12358 27133 12366 27149
rect 12348 27049 12354 27071
rect 12358 27049 12364 27133
rect 12370 27079 12374 27081
rect 12368 27071 12374 27079
rect 12369 27049 12374 27051
rect 12380 27049 12386 27071
rect 12396 27059 12398 27317
rect 12420 27312 12422 27317
rect 12444 27312 12446 27317
rect 12412 27304 12422 27312
rect 12440 27304 12448 27312
rect 12404 27296 12412 27304
rect 12389 27049 12398 27059
rect 12400 27049 12406 27079
rect 12420 27049 12422 27304
rect 12432 27296 12440 27304
rect 12425 27071 12432 27079
rect 12444 27071 12446 27304
rect 12454 27149 12460 27279
rect 12454 27133 12462 27149
rect 12444 27049 12450 27071
rect 12454 27049 12460 27133
rect 12466 27079 12470 27081
rect 12464 27071 12470 27079
rect 12465 27049 12470 27051
rect 12476 27049 12482 27071
rect 12492 27059 12494 27317
rect 12516 27312 12518 27317
rect 12540 27312 12542 27317
rect 12508 27304 12518 27312
rect 12536 27304 12544 27312
rect 12500 27296 12508 27304
rect 12485 27049 12494 27059
rect 12496 27049 12502 27079
rect 12516 27049 12518 27304
rect 12528 27296 12536 27304
rect 12521 27071 12528 27079
rect 12540 27071 12542 27304
rect 12550 27149 12556 27279
rect 12550 27133 12558 27149
rect 12540 27049 12546 27071
rect 12550 27049 12556 27133
rect 12562 27079 12566 27081
rect 12560 27071 12566 27079
rect 12561 27049 12566 27051
rect 12572 27049 12578 27071
rect 12588 27056 12590 27317
rect 12636 27312 12638 27317
rect 12732 27312 12734 27317
rect 12756 27312 12758 27317
rect 12602 27304 12612 27312
rect 12630 27304 12640 27312
rect 12662 27304 12670 27312
rect 12724 27304 12734 27312
rect 12752 27304 12762 27312
rect 12596 27296 12602 27304
rect 12624 27296 12630 27304
rect 12593 27083 12602 27084
rect 12612 27083 12619 27084
rect 12626 27083 12627 27279
rect 12636 27083 12638 27304
rect 12670 27296 12678 27304
rect 12718 27296 12724 27304
rect 12593 27082 12624 27083
rect 12626 27082 12654 27083
rect 12669 27082 12679 27104
rect 12188 27019 12192 27027
rect 12207 27019 12214 27049
rect 12226 27019 12233 27049
rect 12240 27039 12244 27049
rect 12252 27039 12258 27049
rect 12248 27023 12258 27039
rect 12250 27019 12258 27023
rect 12113 27007 12120 27017
rect 12130 26991 12134 27017
rect 12113 26987 12120 26991
rect 12132 26987 12134 26991
rect 12172 26987 12181 27019
rect 12228 26987 12230 27019
rect 12250 27009 12254 27019
rect 12252 27001 12254 27009
rect 12248 26987 12254 27001
rect 12300 26987 12302 27049
rect 12303 27041 12310 27049
rect 12322 27041 12329 27049
rect 12334 27041 12354 27049
rect 12303 27023 12304 27041
rect 12324 26993 12326 27041
rect 12334 27039 12340 27041
rect 12348 27039 12350 27041
rect 12344 27023 12350 27039
rect 12346 27009 12350 27023
rect 12324 26987 12328 26993
rect 12348 26987 12350 27009
rect 12396 26987 12398 27049
rect 12399 27041 12406 27049
rect 12418 27041 12425 27049
rect 12430 27041 12450 27049
rect 12399 27023 12400 27041
rect 12420 26993 12422 27041
rect 12430 27039 12436 27041
rect 12444 27039 12446 27041
rect 12440 27023 12446 27039
rect 12442 27009 12446 27023
rect 12420 26987 12424 26993
rect 12444 26987 12446 27009
rect 12492 26987 12494 27049
rect 12495 27041 12502 27049
rect 12514 27041 12521 27049
rect 12526 27041 12546 27049
rect 12586 27046 12590 27056
rect 12495 27023 12496 27041
rect 12516 26993 12518 27041
rect 12526 27039 12532 27041
rect 12540 27039 12542 27041
rect 12536 27023 12542 27039
rect 12538 27009 12542 27023
rect 12516 26987 12520 26993
rect 12540 26987 12542 27009
rect 12588 26987 12590 27046
rect 12596 27041 12598 27046
rect 12616 27041 12620 27056
rect 12624 27041 12626 27071
rect 12636 27041 12638 27082
rect 12720 27079 12728 27090
rect 12732 27087 12734 27304
rect 12746 27296 12752 27304
rect 12712 27074 12720 27079
rect 12722 27074 12728 27079
rect 12730 27074 12737 27087
rect 12752 27079 12755 27092
rect 12641 27041 12642 27071
rect 12722 27049 12729 27074
rect 12732 27049 12734 27074
rect 12602 27036 12638 27041
rect 12672 27038 12686 27046
rect 12602 27032 12610 27036
rect 12616 27032 12620 27036
rect 12602 27031 12606 27032
rect 12612 27015 12616 27031
rect 12614 27012 12616 27015
rect 12622 27012 12628 27020
rect 12614 27001 12628 27012
rect 12636 27010 12638 27036
rect 12730 27024 12737 27049
rect 12744 27039 12748 27049
rect 12756 27039 12758 27304
rect 12778 27079 12782 27081
rect 12776 27071 12782 27079
rect 12777 27049 12782 27051
rect 12788 27049 12794 27071
rect 12804 27059 12806 27317
rect 12828 27312 12830 27317
rect 12852 27312 12854 27317
rect 12820 27304 12830 27312
rect 12848 27304 12856 27312
rect 12812 27296 12820 27304
rect 12797 27049 12806 27059
rect 12808 27049 12814 27079
rect 12828 27049 12830 27304
rect 12840 27296 12848 27304
rect 12833 27071 12840 27079
rect 12852 27071 12854 27304
rect 12862 27149 12868 27279
rect 12862 27133 12870 27149
rect 12852 27049 12858 27071
rect 12862 27049 12868 27133
rect 12874 27079 12878 27081
rect 12872 27071 12878 27079
rect 12873 27049 12878 27051
rect 12884 27049 12890 27071
rect 12900 27055 12902 27317
rect 12924 27312 12926 27317
rect 12948 27312 12950 27317
rect 12914 27304 12926 27312
rect 12942 27304 12952 27312
rect 12974 27304 12982 27312
rect 13002 27304 13016 27312
rect 12908 27296 12914 27304
rect 12924 27063 12926 27304
rect 12936 27296 12942 27304
rect 12948 27063 12950 27304
rect 12982 27296 12990 27304
rect 13016 27296 13018 27304
rect 13008 27096 13012 27106
rect 13020 27096 13022 27317
rect 13044 27312 13046 27317
rect 13068 27312 13070 27317
rect 13032 27304 13046 27312
rect 13060 27304 13072 27312
rect 13092 27304 13100 27312
rect 13030 27296 13032 27304
rect 13018 27066 13022 27096
rect 12919 27055 12926 27063
rect 12632 26996 12638 27010
rect 12711 27002 12718 27014
rect 12732 27008 12734 27024
rect 12752 27023 12758 27039
rect 12754 27009 12758 27023
rect 12636 26987 12638 26996
rect 12730 26987 12737 27008
rect 12756 26987 12758 27009
rect 12804 26987 12806 27049
rect 12807 27041 12814 27049
rect 12826 27041 12833 27049
rect 12838 27041 12858 27049
rect 12807 27023 12808 27041
rect 12828 26993 12830 27041
rect 12838 27039 12844 27041
rect 12852 27039 12854 27041
rect 12848 27023 12854 27039
rect 12850 27009 12854 27023
rect 12828 26987 12832 26993
rect 12852 26987 12854 27009
rect 12900 27025 12909 27055
rect 12914 27031 12917 27041
rect 12924 27031 12926 27055
rect 12929 27031 12936 27055
rect 12946 27041 12953 27063
rect 12924 27025 12940 27031
rect 12948 27025 12950 27041
rect 12900 27023 12904 27025
rect 12900 26987 12903 27023
rect 12924 27015 12926 27025
rect 12946 27015 12950 27025
rect 12977 27020 12980 27047
rect 12982 27025 12993 27047
rect 12995 27025 12998 27055
rect 12977 27017 12989 27020
rect 12912 27002 12916 27012
rect 12922 27002 12926 27015
rect 12929 27002 12936 27015
rect 12922 27001 12936 27002
rect 12922 26993 12926 27001
rect 12922 26988 12928 26993
rect 12929 26988 12936 27001
rect 12920 26987 12928 26988
rect 12948 26987 12950 27015
rect 13020 27004 13022 27066
rect 13036 27055 13043 27065
rect 13036 27047 13039 27055
rect 13036 27020 13043 27047
rect 13032 27017 13043 27020
rect 13032 27010 13039 27017
rect 13044 27010 13046 27304
rect 13058 27296 13060 27304
rect 13068 27104 13070 27304
rect 13072 27296 13074 27304
rect 13100 27296 13108 27304
rect 13063 27096 13070 27104
rect 13116 27096 13118 27317
rect 13188 27312 13190 27317
rect 13120 27304 13128 27312
rect 13182 27304 13192 27312
rect 13210 27304 13220 27312
rect 13242 27304 13250 27312
rect 13270 27304 13282 27312
rect 13284 27304 13286 27317
rect 13332 27312 13334 27317
rect 13428 27312 13430 27317
rect 13298 27304 13310 27312
rect 13326 27304 13338 27312
rect 13358 27304 13366 27312
rect 13422 27304 13430 27312
rect 13450 27304 13458 27312
rect 13482 27304 13490 27312
rect 13510 27304 13522 27312
rect 13524 27304 13526 27317
rect 13572 27312 13574 27317
rect 13538 27304 13550 27312
rect 13566 27304 13578 27312
rect 13598 27304 13606 27312
rect 13626 27304 13642 27312
rect 13128 27296 13136 27304
rect 13176 27296 13182 27304
rect 13058 27095 13074 27096
rect 13049 27047 13053 27055
rect 13056 27051 13060 27061
rect 13063 27051 13066 27065
rect 13068 27051 13070 27095
rect 13112 27088 13118 27096
rect 13094 27058 13097 27088
rect 13116 27066 13119 27088
rect 13139 27066 13142 27096
rect 13102 27059 13110 27066
rect 13116 27059 13118 27066
rect 13119 27061 13124 27066
rect 13119 27059 13133 27061
rect 13102 27058 13133 27059
rect 13102 27056 13103 27058
rect 13104 27056 13108 27058
rect 13116 27056 13118 27058
rect 13063 27047 13070 27051
rect 13063 27021 13074 27047
rect 13112 27040 13113 27056
rect 13114 27026 13118 27056
rect 13063 27020 13070 27021
rect 13017 26987 13022 27004
rect 13036 26987 13039 27010
rect 13042 27007 13046 27010
rect 13049 27007 13054 27020
rect 13058 27017 13070 27020
rect 13042 26996 13056 27007
rect 13044 26987 13053 26996
rect 13063 26991 13070 27017
rect 13116 27004 13118 27026
rect 13063 26987 13066 26991
rect 13068 26987 13070 26991
rect 13103 26994 13106 26998
rect 13103 26988 13107 26994
rect 13112 26987 13118 27004
rect 13188 27023 13190 27304
rect 13204 27296 13210 27304
rect 13250 27296 13258 27304
rect 13282 27296 13286 27304
rect 13310 27296 13314 27304
rect 13207 27118 13218 27119
rect 13219 27100 13228 27279
rect 13219 27091 13230 27100
rect 13193 27049 13200 27078
rect 13202 27058 13208 27078
rect 13210 27058 13217 27086
rect 13219 27058 13228 27091
rect 13204 27049 13207 27051
rect 13192 27048 13207 27049
rect 13210 27032 13214 27058
rect 13284 27056 13286 27296
rect 13295 27083 13311 27099
rect 13289 27082 13298 27083
rect 13282 27046 13286 27056
rect 13188 27018 13192 27023
rect 13202 27018 13204 27023
rect 13188 27010 13190 27018
rect 13284 27015 13286 27046
rect 13292 27040 13294 27046
rect 13295 27040 13306 27046
rect 13310 27040 13311 27070
rect 13312 27032 13316 27040
rect 13188 26996 13192 27010
rect 13188 26987 13193 26996
rect 13284 26991 13288 27015
rect 13294 27004 13296 27014
rect 13312 27006 13314 27012
rect 13318 27010 13324 27020
rect 13332 27010 13334 27304
rect 13338 27296 13342 27304
rect 13366 27296 13374 27304
rect 13414 27296 13422 27304
rect 13365 27082 13375 27104
rect 13368 27038 13382 27046
rect 13308 27004 13314 27006
rect 13284 26987 13286 26991
rect 13304 26990 13306 27004
rect 13312 26996 13318 27004
rect 13328 26996 13334 27010
rect 13332 26987 13334 26996
rect 13428 27013 13430 27304
rect 13442 27296 13450 27304
rect 13490 27296 13498 27304
rect 13522 27296 13526 27304
rect 13550 27296 13554 27304
rect 13459 27120 13461 27279
rect 13452 27113 13463 27120
rect 13459 27107 13461 27113
rect 13459 27091 13463 27107
rect 13432 27074 13448 27078
rect 13450 27074 13451 27086
rect 13459 27074 13461 27091
rect 13524 27056 13526 27296
rect 13524 27055 13535 27056
rect 13442 27013 13444 27023
rect 13428 27008 13442 27013
rect 13450 27008 13454 27034
rect 13524 27025 13533 27055
rect 13535 27040 13541 27055
rect 13543 27040 13550 27063
rect 13428 26987 13430 27008
rect 13524 26987 13528 27025
rect 13534 27004 13536 27014
rect 13544 27002 13546 27004
rect 13558 27002 13560 27004
rect 13544 26998 13558 27002
rect 13534 26990 13558 26998
rect 13534 26989 13544 26990
rect 13546 26989 13554 26990
rect 13572 26987 13574 27304
rect 13578 27296 13582 27304
rect 13606 27296 13614 27304
rect 13644 27055 13646 27317
rect 13668 27312 13670 27317
rect 13692 27312 13694 27317
rect 13658 27304 13670 27312
rect 13686 27304 13698 27312
rect 13718 27304 13726 27312
rect 13654 27296 13658 27304
rect 13601 27020 13604 27047
rect 13606 27025 13617 27047
rect 13619 27025 13622 27055
rect 13644 27025 13653 27055
rect 13668 27025 13670 27304
rect 13682 27296 13686 27304
rect 13673 27025 13680 27055
rect 13692 27047 13694 27304
rect 13726 27296 13734 27304
rect 13601 27017 13613 27020
rect 13644 26987 13646 27025
rect 13663 27017 13670 27025
rect 13690 27017 13697 27047
rect 13721 27020 13724 27047
rect 13726 27025 13737 27047
rect 13739 27025 13742 27055
rect 13721 27017 13733 27020
rect 13656 27002 13660 27012
rect 13668 27002 13670 27017
rect 13673 27007 13680 27017
rect 13666 26988 13680 27002
rect 13690 26991 13694 27017
rect 13667 26987 13680 26988
rect 13692 26987 13694 26991
rect 13764 26987 13766 27317
rect 13788 27312 13790 27317
rect 13812 27312 13814 27317
rect 13780 27304 13790 27312
rect 13808 27304 13818 27312
rect 13774 27296 13780 27304
rect 13768 27049 13786 27059
rect 13788 27047 13790 27304
rect 13802 27296 13808 27304
rect 13812 27059 13814 27304
rect 13793 27049 13814 27059
rect 13822 27049 13828 27279
rect 13834 27079 13838 27081
rect 13832 27071 13838 27079
rect 13833 27049 13838 27051
rect 13844 27049 13850 27071
rect 13860 27059 13862 27317
rect 13884 27312 13886 27317
rect 13908 27312 13910 27317
rect 13876 27304 13886 27312
rect 13904 27304 13912 27312
rect 13868 27296 13876 27304
rect 13853 27049 13862 27059
rect 13864 27049 13870 27079
rect 13884 27049 13886 27304
rect 13896 27296 13904 27304
rect 13889 27071 13896 27079
rect 13908 27071 13910 27304
rect 13918 27149 13924 27279
rect 13918 27133 13926 27149
rect 13908 27049 13914 27071
rect 13918 27049 13924 27133
rect 13930 27079 13934 27081
rect 13928 27071 13934 27079
rect 13929 27049 13934 27051
rect 13940 27049 13946 27071
rect 13956 27056 13958 27317
rect 14004 27312 14006 27317
rect 14100 27312 14102 27317
rect 13970 27304 13980 27312
rect 13998 27304 14008 27312
rect 14030 27304 14038 27312
rect 14094 27304 14102 27312
rect 14122 27304 14130 27312
rect 14154 27304 14162 27312
rect 14182 27304 14192 27312
rect 14196 27304 14198 27317
rect 14244 27312 14246 27317
rect 14210 27304 14220 27312
rect 14238 27304 14248 27312
rect 14268 27304 14276 27312
rect 13964 27296 13970 27304
rect 13992 27296 13998 27304
rect 13961 27083 13970 27084
rect 13980 27083 13987 27084
rect 13994 27083 13995 27279
rect 14004 27083 14006 27304
rect 14038 27296 14046 27304
rect 14086 27296 14094 27304
rect 13961 27082 13992 27083
rect 13994 27082 14022 27083
rect 14037 27082 14047 27104
rect 13786 27017 13793 27047
rect 13800 27039 13804 27049
rect 13812 27047 13814 27049
rect 13812 27039 13818 27047
rect 13808 27023 13818 27039
rect 13810 27017 13818 27023
rect 13788 26991 13790 27017
rect 13810 27009 13814 27017
rect 13788 26987 13802 26991
rect 13812 26987 13814 27009
rect 13860 26987 13862 27049
rect 13863 27041 13870 27049
rect 13882 27041 13889 27049
rect 13894 27041 13914 27049
rect 13954 27046 13958 27056
rect 13863 27023 13864 27041
rect 13884 26993 13886 27041
rect 13894 27039 13900 27041
rect 13908 27039 13910 27041
rect 13904 27023 13910 27039
rect 13906 27009 13910 27023
rect 13884 26987 13888 26993
rect 13908 26987 13910 27009
rect 13956 26987 13958 27046
rect 13964 27041 13966 27046
rect 13984 27041 13988 27056
rect 13992 27041 13994 27071
rect 14004 27041 14006 27082
rect 14009 27041 14010 27071
rect 13970 27036 14006 27041
rect 14040 27038 14054 27046
rect 13970 27032 13978 27036
rect 13984 27032 13988 27036
rect 13970 27031 13974 27032
rect 13980 27015 13984 27031
rect 13982 27012 13984 27015
rect 13990 27012 13996 27020
rect 13982 27001 13996 27012
rect 14004 27010 14006 27036
rect 14000 26996 14006 27010
rect 14004 26987 14006 26996
rect 14100 27013 14102 27304
rect 14114 27296 14122 27304
rect 14162 27296 14170 27304
rect 14192 27296 14198 27304
rect 14220 27296 14226 27304
rect 14131 27120 14133 27279
rect 14124 27113 14135 27120
rect 14131 27107 14133 27113
rect 14131 27091 14135 27107
rect 14184 27096 14188 27106
rect 14196 27096 14198 27296
rect 14212 27096 14219 27099
rect 14104 27074 14120 27078
rect 14122 27074 14123 27086
rect 14131 27074 14133 27091
rect 14194 27082 14198 27096
rect 14207 27083 14223 27096
rect 14180 27078 14198 27082
rect 14180 27070 14205 27078
rect 14210 27070 14223 27082
rect 14194 27066 14205 27070
rect 14207 27066 14210 27070
rect 14212 27066 14219 27070
rect 14196 27040 14198 27066
rect 14207 27040 14219 27066
rect 14232 27051 14236 27061
rect 14244 27051 14246 27304
rect 14248 27296 14254 27304
rect 14276 27296 14284 27304
rect 14292 27096 14294 27317
rect 14757 27314 14773 27317
rect 14296 27304 14304 27312
rect 14324 27304 14338 27312
rect 14355 27304 14367 27312
rect 14384 27304 14396 27312
rect 14415 27304 14425 27312
rect 14444 27304 14453 27312
rect 14473 27304 14481 27312
rect 14501 27304 14509 27312
rect 14529 27304 14538 27312
rect 14557 27304 14566 27312
rect 14586 27304 14594 27312
rect 14614 27304 14622 27312
rect 14642 27304 14650 27312
rect 14670 27304 14678 27312
rect 14698 27304 14706 27312
rect 14726 27304 14734 27312
rect 14920 27309 14922 27317
rect 15132 27312 15134 27317
rect 15228 27312 15230 27317
rect 15252 27312 15254 27317
rect 14782 27304 14790 27309
rect 14810 27304 14818 27309
rect 14304 27296 14312 27304
rect 14338 27296 14340 27304
rect 14352 27296 14355 27304
rect 14367 27296 14368 27304
rect 14380 27296 14384 27304
rect 14425 27296 14431 27304
rect 14453 27296 14460 27304
rect 14481 27296 14489 27304
rect 14509 27296 14517 27304
rect 14538 27296 14545 27304
rect 14566 27296 14573 27304
rect 14594 27296 14602 27304
rect 14622 27296 14630 27304
rect 14650 27296 14658 27304
rect 14678 27296 14686 27304
rect 14706 27296 14714 27304
rect 14734 27296 14742 27304
rect 14790 27293 14798 27304
rect 14818 27294 14826 27304
rect 14866 27301 14874 27309
rect 14894 27301 14902 27309
rect 14920 27301 14930 27309
rect 14950 27301 14966 27312
rect 14982 27301 14994 27312
rect 15010 27301 15022 27312
rect 15042 27304 15050 27312
rect 15070 27304 15086 27312
rect 15102 27304 15114 27312
rect 15130 27304 15142 27312
rect 15162 27304 15170 27312
rect 15190 27304 15204 27312
rect 15220 27304 15232 27312
rect 15248 27304 15260 27312
rect 14874 27294 14882 27301
rect 14902 27294 14910 27301
rect 14810 27293 14826 27294
rect 14866 27293 14882 27294
rect 14894 27293 14910 27294
rect 14920 27294 14922 27301
rect 14930 27294 14938 27301
rect 14978 27296 14982 27301
rect 15006 27296 15010 27301
rect 15050 27296 15058 27304
rect 15098 27296 15102 27304
rect 15126 27296 15130 27304
rect 14920 27293 14938 27294
rect 14950 27293 14958 27294
rect 14470 27279 14603 27287
rect 14608 27279 14661 27287
rect 14618 27261 14622 27270
rect 14686 27269 14693 27278
rect 14669 27257 14675 27262
rect 14694 27257 14703 27269
rect 14665 27252 14669 27257
rect 14694 27253 14710 27257
rect 14711 27253 14714 27257
rect 14288 27088 14294 27096
rect 14270 27058 14273 27088
rect 14292 27066 14295 27088
rect 14315 27066 14318 27096
rect 14378 27088 14384 27248
rect 14443 27238 14449 27246
rect 14480 27238 14491 27242
rect 14453 27230 14459 27238
rect 14434 27210 14449 27230
rect 14480 27227 14493 27238
rect 14518 27230 14525 27238
rect 14509 27227 14525 27230
rect 14556 27227 14566 27249
rect 14434 27200 14453 27210
rect 14460 27200 14479 27210
rect 14453 27198 14459 27200
rect 14500 27198 14503 27227
rect 14509 27208 14517 27227
rect 14583 27219 14589 27249
rect 14624 27219 14629 27249
rect 14665 27227 14666 27252
rect 14698 27227 14705 27253
rect 14505 27200 14518 27208
rect 14453 27192 14460 27198
rect 14453 27190 14467 27192
rect 14453 27185 14476 27190
rect 14442 27160 14449 27170
rect 14460 27168 14476 27185
rect 14486 27168 14493 27198
rect 14507 27195 14525 27198
rect 14500 27166 14507 27190
rect 14515 27168 14525 27195
rect 14698 27193 14703 27227
rect 14735 27221 14744 27222
rect 14741 27219 14744 27221
rect 14576 27190 14582 27193
rect 14460 27160 14514 27166
rect 14515 27160 14524 27168
rect 14541 27163 14557 27190
rect 14576 27163 14579 27190
rect 14582 27163 14583 27190
rect 14617 27185 14622 27193
rect 14617 27163 14633 27185
rect 14639 27163 14647 27185
rect 14541 27160 14548 27163
rect 14583 27160 14589 27163
rect 14450 27153 14459 27160
rect 14617 27155 14655 27163
rect 14686 27155 14693 27185
rect 14698 27163 14705 27193
rect 14920 27186 14922 27293
rect 14707 27163 14714 27185
rect 14719 27163 14723 27185
rect 14707 27155 14724 27163
rect 14808 27156 14820 27172
rect 14388 27118 14394 27130
rect 14376 27080 14384 27088
rect 14278 27059 14286 27066
rect 14292 27059 14294 27066
rect 14295 27061 14300 27066
rect 14295 27059 14309 27061
rect 14278 27058 14309 27059
rect 14376 27058 14381 27080
rect 14450 27070 14457 27153
rect 14500 27122 14503 27133
rect 14582 27132 14589 27148
rect 14591 27133 14621 27140
rect 14698 27130 14703 27155
rect 14899 27148 14900 27164
rect 14915 27162 14923 27186
rect 14992 27164 14999 27178
rect 14714 27133 14728 27140
rect 14500 27092 14507 27122
rect 14617 27100 14622 27130
rect 14658 27100 14665 27130
rect 14686 27100 14687 27122
rect 14698 27100 14705 27130
rect 14671 27092 14693 27100
rect 14719 27092 14726 27122
rect 14777 27106 14790 27122
rect 14795 27106 14799 27136
rect 14877 27110 14893 27126
rect 14886 27101 14893 27110
rect 14898 27106 14900 27128
rect 14915 27106 14924 27146
rect 14992 27138 15001 27164
rect 14992 27128 15000 27138
rect 14992 27116 15008 27128
rect 14869 27098 14873 27101
rect 14884 27098 14900 27101
rect 14992 27098 15000 27116
rect 14500 27070 14503 27092
rect 14698 27083 14703 27092
rect 14434 27062 14486 27070
rect 14493 27062 14505 27070
rect 14549 27062 14585 27070
rect 14278 27056 14279 27058
rect 14280 27056 14284 27058
rect 14292 27056 14294 27058
rect 14114 27013 14116 27023
rect 14100 27008 14114 27013
rect 14122 27008 14126 27034
rect 14100 26987 14102 27008
rect 14193 26987 14200 27040
rect 14206 27004 14208 27014
rect 14212 27005 14215 27040
rect 14242 27037 14246 27051
rect 14288 27040 14289 27056
rect 14216 27005 14226 27010
rect 14216 27004 14229 27005
rect 14216 26996 14230 27004
rect 14213 26990 14229 26996
rect 14213 26989 14216 26990
rect 14212 26987 14215 26989
rect 14244 26987 14246 27037
rect 14290 27026 14294 27056
rect 14292 27004 14294 27026
rect 14279 26994 14282 26998
rect 14279 26988 14283 26994
rect 14288 26987 14294 27004
rect 14450 26987 14457 27062
rect 14500 27060 14503 27062
rect 14486 27052 14493 27060
rect 14486 27030 14502 27052
rect 14518 27030 14525 27060
rect 14576 27052 14582 27060
rect 14617 27052 14622 27060
rect 14698 27057 14705 27083
rect 14698 27052 14703 27057
rect 14559 27030 14571 27052
rect 14576 27030 14577 27052
rect 14582 27030 14583 27052
rect 14622 27030 14624 27052
rect 14635 27030 14650 27052
rect 14583 27027 14589 27030
rect 14555 27022 14589 27027
rect 14624 27022 14629 27030
rect 14686 27022 14693 27052
rect 14719 27026 14726 27052
rect 14728 27047 14736 27082
rect 14807 27027 14811 27043
rect 14812 27041 14823 27043
rect 14859 27041 14865 27098
rect 14878 27071 14879 27073
rect 14886 27071 14892 27098
rect 14935 27083 14938 27091
rect 14945 27081 14948 27083
rect 14875 27041 14882 27071
rect 14888 27041 14893 27063
rect 14898 27041 14904 27063
rect 14906 27041 14913 27071
rect 14915 27041 14924 27081
rect 14925 27041 14931 27063
rect 14933 27041 14940 27071
rect 14945 27041 14951 27081
rect 14992 27073 14999 27075
rect 14822 27035 14823 27041
rect 14886 27033 14893 27041
rect 14915 27033 14923 27041
rect 14710 27022 14726 27026
rect 14500 26987 14503 27022
rect 14571 26999 14575 27015
rect 14576 26987 14579 26995
rect 14635 26991 14651 26993
rect 14698 26987 14703 27022
rect 14886 27018 14892 27033
rect 14785 27008 14793 27018
rect 14886 27013 14901 27018
rect 14795 27008 14804 27011
rect 14795 26992 14803 27008
rect 14804 26995 14811 27008
rect 14886 27003 14892 27013
rect 14916 26987 14923 27033
rect 14965 27027 14969 27057
rect 14974 27033 14981 27057
rect 14983 27033 14990 27063
rect 14992 27033 15000 27073
rect 15001 27033 15008 27057
rect 15010 27033 15017 27063
rect 15075 27057 15084 27067
rect 14977 27000 14985 27027
rect 14992 26987 14999 27033
rect 15041 27019 15044 27049
rect 15046 27027 15057 27049
rect 15059 27027 15062 27057
rect 15068 27019 15072 27027
rect 15085 27019 15094 27057
rect 15113 27027 15120 27057
rect 15132 27049 15134 27304
rect 15170 27296 15178 27304
rect 15204 27296 15206 27304
rect 15218 27296 15220 27304
rect 15198 27079 15204 27089
rect 15122 27027 15128 27049
rect 15103 27019 15110 27027
rect 15130 27019 15137 27049
rect 15161 27019 15164 27049
rect 15166 27027 15177 27049
rect 15179 27027 15182 27057
rect 15197 27049 15204 27059
rect 15208 27049 15214 27079
rect 15228 27049 15230 27304
rect 15232 27296 15234 27304
rect 15246 27296 15248 27304
rect 15233 27049 15240 27057
rect 15252 27049 15254 27304
rect 15260 27296 15262 27304
rect 15274 27079 15278 27081
rect 15272 27071 15278 27079
rect 15262 27049 15268 27059
rect 15273 27049 15278 27051
rect 15284 27049 15290 27071
rect 15300 27059 15302 27317
rect 15324 27312 15326 27317
rect 15348 27312 15350 27317
rect 15316 27304 15326 27312
rect 15344 27304 15352 27312
rect 15308 27296 15316 27304
rect 15293 27049 15302 27059
rect 15304 27049 15310 27079
rect 15324 27049 15326 27304
rect 15336 27296 15344 27304
rect 15329 27071 15336 27079
rect 15348 27071 15350 27304
rect 15358 27149 15364 27279
rect 15358 27133 15366 27149
rect 15348 27049 15354 27071
rect 15358 27049 15364 27133
rect 15370 27079 15374 27081
rect 15368 27071 15374 27079
rect 15369 27049 15374 27051
rect 15380 27049 15386 27071
rect 15396 27059 15398 27317
rect 15420 27312 15422 27317
rect 15444 27312 15446 27317
rect 15412 27304 15422 27312
rect 15440 27304 15448 27312
rect 15404 27296 15412 27304
rect 15389 27049 15398 27059
rect 15400 27049 15406 27079
rect 15420 27049 15422 27304
rect 15432 27296 15440 27304
rect 15425 27071 15432 27079
rect 15444 27071 15446 27304
rect 15454 27149 15460 27279
rect 15454 27133 15462 27149
rect 15444 27049 15450 27071
rect 15454 27049 15460 27133
rect 15466 27079 15470 27081
rect 15464 27071 15470 27079
rect 15465 27049 15470 27051
rect 15476 27049 15482 27071
rect 15492 27067 15494 27317
rect 15540 27312 15542 27317
rect 15636 27312 15638 27317
rect 15660 27312 15662 27317
rect 15510 27304 15516 27312
rect 15538 27304 15544 27312
rect 15570 27304 15578 27312
rect 15598 27304 15612 27312
rect 15628 27304 15640 27312
rect 15656 27304 15668 27312
rect 15500 27296 15510 27304
rect 15528 27296 15538 27304
rect 15520 27132 15530 27141
rect 15530 27125 15536 27132
rect 15483 27057 15494 27067
rect 15540 27065 15542 27304
rect 15578 27296 15586 27304
rect 15612 27296 15614 27304
rect 15626 27296 15628 27304
rect 15606 27079 15612 27089
rect 15511 27057 15518 27065
rect 15188 27019 15192 27027
rect 15207 27019 15214 27049
rect 15226 27019 15233 27049
rect 15240 27039 15244 27049
rect 15252 27039 15258 27049
rect 15248 27023 15258 27039
rect 15250 27019 15258 27023
rect 15052 26987 15061 27019
rect 15113 26987 15120 27019
rect 15132 26987 15134 27019
rect 15172 26987 15181 27019
rect 15228 26987 15230 27019
rect 15250 27009 15254 27019
rect 15252 27001 15254 27009
rect 15248 26987 15254 27001
rect 15300 26987 15302 27049
rect 15303 27041 15310 27049
rect 15322 27041 15329 27049
rect 15334 27041 15354 27049
rect 15303 27023 15304 27041
rect 15324 26993 15326 27041
rect 15334 27039 15340 27041
rect 15348 27039 15350 27041
rect 15344 27023 15350 27039
rect 15346 27009 15350 27023
rect 15324 26987 15328 26993
rect 15348 26987 15350 27009
rect 15396 26987 15398 27049
rect 15399 27041 15406 27049
rect 15418 27041 15425 27049
rect 15430 27041 15450 27049
rect 15492 27041 15502 27057
rect 15399 27023 15400 27041
rect 15420 26993 15422 27041
rect 15430 27039 15436 27041
rect 15444 27039 15446 27041
rect 15440 27023 15446 27039
rect 15442 27009 15446 27023
rect 15420 26987 15424 26993
rect 15444 26987 15446 27009
rect 15492 27027 15501 27041
rect 15506 27031 15509 27041
rect 15521 27031 15528 27057
rect 15530 27041 15536 27057
rect 15538 27041 15545 27065
rect 15516 27027 15532 27031
rect 15540 27027 15542 27041
rect 15492 27023 15496 27027
rect 15492 26987 15495 27023
rect 15538 27015 15542 27027
rect 15569 27019 15572 27049
rect 15574 27027 15585 27049
rect 15587 27027 15590 27057
rect 15605 27049 15612 27059
rect 15616 27049 15622 27079
rect 15636 27049 15638 27304
rect 15640 27296 15642 27304
rect 15654 27296 15656 27304
rect 15641 27049 15648 27057
rect 15660 27049 15662 27304
rect 15668 27296 15670 27304
rect 15682 27079 15686 27081
rect 15680 27071 15686 27079
rect 15670 27049 15676 27059
rect 15681 27049 15686 27051
rect 15692 27049 15698 27071
rect 15708 27059 15710 27317
rect 15732 27312 15734 27317
rect 15756 27312 15758 27317
rect 15724 27304 15734 27312
rect 15752 27304 15760 27312
rect 15716 27296 15724 27304
rect 15701 27049 15710 27059
rect 15712 27049 15718 27079
rect 15732 27049 15734 27304
rect 15744 27296 15752 27304
rect 15737 27071 15744 27079
rect 15756 27071 15758 27304
rect 15766 27149 15772 27279
rect 15766 27133 15774 27149
rect 15756 27049 15762 27071
rect 15766 27049 15772 27133
rect 15778 27079 15782 27081
rect 15776 27071 15782 27079
rect 15777 27049 15782 27051
rect 15788 27049 15794 27071
rect 15804 27059 15806 27317
rect 15828 27312 15830 27317
rect 15852 27312 15854 27317
rect 15820 27304 15830 27312
rect 15848 27304 15856 27312
rect 15812 27296 15820 27304
rect 15797 27049 15806 27059
rect 15808 27049 15814 27079
rect 15828 27049 15830 27304
rect 15840 27296 15848 27304
rect 15833 27071 15840 27079
rect 15852 27071 15854 27304
rect 15862 27149 15868 27279
rect 15862 27133 15870 27149
rect 15852 27049 15858 27071
rect 15862 27049 15868 27133
rect 15874 27079 15878 27081
rect 15872 27071 15878 27079
rect 15873 27049 15878 27051
rect 15884 27049 15890 27071
rect 15900 27059 15902 27317
rect 15924 27312 15926 27317
rect 15948 27312 15950 27317
rect 15916 27304 15926 27312
rect 15944 27304 15952 27312
rect 15908 27296 15916 27304
rect 15893 27049 15902 27059
rect 15904 27049 15910 27079
rect 15924 27049 15926 27304
rect 15936 27296 15944 27304
rect 15929 27071 15936 27079
rect 15948 27071 15950 27304
rect 15958 27149 15964 27279
rect 15958 27133 15966 27149
rect 15948 27049 15954 27071
rect 15958 27049 15964 27133
rect 15970 27079 15974 27081
rect 15968 27071 15974 27079
rect 15969 27049 15974 27051
rect 15980 27049 15986 27071
rect 15996 27059 15998 27317
rect 16020 27312 16022 27317
rect 16044 27312 16046 27317
rect 16012 27304 16022 27312
rect 16040 27304 16048 27312
rect 16004 27296 16012 27304
rect 15989 27049 15998 27059
rect 16000 27049 16006 27079
rect 16020 27049 16022 27304
rect 16032 27296 16040 27304
rect 16025 27071 16032 27079
rect 16044 27071 16046 27304
rect 16054 27149 16060 27279
rect 16054 27133 16062 27149
rect 16044 27049 16050 27071
rect 16054 27049 16060 27133
rect 16066 27079 16070 27081
rect 16064 27071 16070 27079
rect 16065 27049 16070 27051
rect 16076 27049 16082 27071
rect 16092 27067 16094 27317
rect 16140 27312 16142 27317
rect 16236 27312 16238 27317
rect 16260 27312 16262 27317
rect 16110 27304 16116 27312
rect 16138 27304 16144 27312
rect 16170 27304 16178 27312
rect 16198 27304 16212 27312
rect 16228 27304 16240 27312
rect 16256 27304 16268 27312
rect 16100 27296 16110 27304
rect 16128 27296 16138 27304
rect 16120 27132 16130 27141
rect 16130 27125 16136 27132
rect 16083 27057 16094 27067
rect 16140 27065 16142 27304
rect 16178 27296 16186 27304
rect 16212 27296 16214 27304
rect 16226 27296 16228 27304
rect 16206 27079 16212 27089
rect 16111 27057 16118 27065
rect 15596 27019 15600 27027
rect 15615 27019 15622 27049
rect 15634 27019 15641 27049
rect 15648 27039 15652 27049
rect 15660 27039 15666 27049
rect 15656 27023 15666 27039
rect 15658 27019 15666 27023
rect 15521 26987 15528 27015
rect 15540 26987 15542 27015
rect 15580 26987 15589 27019
rect 15636 26987 15638 27019
rect 15658 27009 15662 27019
rect 15660 27001 15662 27009
rect 15656 26987 15662 27001
rect 15708 26987 15710 27049
rect 15711 27041 15718 27049
rect 15730 27041 15737 27049
rect 15742 27041 15762 27049
rect 15711 27023 15712 27041
rect 15732 26993 15734 27041
rect 15742 27039 15748 27041
rect 15756 27039 15758 27041
rect 15752 27023 15758 27039
rect 15754 27009 15758 27023
rect 15732 26987 15736 26993
rect 15756 26987 15758 27009
rect 15804 26987 15806 27049
rect 15807 27041 15814 27049
rect 15826 27041 15833 27049
rect 15838 27041 15858 27049
rect 15807 27023 15808 27041
rect 15828 26993 15830 27041
rect 15838 27039 15844 27041
rect 15852 27039 15854 27041
rect 15848 27023 15854 27039
rect 15850 27009 15854 27023
rect 15828 26987 15832 26993
rect 15852 26987 15854 27009
rect 15900 26987 15902 27049
rect 15903 27041 15910 27049
rect 15922 27041 15929 27049
rect 15934 27041 15954 27049
rect 15903 27023 15904 27041
rect 15924 26993 15926 27041
rect 15934 27039 15940 27041
rect 15948 27039 15950 27041
rect 15944 27023 15950 27039
rect 15946 27009 15950 27023
rect 15924 26987 15928 26993
rect 15948 26987 15950 27009
rect 15996 26987 15998 27049
rect 15999 27041 16006 27049
rect 16018 27041 16025 27049
rect 16030 27041 16050 27049
rect 16092 27041 16102 27057
rect 15999 27023 16000 27041
rect 16020 26993 16022 27041
rect 16030 27039 16036 27041
rect 16044 27039 16046 27041
rect 16040 27023 16046 27039
rect 16042 27009 16046 27023
rect 16020 26987 16024 26993
rect 16044 26987 16046 27009
rect 16092 27027 16101 27041
rect 16106 27031 16109 27041
rect 16121 27031 16128 27057
rect 16130 27041 16136 27057
rect 16138 27041 16145 27065
rect 16116 27027 16132 27031
rect 16140 27027 16142 27041
rect 16092 27023 16096 27027
rect 16092 26987 16095 27023
rect 16138 27015 16142 27027
rect 16169 27019 16172 27049
rect 16174 27027 16185 27049
rect 16187 27027 16190 27057
rect 16205 27049 16212 27059
rect 16216 27049 16222 27079
rect 16236 27049 16238 27304
rect 16240 27296 16242 27304
rect 16254 27296 16256 27304
rect 16241 27049 16248 27057
rect 16260 27049 16262 27304
rect 16268 27296 16270 27304
rect 16282 27079 16286 27081
rect 16280 27071 16286 27079
rect 16270 27049 16276 27059
rect 16281 27049 16286 27051
rect 16292 27049 16298 27071
rect 16308 27059 16310 27317
rect 16332 27312 16334 27317
rect 16356 27312 16358 27317
rect 16324 27304 16334 27312
rect 16352 27304 16360 27312
rect 16316 27296 16324 27304
rect 16301 27049 16310 27059
rect 16312 27049 16318 27079
rect 16332 27049 16334 27304
rect 16344 27296 16352 27304
rect 16337 27071 16344 27079
rect 16356 27071 16358 27304
rect 16366 27149 16372 27279
rect 16366 27133 16374 27149
rect 16356 27049 16362 27071
rect 16366 27049 16372 27133
rect 16378 27079 16382 27081
rect 16376 27071 16382 27079
rect 16377 27049 16382 27051
rect 16388 27049 16394 27071
rect 16404 27056 16406 27317
rect 16452 27312 16454 27317
rect 16548 27312 16550 27317
rect 16572 27312 16574 27317
rect 16418 27304 16428 27312
rect 16446 27304 16456 27312
rect 16478 27304 16486 27312
rect 16540 27304 16550 27312
rect 16568 27304 16578 27312
rect 16412 27296 16418 27304
rect 16440 27296 16446 27304
rect 16409 27083 16418 27084
rect 16428 27083 16435 27084
rect 16442 27083 16443 27279
rect 16452 27083 16454 27304
rect 16486 27296 16494 27304
rect 16534 27296 16540 27304
rect 16409 27082 16440 27083
rect 16442 27082 16470 27083
rect 16485 27082 16495 27104
rect 16196 27019 16200 27027
rect 16215 27019 16222 27049
rect 16234 27019 16241 27049
rect 16248 27039 16252 27049
rect 16260 27039 16266 27049
rect 16256 27023 16266 27039
rect 16258 27019 16266 27023
rect 16121 26987 16128 27015
rect 16140 26987 16142 27015
rect 16180 26987 16189 27019
rect 16236 26987 16238 27019
rect 16258 27009 16262 27019
rect 16260 27001 16262 27009
rect 16256 26987 16262 27001
rect 16308 26987 16310 27049
rect 16311 27041 16318 27049
rect 16330 27041 16337 27049
rect 16342 27041 16362 27049
rect 16402 27046 16406 27056
rect 16311 27023 16312 27041
rect 16332 26993 16334 27041
rect 16342 27039 16348 27041
rect 16356 27039 16358 27041
rect 16352 27023 16358 27039
rect 16354 27009 16358 27023
rect 16332 26987 16336 26993
rect 16356 26987 16358 27009
rect 16404 26987 16406 27046
rect 16412 27041 16414 27046
rect 16432 27041 16436 27056
rect 16440 27041 16442 27071
rect 16452 27041 16454 27082
rect 16536 27079 16544 27090
rect 16548 27087 16550 27304
rect 16562 27296 16568 27304
rect 16528 27074 16536 27079
rect 16538 27074 16544 27079
rect 16546 27074 16553 27087
rect 16568 27079 16571 27092
rect 16457 27041 16458 27071
rect 16538 27049 16545 27074
rect 16548 27049 16550 27074
rect 16418 27036 16454 27041
rect 16488 27038 16502 27046
rect 16418 27032 16426 27036
rect 16432 27032 16436 27036
rect 16418 27031 16422 27032
rect 16428 27015 16432 27031
rect 16430 27012 16432 27015
rect 16438 27012 16444 27020
rect 16430 27001 16444 27012
rect 16452 27010 16454 27036
rect 16546 27024 16553 27049
rect 16560 27039 16564 27049
rect 16572 27039 16574 27304
rect 16594 27079 16598 27081
rect 16592 27071 16598 27079
rect 16593 27049 16598 27051
rect 16604 27049 16610 27071
rect 16620 27059 16622 27317
rect 16644 27312 16646 27317
rect 16668 27312 16670 27317
rect 16636 27304 16646 27312
rect 16664 27304 16672 27312
rect 16628 27296 16636 27304
rect 16613 27049 16622 27059
rect 16624 27049 16630 27079
rect 16644 27049 16646 27304
rect 16656 27296 16664 27304
rect 16649 27071 16656 27079
rect 16668 27071 16670 27304
rect 16678 27149 16684 27279
rect 16678 27133 16686 27149
rect 16668 27049 16674 27071
rect 16678 27049 16684 27133
rect 16690 27079 16694 27081
rect 16688 27071 16694 27079
rect 16689 27049 16694 27051
rect 16700 27049 16706 27071
rect 16716 27055 16718 27317
rect 16740 27312 16742 27317
rect 16764 27312 16766 27317
rect 16730 27304 16742 27312
rect 16758 27304 16768 27312
rect 16790 27304 16798 27312
rect 16818 27304 16834 27312
rect 16724 27296 16730 27304
rect 16740 27063 16742 27304
rect 16752 27296 16758 27304
rect 16764 27063 16766 27304
rect 16798 27296 16806 27304
rect 16735 27055 16742 27063
rect 16448 26996 16454 27010
rect 16527 27002 16534 27014
rect 16548 27008 16550 27024
rect 16568 27023 16574 27039
rect 16570 27009 16574 27023
rect 16452 26987 16454 26996
rect 16546 26987 16553 27008
rect 16572 26987 16574 27009
rect 16620 26987 16622 27049
rect 16623 27041 16630 27049
rect 16642 27041 16649 27049
rect 16654 27041 16674 27049
rect 16623 27023 16624 27041
rect 16644 26993 16646 27041
rect 16654 27039 16660 27041
rect 16668 27039 16670 27041
rect 16664 27023 16670 27039
rect 16666 27009 16670 27023
rect 16644 26987 16648 26993
rect 16668 26987 16670 27009
rect 16716 27025 16725 27055
rect 16730 27031 16733 27041
rect 16740 27031 16742 27055
rect 16745 27031 16752 27055
rect 16762 27041 16769 27063
rect 16740 27025 16756 27031
rect 16764 27025 16766 27041
rect 16716 27023 16720 27025
rect 16716 26987 16719 27023
rect 16740 27015 16742 27025
rect 16762 27015 16766 27025
rect 16793 27020 16796 27047
rect 16798 27025 16809 27047
rect 16811 27025 16814 27055
rect 16793 27017 16805 27020
rect 16728 27002 16732 27012
rect 16738 27002 16742 27015
rect 16745 27002 16752 27015
rect 16738 27001 16752 27002
rect 16738 26993 16742 27001
rect 16738 26988 16744 26993
rect 16745 26988 16752 27001
rect 16736 26987 16744 26988
rect 16764 26987 16766 27015
rect 16836 26987 16838 27317
rect 16884 27312 16886 27317
rect 16980 27312 16982 27317
rect 17004 27312 17006 27317
rect 16850 27304 16862 27312
rect 16878 27304 16890 27312
rect 16910 27304 16918 27312
rect 16972 27304 16982 27312
rect 17000 27304 17010 27312
rect 16846 27296 16850 27304
rect 16874 27296 16878 27304
rect 16874 27111 16875 27279
rect 16884 27111 16886 27304
rect 16918 27296 16926 27304
rect 16966 27296 16972 27304
rect 16874 27095 16890 27111
rect 16874 27082 16875 27095
rect 16864 27032 16868 27056
rect 16872 27022 16874 27047
rect 16884 27022 16886 27095
rect 16917 27082 16927 27104
rect 16968 27079 16976 27090
rect 16980 27087 16982 27304
rect 16994 27296 17000 27304
rect 16960 27074 16968 27079
rect 16970 27074 16976 27079
rect 16978 27074 16985 27087
rect 17000 27079 17003 27092
rect 16970 27049 16977 27074
rect 16980 27049 16982 27074
rect 16889 27022 16890 27047
rect 16920 27038 16934 27046
rect 16978 27024 16985 27049
rect 16992 27039 16996 27049
rect 17004 27039 17006 27304
rect 17026 27079 17030 27081
rect 17024 27071 17030 27079
rect 17025 27049 17030 27051
rect 17036 27049 17042 27071
rect 17052 27067 17054 27317
rect 17100 27312 17102 27317
rect 17196 27312 17198 27317
rect 17220 27312 17222 27317
rect 17070 27304 17076 27312
rect 17098 27304 17104 27312
rect 17130 27304 17138 27312
rect 17158 27304 17172 27312
rect 17188 27304 17200 27312
rect 17216 27304 17228 27312
rect 17060 27296 17070 27304
rect 17088 27296 17098 27304
rect 17080 27132 17090 27141
rect 17090 27125 17096 27132
rect 17043 27057 17054 27067
rect 17100 27065 17102 27304
rect 17138 27296 17146 27304
rect 17172 27296 17174 27304
rect 17186 27296 17188 27304
rect 17166 27079 17172 27089
rect 17071 27057 17078 27065
rect 16872 27020 16890 27022
rect 16870 27017 16890 27020
rect 16850 27007 16854 27017
rect 16860 27007 16864 27012
rect 16870 27010 16876 27017
rect 16884 27010 16886 27017
rect 16860 26996 16876 27007
rect 16880 26996 16886 27010
rect 16959 27002 16966 27014
rect 16980 27008 16982 27024
rect 17000 27023 17006 27039
rect 17002 27009 17006 27023
rect 16860 26991 16864 26996
rect 16862 26987 16864 26991
rect 16884 26987 16886 26996
rect 16978 26987 16985 27008
rect 17004 26987 17006 27009
rect 17052 27041 17062 27057
rect 17052 27027 17061 27041
rect 17066 27031 17069 27041
rect 17081 27031 17088 27057
rect 17090 27041 17096 27057
rect 17098 27041 17105 27065
rect 17076 27027 17092 27031
rect 17100 27027 17102 27041
rect 17052 27023 17056 27027
rect 17052 26987 17055 27023
rect 17098 27015 17102 27027
rect 17129 27019 17132 27049
rect 17134 27027 17145 27049
rect 17147 27027 17150 27057
rect 17165 27049 17172 27059
rect 17176 27049 17182 27079
rect 17196 27049 17198 27304
rect 17200 27296 17202 27304
rect 17214 27296 17216 27304
rect 17201 27049 17208 27057
rect 17220 27049 17222 27304
rect 17228 27296 17230 27304
rect 17242 27079 17246 27081
rect 17240 27071 17246 27079
rect 17230 27049 17236 27059
rect 17241 27049 17246 27051
rect 17252 27049 17258 27071
rect 17268 27059 17270 27317
rect 17292 27312 17294 27317
rect 17316 27312 17318 27317
rect 17781 27314 17797 27317
rect 17284 27304 17294 27312
rect 17312 27304 17320 27312
rect 17379 27304 17388 27312
rect 17408 27304 17416 27312
rect 17439 27304 17449 27312
rect 17468 27304 17477 27312
rect 17497 27304 17505 27312
rect 17525 27304 17533 27312
rect 17553 27304 17562 27312
rect 17581 27304 17590 27312
rect 17610 27304 17618 27312
rect 17638 27304 17646 27312
rect 17666 27304 17674 27312
rect 17694 27304 17702 27312
rect 17722 27304 17730 27312
rect 17750 27304 17758 27312
rect 17944 27309 17946 27317
rect 17806 27304 17814 27309
rect 17834 27304 17842 27309
rect 17276 27296 17284 27304
rect 17261 27049 17270 27059
rect 17272 27049 17278 27079
rect 17292 27049 17294 27304
rect 17304 27296 17312 27304
rect 17297 27071 17304 27079
rect 17316 27071 17318 27304
rect 17372 27296 17379 27304
rect 17400 27296 17408 27304
rect 17449 27296 17455 27304
rect 17477 27296 17484 27304
rect 17505 27296 17513 27304
rect 17533 27296 17541 27304
rect 17562 27296 17569 27304
rect 17590 27296 17597 27304
rect 17618 27296 17626 27304
rect 17646 27296 17654 27304
rect 17674 27296 17682 27304
rect 17702 27296 17710 27304
rect 17730 27296 17738 27304
rect 17758 27296 17766 27304
rect 17814 27293 17822 27304
rect 17842 27294 17850 27304
rect 17890 27301 17898 27309
rect 17918 27301 17926 27309
rect 17944 27301 17954 27309
rect 17974 27301 17988 27312
rect 18004 27301 18016 27312
rect 18032 27301 18044 27312
rect 18064 27304 18080 27312
rect 17898 27294 17906 27301
rect 17926 27294 17934 27301
rect 17834 27293 17850 27294
rect 17890 27293 17906 27294
rect 17918 27293 17934 27294
rect 17944 27294 17946 27301
rect 17954 27294 17962 27301
rect 17988 27296 17990 27301
rect 18002 27296 18004 27301
rect 18016 27296 18018 27301
rect 18030 27296 18032 27301
rect 18044 27296 18046 27301
rect 17944 27293 17962 27294
rect 17974 27293 17982 27294
rect 17494 27279 17627 27287
rect 17632 27279 17685 27287
rect 17326 27149 17332 27279
rect 17642 27261 17646 27270
rect 17710 27269 17717 27278
rect 17693 27257 17699 27262
rect 17718 27257 17727 27269
rect 17689 27252 17693 27257
rect 17718 27253 17734 27257
rect 17735 27253 17738 27257
rect 17326 27133 17334 27149
rect 17316 27049 17322 27071
rect 17326 27049 17332 27133
rect 17338 27079 17342 27081
rect 17402 27080 17408 27248
rect 17467 27238 17473 27246
rect 17504 27238 17515 27242
rect 17477 27230 17483 27238
rect 17458 27210 17473 27230
rect 17504 27227 17517 27238
rect 17542 27230 17549 27238
rect 17533 27227 17549 27230
rect 17580 27227 17590 27249
rect 17458 27200 17477 27210
rect 17484 27200 17503 27210
rect 17477 27198 17483 27200
rect 17524 27198 17527 27227
rect 17533 27208 17541 27227
rect 17607 27219 17613 27249
rect 17648 27219 17653 27249
rect 17689 27227 17690 27252
rect 17722 27227 17729 27253
rect 17529 27200 17542 27208
rect 17477 27192 17484 27198
rect 17477 27190 17491 27192
rect 17477 27185 17500 27190
rect 17466 27160 17473 27170
rect 17484 27168 17500 27185
rect 17510 27168 17517 27198
rect 17531 27195 17549 27198
rect 17524 27166 17531 27190
rect 17539 27168 17549 27195
rect 17722 27193 17727 27227
rect 17759 27221 17768 27222
rect 17765 27219 17768 27221
rect 17600 27190 17606 27193
rect 17484 27160 17538 27166
rect 17539 27160 17548 27168
rect 17565 27163 17581 27190
rect 17600 27163 17603 27190
rect 17606 27163 17607 27190
rect 17641 27185 17646 27193
rect 17641 27163 17657 27185
rect 17663 27163 17671 27185
rect 17565 27160 17572 27163
rect 17607 27160 17613 27163
rect 17474 27153 17483 27160
rect 17641 27155 17679 27163
rect 17710 27155 17717 27185
rect 17722 27163 17729 27193
rect 17944 27186 17946 27293
rect 17731 27163 17738 27185
rect 17743 27163 17747 27185
rect 17731 27155 17748 27163
rect 17832 27156 17844 27172
rect 17412 27125 17418 27130
rect 17336 27071 17342 27079
rect 17337 27049 17342 27051
rect 17348 27049 17354 27071
rect 17156 27019 17160 27027
rect 17175 27019 17182 27049
rect 17194 27019 17201 27049
rect 17208 27039 17212 27049
rect 17220 27039 17226 27049
rect 17216 27023 17226 27039
rect 17218 27019 17226 27023
rect 17081 26987 17088 27015
rect 17100 26987 17102 27015
rect 17140 26987 17149 27019
rect 17196 26987 17198 27019
rect 17218 27009 17222 27019
rect 17220 27001 17222 27009
rect 17216 26987 17222 27001
rect 17268 26987 17270 27049
rect 17271 27041 17278 27049
rect 17290 27041 17297 27049
rect 17302 27041 17322 27049
rect 17400 27041 17405 27071
rect 17474 27070 17481 27153
rect 17524 27122 17527 27133
rect 17606 27132 17613 27148
rect 17615 27133 17645 27140
rect 17722 27130 17727 27155
rect 17923 27148 17924 27164
rect 17939 27162 17947 27186
rect 17738 27133 17752 27140
rect 17524 27092 17531 27122
rect 17641 27100 17646 27130
rect 17682 27100 17689 27130
rect 17710 27100 17711 27122
rect 17722 27100 17729 27130
rect 17695 27092 17717 27100
rect 17743 27092 17750 27122
rect 17801 27106 17814 27122
rect 17819 27106 17823 27136
rect 17901 27110 17917 27126
rect 17910 27101 17917 27110
rect 17922 27106 17924 27128
rect 17939 27106 17948 27146
rect 18046 27140 18051 27279
rect 18046 27133 18053 27140
rect 17893 27098 17897 27101
rect 17908 27098 17924 27101
rect 18046 27098 18051 27133
rect 17524 27070 17527 27092
rect 17722 27083 17727 27092
rect 17458 27062 17510 27070
rect 17517 27062 17529 27070
rect 17573 27062 17609 27070
rect 17271 27023 17272 27041
rect 17292 26993 17294 27041
rect 17302 27039 17308 27041
rect 17316 27039 17318 27041
rect 17312 27023 17318 27039
rect 17314 27009 17318 27023
rect 17292 26987 17296 26993
rect 17316 26987 17318 27009
rect 17474 26987 17481 27062
rect 17524 27060 17527 27062
rect 17510 27052 17517 27060
rect 17510 27030 17526 27052
rect 17542 27030 17549 27060
rect 17600 27052 17606 27060
rect 17641 27052 17646 27060
rect 17722 27057 17729 27083
rect 17722 27052 17727 27057
rect 17583 27030 17595 27052
rect 17600 27030 17601 27052
rect 17606 27030 17607 27052
rect 17646 27030 17648 27052
rect 17659 27030 17674 27052
rect 17607 27027 17613 27030
rect 17579 27022 17613 27027
rect 17648 27022 17653 27030
rect 17710 27022 17717 27052
rect 17743 27026 17750 27052
rect 17752 27047 17760 27082
rect 17831 27027 17835 27043
rect 17836 27041 17847 27043
rect 17883 27041 17889 27098
rect 17902 27071 17903 27073
rect 17910 27071 17916 27098
rect 18072 27096 18076 27106
rect 18084 27096 18086 27317
rect 18108 27312 18110 27317
rect 18132 27312 18134 27317
rect 18096 27304 18110 27312
rect 18124 27304 18136 27312
rect 18156 27304 18164 27312
rect 18092 27296 18096 27304
rect 17959 27083 17962 27091
rect 17969 27081 17972 27083
rect 17899 27041 17906 27071
rect 17912 27041 17917 27063
rect 17922 27041 17928 27063
rect 17930 27041 17937 27071
rect 17939 27041 17948 27081
rect 17949 27041 17955 27063
rect 17957 27041 17964 27071
rect 17969 27041 17975 27081
rect 17992 27049 17993 27079
rect 18008 27063 18014 27065
rect 18017 27063 18023 27079
rect 18046 27073 18048 27093
rect 18082 27082 18086 27096
rect 18058 27079 18062 27081
rect 17998 27049 18008 27063
rect 18010 27049 18014 27063
rect 18016 27049 18017 27063
rect 17846 27035 17847 27041
rect 17910 27033 17917 27041
rect 17939 27033 17947 27041
rect 18010 27033 18016 27049
rect 18037 27043 18041 27063
rect 18046 27049 18051 27073
rect 18056 27071 18062 27079
rect 18068 27079 18086 27082
rect 18068 27071 18093 27079
rect 18057 27049 18062 27051
rect 18068 27049 18074 27071
rect 18082 27066 18093 27071
rect 18037 27039 18042 27043
rect 18084 27041 18086 27066
rect 18032 27033 18041 27039
rect 17734 27022 17750 27026
rect 17524 26987 17527 27022
rect 17595 26999 17599 27015
rect 17600 26987 17603 26995
rect 17659 26991 17675 26993
rect 17722 26987 17727 27022
rect 17910 27018 17916 27033
rect 17809 27008 17817 27018
rect 17910 27013 17925 27018
rect 17819 27008 17828 27011
rect 17819 26992 17827 27008
rect 17828 26995 17835 27008
rect 17910 27003 17916 27013
rect 17940 26987 17947 27033
rect 18032 27023 18033 27033
rect 18081 27023 18088 27041
rect 18100 27031 18107 27066
rect 18108 27031 18110 27304
rect 18120 27296 18124 27304
rect 18113 27071 18120 27079
rect 18132 27071 18134 27304
rect 18164 27296 18172 27304
rect 18180 27096 18182 27317
rect 18252 27312 18254 27317
rect 18348 27312 18350 27317
rect 18396 27312 18398 27317
rect 18492 27312 18494 27317
rect 18516 27312 18518 27317
rect 18184 27304 18192 27312
rect 18246 27304 18256 27312
rect 18274 27304 18284 27312
rect 18306 27304 18314 27312
rect 18334 27304 18350 27312
rect 18366 27304 18378 27312
rect 18394 27304 18406 27312
rect 18426 27304 18434 27312
rect 18454 27304 18468 27312
rect 18484 27304 18496 27312
rect 18512 27304 18524 27312
rect 18192 27296 18200 27304
rect 18240 27296 18246 27304
rect 18176 27088 18182 27096
rect 18113 27066 18117 27071
rect 18127 27051 18134 27071
rect 18158 27058 18161 27088
rect 18180 27066 18183 27088
rect 18203 27066 18206 27096
rect 18166 27059 18174 27066
rect 18180 27059 18182 27066
rect 18183 27061 18188 27066
rect 18183 27059 18197 27061
rect 18166 27058 18197 27059
rect 18166 27056 18167 27058
rect 18168 27056 18172 27058
rect 18180 27056 18182 27058
rect 18127 27047 18138 27051
rect 18122 27041 18138 27047
rect 18113 27031 18117 27041
rect 18002 26991 18011 27001
rect 18012 26990 18021 26991
rect 18081 26987 18087 27023
rect 18100 27020 18103 27031
rect 18096 27010 18103 27020
rect 18108 27020 18117 27031
rect 18108 27015 18118 27020
rect 18100 26990 18103 27010
rect 18106 27010 18110 27015
rect 18113 27010 18118 27015
rect 18127 27015 18134 27041
rect 18176 27040 18177 27056
rect 18178 27026 18182 27056
rect 18106 27001 18120 27010
rect 18106 26996 18110 27001
rect 18113 26996 18118 27001
rect 18092 26987 18103 26990
rect 18108 26993 18110 26996
rect 18108 26987 18112 26993
rect 18127 26987 18130 27015
rect 18132 26987 18134 27015
rect 18180 27004 18182 27026
rect 18167 26994 18170 26998
rect 18167 26988 18171 26994
rect 18176 26987 18182 27004
rect 18252 27023 18254 27304
rect 18268 27296 18274 27304
rect 18314 27296 18322 27304
rect 18271 27118 18282 27119
rect 18283 27100 18292 27279
rect 18283 27091 18294 27100
rect 18257 27049 18264 27078
rect 18266 27058 18272 27078
rect 18274 27058 18281 27086
rect 18283 27058 18292 27091
rect 18348 27067 18350 27304
rect 18362 27296 18366 27304
rect 18390 27296 18394 27304
rect 18268 27049 18271 27051
rect 18256 27048 18271 27049
rect 18274 27032 18278 27058
rect 18339 27057 18350 27067
rect 18348 27040 18358 27057
rect 18359 27040 18365 27057
rect 18367 27040 18374 27065
rect 18376 27040 18385 27279
rect 18348 27027 18357 27040
rect 18252 27018 18256 27023
rect 18266 27018 18268 27023
rect 18252 27010 18254 27018
rect 18252 26996 18256 27010
rect 18252 26987 18257 26996
rect 18348 26987 18352 27027
rect 18358 27004 18360 27014
rect 18368 26990 18370 27004
rect 18396 26987 18398 27304
rect 18434 27296 18442 27304
rect 18468 27296 18470 27304
rect 18482 27296 18484 27304
rect 18462 27079 18468 27089
rect 18425 27019 18428 27049
rect 18430 27027 18441 27049
rect 18443 27027 18446 27057
rect 18461 27049 18468 27059
rect 18472 27049 18478 27079
rect 18492 27049 18494 27304
rect 18496 27296 18498 27304
rect 18510 27296 18512 27304
rect 18497 27049 18504 27057
rect 18516 27049 18518 27304
rect 18524 27296 18526 27304
rect 18538 27079 18542 27081
rect 18536 27071 18542 27079
rect 18526 27049 18532 27059
rect 18537 27049 18542 27051
rect 18548 27049 18554 27071
rect 18564 27059 18566 27317
rect 18588 27312 18590 27317
rect 18612 27312 18614 27317
rect 18580 27304 18590 27312
rect 18608 27304 18616 27312
rect 18572 27296 18580 27304
rect 18557 27049 18566 27059
rect 18568 27049 18574 27079
rect 18588 27049 18590 27304
rect 18600 27296 18608 27304
rect 18593 27071 18600 27079
rect 18612 27071 18614 27304
rect 18622 27149 18628 27279
rect 18622 27133 18630 27149
rect 18612 27049 18618 27071
rect 18622 27049 18628 27133
rect 18634 27079 18638 27081
rect 18632 27071 18638 27079
rect 18633 27049 18638 27051
rect 18644 27049 18650 27071
rect 18660 27059 18662 27317
rect 18684 27312 18686 27317
rect 18708 27312 18710 27317
rect 18676 27304 18686 27312
rect 18704 27304 18712 27312
rect 18668 27296 18676 27304
rect 18653 27049 18662 27059
rect 18664 27049 18670 27079
rect 18684 27049 18686 27304
rect 18696 27296 18704 27304
rect 18689 27071 18696 27079
rect 18708 27071 18710 27304
rect 18718 27149 18724 27279
rect 18718 27133 18726 27149
rect 18708 27049 18714 27071
rect 18718 27049 18724 27133
rect 18730 27079 18734 27081
rect 18728 27071 18734 27079
rect 18729 27049 18734 27051
rect 18740 27049 18746 27071
rect 18756 27059 18758 27317
rect 18780 27312 18782 27317
rect 18804 27312 18806 27317
rect 18772 27304 18782 27312
rect 18800 27304 18808 27312
rect 18832 27304 18848 27312
rect 18764 27296 18772 27304
rect 18749 27049 18758 27059
rect 18760 27049 18766 27079
rect 18780 27049 18782 27304
rect 18792 27296 18800 27304
rect 18785 27071 18792 27079
rect 18804 27071 18806 27304
rect 18814 27149 18820 27279
rect 18814 27133 18822 27149
rect 18804 27049 18810 27071
rect 18814 27049 18820 27133
rect 18840 27096 18844 27106
rect 18852 27096 18854 27317
rect 18876 27312 18878 27317
rect 18900 27312 18902 27317
rect 18864 27304 18878 27312
rect 18892 27304 18904 27312
rect 18924 27304 18932 27312
rect 18860 27296 18864 27304
rect 18850 27082 18854 27096
rect 18826 27079 18830 27081
rect 18824 27071 18830 27079
rect 18836 27079 18854 27082
rect 18836 27071 18861 27079
rect 18825 27049 18830 27051
rect 18836 27049 18842 27071
rect 18850 27066 18861 27071
rect 18452 27019 18456 27027
rect 18471 27019 18478 27049
rect 18490 27019 18497 27049
rect 18504 27039 18508 27049
rect 18516 27039 18522 27049
rect 18512 27023 18522 27039
rect 18514 27019 18522 27023
rect 18436 26987 18445 27019
rect 18492 26987 18494 27019
rect 18514 27009 18518 27019
rect 18516 27001 18518 27009
rect 18512 26987 18518 27001
rect 18564 26987 18566 27049
rect 18567 27041 18574 27049
rect 18586 27041 18593 27049
rect 18598 27041 18618 27049
rect 18567 27023 18568 27041
rect 18588 26993 18590 27041
rect 18598 27039 18604 27041
rect 18612 27039 18614 27041
rect 18608 27023 18614 27039
rect 18610 27009 18614 27023
rect 18588 26987 18592 26993
rect 18612 26987 18614 27009
rect 18660 26987 18662 27049
rect 18663 27041 18670 27049
rect 18682 27041 18689 27049
rect 18694 27041 18714 27049
rect 18663 27023 18664 27041
rect 18684 26993 18686 27041
rect 18694 27039 18700 27041
rect 18708 27039 18710 27041
rect 18704 27023 18710 27039
rect 18706 27009 18710 27023
rect 18684 26987 18688 26993
rect 18708 26987 18710 27009
rect 18756 26987 18758 27049
rect 18759 27041 18766 27049
rect 18778 27041 18785 27049
rect 18790 27041 18810 27049
rect 18852 27041 18854 27066
rect 18759 27023 18760 27041
rect 18780 26993 18782 27041
rect 18790 27039 18796 27041
rect 18804 27039 18806 27041
rect 18800 27023 18806 27039
rect 18802 27009 18806 27023
rect 18780 26987 18784 26993
rect 18804 26987 18806 27009
rect 18849 27023 18856 27041
rect 18868 27031 18875 27066
rect 18876 27031 18878 27304
rect 18888 27296 18892 27304
rect 18881 27071 18888 27079
rect 18900 27071 18902 27304
rect 18932 27296 18940 27304
rect 18948 27096 18950 27317
rect 18996 27312 18998 27317
rect 19020 27312 19022 27317
rect 19044 27312 19046 27317
rect 18952 27304 18960 27312
rect 18980 27304 18998 27312
rect 19012 27304 19024 27312
rect 19040 27304 19052 27312
rect 18960 27296 18968 27304
rect 18944 27088 18950 27096
rect 18881 27066 18885 27071
rect 18895 27051 18902 27071
rect 18926 27058 18929 27088
rect 18948 27066 18951 27088
rect 18971 27066 18974 27096
rect 18934 27059 18942 27066
rect 18948 27059 18950 27066
rect 18951 27061 18956 27066
rect 18951 27059 18965 27061
rect 18934 27058 18965 27059
rect 18934 27056 18935 27058
rect 18936 27056 18940 27058
rect 18948 27056 18950 27058
rect 18895 27047 18906 27051
rect 18890 27041 18906 27047
rect 18881 27031 18885 27041
rect 18849 26987 18855 27023
rect 18868 27020 18871 27031
rect 18864 27010 18871 27020
rect 18876 27020 18885 27031
rect 18876 27015 18886 27020
rect 18868 26990 18871 27010
rect 18874 27010 18878 27015
rect 18881 27010 18886 27015
rect 18895 27015 18902 27041
rect 18944 27040 18945 27056
rect 18946 27026 18950 27056
rect 18874 27001 18888 27010
rect 18874 26996 18878 27001
rect 18881 26996 18886 27001
rect 18860 26987 18871 26990
rect 18876 26993 18878 26996
rect 18876 26987 18880 26993
rect 18895 26987 18898 27015
rect 18900 26987 18902 27015
rect 18948 27004 18950 27026
rect 18935 26994 18938 26998
rect 18935 26988 18939 26994
rect 18944 26987 18950 27004
rect 18996 26987 18998 27304
rect 19008 27296 19012 27304
rect 19020 27087 19022 27304
rect 19036 27296 19040 27304
rect 19044 27087 19046 27304
rect 19054 27146 19060 27279
rect 19054 27133 19062 27146
rect 19018 27079 19025 27087
rect 19000 27049 19005 27079
rect 19010 27049 19016 27058
rect 19020 27051 19022 27079
rect 19044 27058 19050 27087
rect 19054 27058 19060 27133
rect 19066 27079 19070 27081
rect 19064 27071 19070 27079
rect 19025 27053 19032 27058
rect 19025 27051 19041 27053
rect 19017 27049 19041 27051
rect 19020 27010 19022 27049
rect 19030 27039 19036 27049
rect 19044 27039 19046 27058
rect 19065 27049 19070 27051
rect 19076 27049 19082 27071
rect 19092 27059 19094 27317
rect 19116 27312 19118 27317
rect 19140 27312 19142 27317
rect 19108 27304 19118 27312
rect 19136 27304 19144 27312
rect 19100 27296 19108 27304
rect 19085 27049 19094 27059
rect 19096 27049 19102 27079
rect 19116 27049 19118 27304
rect 19128 27296 19136 27304
rect 19121 27071 19128 27079
rect 19140 27071 19142 27304
rect 19150 27149 19156 27279
rect 19150 27133 19158 27149
rect 19140 27049 19146 27071
rect 19150 27049 19156 27133
rect 19162 27079 19166 27081
rect 19160 27071 19166 27079
rect 19161 27049 19166 27051
rect 19172 27049 19178 27071
rect 19188 27056 19190 27317
rect 19236 27312 19238 27317
rect 19332 27312 19334 27317
rect 19202 27304 19212 27312
rect 19230 27304 19240 27312
rect 19262 27304 19270 27312
rect 19326 27304 19334 27312
rect 19354 27304 19362 27312
rect 19386 27304 19394 27312
rect 19414 27304 19424 27312
rect 19428 27304 19430 27317
rect 19476 27312 19478 27317
rect 19442 27304 19452 27312
rect 19470 27304 19480 27312
rect 19500 27304 19508 27312
rect 19196 27296 19202 27304
rect 19224 27296 19230 27304
rect 19193 27083 19202 27084
rect 19212 27083 19219 27084
rect 19226 27083 19227 27279
rect 19236 27083 19238 27304
rect 19270 27296 19278 27304
rect 19318 27296 19326 27304
rect 19193 27082 19224 27083
rect 19226 27082 19254 27083
rect 19269 27082 19279 27104
rect 19040 27023 19046 27039
rect 19010 26991 19014 27000
rect 19020 26996 19024 27010
rect 19042 27009 19046 27023
rect 19018 26987 19025 26996
rect 19044 26987 19046 27009
rect 19092 26987 19094 27049
rect 19095 27041 19102 27049
rect 19114 27041 19121 27049
rect 19126 27041 19146 27049
rect 19186 27046 19190 27056
rect 19095 27023 19096 27041
rect 19116 26993 19118 27041
rect 19126 27039 19132 27041
rect 19140 27039 19142 27041
rect 19136 27023 19142 27039
rect 19138 27009 19142 27023
rect 19116 26987 19120 26993
rect 19140 26987 19142 27009
rect 19188 26987 19190 27046
rect 19196 27041 19198 27046
rect 19216 27041 19220 27056
rect 19224 27041 19226 27071
rect 19236 27041 19238 27082
rect 19241 27041 19242 27071
rect 19202 27036 19238 27041
rect 19272 27038 19286 27046
rect 19202 27032 19210 27036
rect 19216 27032 19220 27036
rect 19202 27031 19206 27032
rect 19212 27015 19216 27031
rect 19214 27012 19216 27015
rect 19222 27012 19228 27020
rect 19214 27001 19228 27012
rect 19236 27010 19238 27036
rect 19232 26996 19238 27010
rect 19236 26987 19238 26996
rect 19332 27013 19334 27304
rect 19346 27296 19354 27304
rect 19394 27296 19402 27304
rect 19424 27296 19430 27304
rect 19452 27296 19458 27304
rect 19363 27120 19365 27279
rect 19356 27113 19367 27120
rect 19363 27107 19365 27113
rect 19363 27091 19367 27107
rect 19416 27096 19420 27106
rect 19428 27096 19430 27296
rect 19444 27096 19451 27099
rect 19336 27074 19352 27078
rect 19354 27074 19355 27086
rect 19363 27074 19365 27091
rect 19426 27082 19430 27096
rect 19439 27083 19455 27096
rect 19412 27078 19430 27082
rect 19412 27070 19437 27078
rect 19442 27070 19455 27082
rect 19426 27066 19437 27070
rect 19439 27066 19442 27070
rect 19444 27066 19451 27070
rect 19428 27040 19430 27066
rect 19439 27040 19451 27066
rect 19464 27051 19468 27061
rect 19476 27051 19478 27304
rect 19480 27296 19486 27304
rect 19508 27296 19516 27304
rect 19524 27096 19526 27317
rect 19572 27312 19574 27317
rect 19596 27312 19598 27317
rect 19620 27312 19622 27317
rect 19528 27304 19536 27312
rect 19556 27304 19574 27312
rect 19588 27304 19600 27312
rect 19616 27304 19628 27312
rect 19648 27304 19664 27312
rect 19536 27296 19544 27304
rect 19520 27088 19526 27096
rect 19502 27058 19505 27088
rect 19524 27066 19527 27088
rect 19547 27066 19550 27096
rect 19510 27059 19518 27066
rect 19524 27059 19526 27066
rect 19527 27061 19532 27066
rect 19527 27059 19541 27061
rect 19510 27058 19541 27059
rect 19510 27056 19511 27058
rect 19512 27056 19516 27058
rect 19524 27056 19526 27058
rect 19346 27013 19348 27023
rect 19332 27008 19346 27013
rect 19354 27008 19358 27034
rect 19332 26987 19334 27008
rect 19425 26987 19432 27040
rect 19438 27004 19440 27014
rect 19444 27005 19447 27040
rect 19474 27037 19478 27051
rect 19520 27040 19521 27056
rect 19448 27005 19458 27010
rect 19448 27004 19461 27005
rect 19448 26996 19462 27004
rect 19445 26990 19461 26996
rect 19445 26989 19448 26990
rect 19444 26987 19447 26989
rect 19476 26987 19478 27037
rect 19522 27026 19526 27056
rect 19524 27004 19526 27026
rect 19511 26994 19514 26998
rect 19511 26988 19515 26994
rect 19520 26987 19526 27004
rect 19572 26987 19574 27304
rect 19584 27296 19588 27304
rect 19596 27087 19598 27304
rect 19612 27296 19616 27304
rect 19620 27087 19622 27304
rect 19630 27146 19636 27279
rect 19630 27133 19638 27146
rect 19594 27079 19601 27087
rect 19576 27049 19581 27079
rect 19586 27049 19592 27058
rect 19596 27051 19598 27079
rect 19620 27058 19626 27087
rect 19630 27058 19636 27133
rect 19656 27096 19660 27106
rect 19668 27096 19670 27317
rect 19692 27312 19694 27317
rect 19716 27312 19718 27317
rect 19680 27304 19694 27312
rect 19708 27304 19720 27312
rect 19740 27304 19748 27312
rect 19676 27296 19680 27304
rect 19666 27082 19670 27096
rect 19642 27079 19646 27081
rect 19640 27071 19646 27079
rect 19652 27079 19670 27082
rect 19652 27071 19677 27079
rect 19601 27053 19608 27058
rect 19601 27051 19617 27053
rect 19593 27049 19617 27051
rect 19596 27010 19598 27049
rect 19606 27039 19612 27049
rect 19620 27039 19622 27058
rect 19641 27049 19646 27051
rect 19652 27049 19658 27071
rect 19666 27066 19677 27071
rect 19668 27041 19670 27066
rect 19616 27023 19622 27039
rect 19586 26991 19590 27000
rect 19596 26996 19600 27010
rect 19618 27009 19622 27023
rect 19594 26987 19601 26996
rect 19620 26987 19622 27009
rect 19665 27023 19672 27041
rect 19684 27031 19691 27066
rect 19692 27031 19694 27304
rect 19704 27296 19708 27304
rect 19697 27071 19704 27079
rect 19716 27071 19718 27304
rect 19748 27296 19756 27304
rect 19764 27096 19766 27317
rect 19768 27304 19776 27312
rect 19796 27304 19810 27312
rect 19812 27304 19814 27317
rect 19836 27312 19838 27317
rect 19860 27312 19862 27317
rect 19826 27304 19838 27312
rect 19854 27304 19866 27312
rect 19886 27304 19894 27312
rect 19776 27296 19784 27304
rect 19810 27296 19814 27304
rect 19824 27296 19826 27304
rect 19836 27296 19840 27304
rect 19852 27296 19854 27304
rect 19760 27088 19766 27096
rect 19697 27066 19701 27071
rect 19711 27051 19718 27071
rect 19742 27058 19745 27088
rect 19764 27066 19767 27088
rect 19787 27066 19790 27096
rect 19812 27067 19814 27296
rect 19836 27067 19838 27296
rect 19860 27067 19862 27304
rect 19866 27296 19868 27304
rect 19894 27296 19902 27304
rect 19750 27059 19758 27066
rect 19764 27059 19766 27066
rect 19767 27061 19772 27066
rect 19767 27059 19781 27061
rect 19750 27058 19781 27059
rect 19801 27058 19814 27067
rect 19821 27058 19841 27067
rect 19848 27058 19866 27067
rect 19750 27056 19751 27058
rect 19752 27056 19756 27058
rect 19764 27056 19766 27058
rect 19711 27047 19722 27051
rect 19706 27041 19722 27047
rect 19697 27031 19701 27041
rect 19665 26987 19671 27023
rect 19684 27020 19687 27031
rect 19680 27010 19687 27020
rect 19692 27020 19701 27031
rect 19692 27015 19702 27020
rect 19684 26990 19687 27010
rect 19690 27010 19694 27015
rect 19697 27010 19702 27015
rect 19711 27015 19718 27041
rect 19760 27040 19761 27056
rect 19762 27026 19766 27056
rect 19690 27001 19704 27010
rect 19690 26996 19694 27001
rect 19697 26996 19702 27001
rect 19676 26987 19687 26990
rect 19692 26993 19694 26996
rect 19692 26987 19696 26993
rect 19711 26987 19714 27015
rect 19716 26987 19718 27015
rect 19764 27004 19766 27026
rect 19751 26994 19754 26998
rect 19751 26988 19755 26994
rect 19760 26987 19766 27004
rect 19812 27055 19814 27058
rect 19812 27025 19821 27055
rect 19826 27048 19829 27055
rect 19836 27048 19838 27058
rect 19841 27048 19848 27058
rect 19836 27032 19852 27048
rect 19836 27025 19839 27032
rect 19812 26987 19814 27025
rect 19824 27002 19828 27012
rect 19836 27010 19838 27025
rect 19836 27002 19840 27010
rect 19822 26988 19830 26998
rect 19834 26996 19840 27002
rect 19841 26996 19848 27032
rect 19834 26988 19848 26996
rect 19832 26987 19841 26988
rect 19860 26987 19862 27058
rect 19889 27020 19892 27047
rect 19894 27025 19905 27047
rect 19907 27025 19910 27055
rect 19889 27017 19901 27020
rect 19932 26987 19934 27317
rect 19956 27312 19958 27317
rect 19980 27312 19982 27317
rect 19948 27304 19958 27312
rect 19976 27304 19986 27312
rect 19942 27296 19948 27304
rect 19936 27049 19954 27059
rect 19956 27047 19958 27304
rect 19970 27296 19976 27304
rect 19980 27059 19982 27304
rect 19961 27049 19982 27059
rect 19990 27049 19996 27279
rect 20002 27079 20006 27081
rect 20000 27071 20006 27079
rect 20001 27049 20006 27051
rect 20012 27049 20018 27071
rect 20028 27055 20030 27317
rect 20052 27312 20054 27317
rect 20076 27312 20078 27317
rect 20042 27304 20054 27312
rect 20070 27304 20080 27312
rect 20102 27304 20110 27312
rect 20036 27296 20042 27304
rect 20052 27063 20054 27304
rect 20064 27296 20070 27304
rect 20076 27063 20078 27304
rect 20110 27296 20118 27304
rect 20047 27055 20054 27063
rect 19954 27017 19961 27047
rect 19968 27039 19972 27049
rect 19980 27047 19982 27049
rect 19980 27039 19986 27047
rect 19976 27023 19986 27039
rect 19978 27017 19986 27023
rect 20028 27025 20037 27055
rect 20042 27031 20045 27041
rect 20052 27031 20054 27055
rect 20057 27031 20064 27055
rect 20074 27041 20081 27063
rect 20052 27025 20068 27031
rect 20076 27025 20078 27041
rect 20028 27023 20032 27025
rect 19956 26991 19958 27017
rect 19978 27009 19982 27017
rect 19956 26987 19970 26991
rect 19980 26987 19982 27009
rect 20028 26987 20031 27023
rect 20052 27015 20054 27025
rect 20074 27015 20078 27025
rect 20105 27020 20108 27047
rect 20110 27025 20121 27047
rect 20123 27025 20126 27055
rect 20105 27017 20117 27020
rect 20040 27002 20044 27012
rect 20050 27002 20054 27015
rect 20057 27002 20064 27015
rect 20050 27001 20064 27002
rect 20050 26993 20054 27001
rect 20050 26988 20056 26993
rect 20057 26988 20064 27001
rect 20048 26987 20056 26988
rect 20076 26987 20078 27015
rect 20148 26987 20150 27317
rect 20172 27312 20174 27317
rect 20196 27312 20198 27317
rect 20164 27304 20174 27312
rect 20192 27304 20202 27312
rect 20158 27296 20164 27304
rect 20152 27049 20170 27059
rect 20172 27047 20174 27304
rect 20186 27296 20192 27304
rect 20196 27059 20198 27304
rect 20177 27049 20198 27059
rect 20206 27049 20212 27279
rect 20218 27079 20222 27081
rect 20216 27071 20222 27079
rect 20217 27049 20222 27051
rect 20228 27049 20234 27071
rect 20244 27059 20246 27317
rect 20268 27312 20270 27317
rect 20292 27312 20294 27317
rect 20260 27304 20270 27312
rect 20288 27304 20296 27312
rect 20252 27296 20260 27304
rect 20237 27049 20246 27059
rect 20248 27049 20254 27079
rect 20268 27049 20270 27304
rect 20280 27296 20288 27304
rect 20273 27071 20280 27079
rect 20292 27071 20294 27304
rect 20302 27149 20308 27279
rect 20302 27133 20310 27149
rect 20292 27049 20298 27071
rect 20302 27049 20308 27133
rect 20314 27079 20318 27081
rect 20312 27071 20318 27079
rect 20313 27049 20318 27051
rect 20324 27049 20330 27071
rect 20340 27056 20342 27317
rect 20388 27312 20390 27317
rect 20484 27312 20486 27317
rect 20508 27312 20510 27317
rect 20354 27304 20364 27312
rect 20382 27304 20392 27312
rect 20414 27304 20422 27312
rect 20476 27304 20486 27312
rect 20504 27304 20514 27312
rect 20348 27296 20354 27304
rect 20376 27296 20382 27304
rect 20345 27083 20354 27084
rect 20364 27083 20371 27084
rect 20378 27083 20379 27279
rect 20388 27083 20390 27304
rect 20422 27296 20430 27304
rect 20470 27296 20476 27304
rect 20345 27082 20376 27083
rect 20378 27082 20406 27083
rect 20421 27082 20431 27104
rect 20170 27017 20177 27047
rect 20184 27039 20188 27049
rect 20196 27047 20198 27049
rect 20196 27039 20202 27047
rect 20192 27023 20202 27039
rect 20194 27017 20202 27023
rect 20172 26991 20174 27017
rect 20194 27009 20198 27017
rect 20172 26987 20186 26991
rect 20196 26987 20198 27009
rect 20244 26987 20246 27049
rect 20247 27041 20254 27049
rect 20266 27041 20273 27049
rect 20278 27041 20298 27049
rect 20338 27046 20342 27056
rect 20247 27023 20248 27041
rect 20268 26993 20270 27041
rect 20278 27039 20284 27041
rect 20292 27039 20294 27041
rect 20288 27023 20294 27039
rect 20290 27009 20294 27023
rect 20268 26987 20272 26993
rect 20292 26987 20294 27009
rect 20340 26987 20342 27046
rect 20348 27041 20350 27046
rect 20368 27041 20372 27056
rect 20376 27041 20378 27071
rect 20388 27041 20390 27082
rect 20472 27079 20480 27090
rect 20484 27087 20486 27304
rect 20498 27296 20504 27304
rect 20464 27074 20472 27079
rect 20474 27074 20480 27079
rect 20482 27074 20489 27087
rect 20504 27079 20507 27092
rect 20393 27041 20394 27071
rect 20474 27049 20481 27074
rect 20484 27049 20486 27074
rect 20354 27036 20390 27041
rect 20424 27038 20438 27046
rect 20354 27032 20362 27036
rect 20368 27032 20372 27036
rect 20354 27031 20358 27032
rect 20364 27015 20368 27031
rect 20366 27012 20368 27015
rect 20374 27012 20380 27020
rect 20366 27001 20380 27012
rect 20388 27010 20390 27036
rect 20482 27024 20489 27049
rect 20496 27039 20500 27049
rect 20508 27039 20510 27304
rect 20530 27079 20534 27081
rect 20528 27071 20534 27079
rect 20529 27049 20534 27051
rect 20540 27049 20546 27071
rect 20556 27055 20558 27317
rect 20580 27312 20582 27317
rect 20604 27312 20606 27317
rect 20700 27312 20702 27317
rect 20570 27304 20582 27312
rect 20598 27304 20608 27312
rect 20630 27304 20638 27312
rect 20694 27304 20702 27312
rect 20722 27304 20730 27312
rect 20754 27304 20762 27312
rect 20782 27304 20798 27312
rect 20814 27304 20826 27312
rect 20842 27304 20854 27312
rect 20874 27304 20882 27312
rect 20902 27304 20912 27312
rect 20916 27304 20918 27317
rect 20964 27312 20966 27317
rect 20930 27304 20940 27312
rect 20958 27304 20968 27312
rect 20988 27304 20996 27312
rect 20564 27296 20570 27304
rect 20580 27063 20582 27304
rect 20592 27296 20598 27304
rect 20604 27063 20606 27304
rect 20638 27296 20646 27304
rect 20686 27296 20694 27304
rect 20575 27055 20582 27063
rect 20384 26996 20390 27010
rect 20463 27002 20470 27014
rect 20484 27008 20486 27024
rect 20504 27023 20510 27039
rect 20506 27009 20510 27023
rect 20388 26987 20390 26996
rect 20482 26987 20489 27008
rect 20508 26987 20510 27009
rect 20556 27025 20565 27055
rect 20570 27031 20573 27041
rect 20580 27031 20582 27055
rect 20585 27031 20592 27055
rect 20602 27041 20609 27063
rect 20580 27025 20596 27031
rect 20604 27025 20606 27041
rect 20556 27023 20560 27025
rect 20556 26987 20559 27023
rect 20580 27015 20582 27025
rect 20602 27015 20606 27025
rect 20633 27020 20636 27047
rect 20638 27025 20649 27047
rect 20651 27025 20654 27055
rect 20633 27017 20645 27020
rect 20568 27002 20572 27012
rect 20578 27002 20582 27015
rect 20585 27002 20592 27015
rect 20578 27001 20592 27002
rect 20578 26993 20582 27001
rect 20578 26988 20584 26993
rect 20585 26988 20592 27001
rect 20576 26987 20584 26988
rect 20604 26987 20606 27015
rect 20700 27007 20702 27304
rect 20714 27296 20722 27304
rect 20762 27296 20770 27304
rect 20810 27296 20814 27304
rect 20838 27296 20842 27304
rect 20882 27296 20890 27304
rect 20912 27296 20918 27304
rect 20940 27296 20946 27304
rect 20719 27107 20730 27111
rect 20731 27107 20740 27279
rect 20731 27095 20742 27107
rect 20904 27096 20908 27106
rect 20916 27096 20918 27296
rect 20932 27096 20939 27099
rect 20731 27059 20740 27095
rect 20812 27083 20823 27090
rect 20814 27078 20823 27083
rect 20914 27082 20918 27096
rect 20927 27083 20943 27096
rect 20900 27078 20918 27082
rect 20704 27048 20722 27059
rect 20729 27048 20742 27059
rect 20824 27048 20835 27078
rect 20900 27070 20925 27078
rect 20930 27070 20943 27082
rect 20914 27066 20925 27070
rect 20927 27066 20930 27070
rect 20932 27066 20939 27070
rect 20722 27023 20729 27047
rect 20824 27040 20833 27048
rect 20916 27040 20918 27066
rect 20927 27040 20939 27066
rect 20952 27051 20956 27061
rect 20964 27051 20966 27304
rect 20968 27296 20974 27304
rect 20996 27296 21004 27304
rect 21012 27096 21014 27317
rect 21060 27312 21062 27317
rect 21084 27312 21086 27317
rect 21108 27312 21110 27317
rect 21016 27304 21024 27312
rect 21044 27304 21062 27312
rect 21076 27304 21088 27312
rect 21104 27304 21116 27312
rect 21024 27296 21032 27304
rect 21008 27088 21014 27096
rect 20990 27058 20993 27088
rect 21012 27066 21015 27088
rect 21035 27066 21038 27096
rect 20998 27059 21006 27066
rect 21012 27059 21014 27066
rect 21015 27061 21020 27066
rect 21015 27059 21029 27061
rect 20998 27058 21029 27059
rect 20998 27056 20999 27058
rect 21000 27056 21004 27058
rect 21012 27056 21014 27058
rect 20714 27017 20730 27023
rect 20700 26999 20714 27007
rect 20700 26987 20702 26999
rect 20722 26991 20726 27017
rect 20824 27013 20826 27015
rect 20816 27004 20826 27013
rect 20820 26999 20830 27004
rect 20824 26989 20826 26990
rect 20913 26987 20920 27040
rect 20926 27004 20928 27014
rect 20932 27005 20935 27040
rect 20962 27037 20966 27051
rect 21008 27040 21009 27056
rect 20936 27005 20946 27010
rect 20936 27004 20949 27005
rect 20936 26996 20950 27004
rect 20933 26990 20949 26996
rect 20933 26989 20936 26990
rect 20932 26987 20935 26989
rect 20964 26987 20966 27037
rect 21010 27026 21014 27056
rect 21012 27004 21014 27026
rect 20999 26994 21002 26998
rect 20999 26988 21003 26994
rect 21008 26987 21014 27004
rect 21060 26987 21062 27304
rect 21072 27296 21076 27304
rect 21084 27087 21086 27304
rect 21100 27296 21104 27304
rect 21108 27087 21110 27304
rect 21118 27146 21124 27279
rect 21118 27133 21126 27146
rect 21082 27079 21089 27087
rect 21064 27049 21069 27079
rect 21074 27049 21080 27058
rect 21084 27051 21086 27079
rect 21108 27058 21114 27087
rect 21118 27058 21124 27133
rect 21130 27079 21134 27081
rect 21128 27071 21134 27079
rect 21089 27053 21096 27058
rect 21089 27051 21105 27053
rect 21081 27049 21105 27051
rect 21084 27010 21086 27049
rect 21094 27039 21100 27049
rect 21108 27039 21110 27058
rect 21129 27049 21134 27051
rect 21140 27049 21146 27071
rect 21156 27056 21158 27317
rect 21204 27312 21206 27317
rect 21300 27312 21302 27317
rect 21324 27312 21326 27317
rect 21170 27304 21180 27312
rect 21198 27304 21208 27312
rect 21230 27304 21238 27312
rect 21258 27304 21272 27312
rect 21288 27304 21302 27312
rect 21316 27304 21328 27312
rect 21348 27304 21356 27312
rect 21164 27296 21170 27304
rect 21192 27296 21198 27304
rect 21161 27083 21170 27084
rect 21180 27083 21187 27084
rect 21194 27083 21195 27279
rect 21204 27083 21206 27304
rect 21238 27296 21246 27304
rect 21272 27296 21274 27304
rect 21286 27296 21288 27304
rect 21300 27106 21302 27304
rect 21314 27296 21316 27304
rect 21299 27104 21302 27106
rect 21161 27082 21192 27083
rect 21194 27082 21222 27083
rect 21237 27082 21247 27104
rect 21290 27096 21292 27098
rect 21297 27096 21302 27104
rect 21154 27046 21158 27056
rect 21104 27023 21110 27039
rect 21074 26991 21078 27000
rect 21084 26996 21088 27010
rect 21106 27009 21110 27023
rect 21082 26987 21089 26996
rect 21108 26987 21110 27009
rect 21156 26987 21158 27046
rect 21164 27041 21166 27046
rect 21184 27041 21188 27056
rect 21192 27041 21194 27071
rect 21204 27041 21206 27082
rect 21274 27074 21288 27096
rect 21290 27074 21297 27096
rect 21299 27074 21302 27096
rect 21319 27074 21323 27104
rect 21209 27041 21210 27071
rect 21274 27066 21275 27074
rect 21290 27066 21292 27074
rect 21170 27036 21206 27041
rect 21240 27038 21254 27046
rect 21170 27032 21178 27036
rect 21184 27032 21188 27036
rect 21170 27031 21174 27032
rect 21180 27015 21184 27031
rect 21182 27012 21184 27015
rect 21190 27012 21196 27020
rect 21182 27001 21196 27012
rect 21204 27010 21206 27036
rect 21288 27010 21292 27020
rect 21300 27010 21302 27074
rect 21312 27051 21316 27061
rect 21324 27051 21326 27304
rect 21328 27296 21330 27304
rect 21356 27296 21364 27304
rect 21372 27096 21374 27317
rect 21420 27312 21422 27317
rect 21444 27312 21446 27317
rect 21468 27312 21470 27317
rect 21376 27304 21384 27312
rect 21404 27304 21422 27312
rect 21436 27304 21448 27312
rect 21464 27304 21476 27312
rect 21496 27304 21512 27312
rect 21384 27296 21392 27304
rect 21368 27088 21374 27096
rect 21350 27058 21353 27088
rect 21372 27066 21375 27088
rect 21395 27066 21398 27096
rect 21358 27059 21366 27066
rect 21372 27059 21374 27066
rect 21375 27061 21380 27066
rect 21375 27059 21389 27061
rect 21358 27058 21389 27059
rect 21358 27056 21359 27058
rect 21360 27056 21364 27058
rect 21372 27056 21374 27058
rect 21310 27037 21316 27038
rect 21322 27037 21326 27051
rect 21368 27040 21369 27056
rect 21320 27034 21326 27037
rect 21200 26996 21206 27010
rect 21298 27008 21312 27010
rect 21319 27008 21326 27034
rect 21370 27026 21374 27056
rect 21283 26996 21290 27002
rect 21298 26996 21302 27008
rect 21204 26987 21206 26996
rect 21293 26988 21302 26996
rect 21300 26987 21302 26988
rect 21324 26987 21326 27008
rect 21372 27004 21374 27026
rect 21359 26994 21362 26998
rect 21359 26988 21363 26994
rect 21368 26987 21374 27004
rect 21420 26987 21422 27304
rect 21432 27296 21436 27304
rect 21444 27087 21446 27304
rect 21460 27296 21464 27304
rect 21468 27087 21470 27304
rect 21478 27146 21484 27279
rect 21478 27133 21486 27146
rect 21442 27079 21449 27087
rect 21424 27049 21429 27079
rect 21434 27049 21440 27058
rect 21444 27051 21446 27079
rect 21468 27058 21474 27087
rect 21478 27058 21484 27133
rect 21504 27096 21508 27106
rect 21516 27096 21518 27317
rect 21540 27312 21542 27317
rect 21564 27312 21566 27317
rect 21528 27304 21542 27312
rect 21556 27304 21568 27312
rect 21588 27304 21596 27312
rect 21524 27296 21528 27304
rect 21514 27082 21518 27096
rect 21490 27079 21494 27081
rect 21488 27071 21494 27079
rect 21500 27079 21518 27082
rect 21500 27071 21525 27079
rect 21449 27053 21456 27058
rect 21449 27051 21465 27053
rect 21441 27049 21465 27051
rect 21444 27010 21446 27049
rect 21454 27039 21460 27049
rect 21468 27039 21470 27058
rect 21489 27049 21494 27051
rect 21500 27049 21506 27071
rect 21514 27066 21525 27071
rect 21516 27041 21518 27066
rect 21464 27023 21470 27039
rect 21434 26991 21438 27000
rect 21444 26996 21448 27010
rect 21466 27009 21470 27023
rect 21442 26987 21449 26996
rect 21468 26987 21470 27009
rect 21513 27023 21520 27041
rect 21532 27031 21539 27066
rect 21540 27031 21542 27304
rect 21552 27296 21556 27304
rect 21545 27071 21552 27079
rect 21564 27071 21566 27304
rect 21596 27296 21604 27304
rect 21612 27096 21614 27317
rect 21616 27304 21624 27312
rect 21644 27304 21658 27312
rect 21660 27304 21662 27317
rect 21684 27312 21686 27317
rect 21708 27312 21710 27317
rect 21674 27304 21686 27312
rect 21702 27304 21714 27312
rect 21734 27304 21742 27312
rect 21762 27304 21778 27312
rect 21624 27296 21632 27304
rect 21658 27296 21662 27304
rect 21672 27296 21674 27304
rect 21684 27296 21688 27304
rect 21700 27296 21702 27304
rect 21608 27088 21614 27096
rect 21545 27066 21549 27071
rect 21559 27051 21566 27071
rect 21590 27058 21593 27088
rect 21612 27066 21615 27088
rect 21635 27066 21638 27096
rect 21660 27067 21662 27296
rect 21684 27067 21686 27296
rect 21708 27067 21710 27304
rect 21714 27296 21716 27304
rect 21742 27296 21750 27304
rect 21598 27059 21606 27066
rect 21612 27059 21614 27066
rect 21615 27061 21620 27066
rect 21615 27059 21629 27061
rect 21598 27058 21629 27059
rect 21649 27058 21662 27067
rect 21669 27058 21689 27067
rect 21696 27058 21714 27067
rect 21598 27056 21599 27058
rect 21600 27056 21604 27058
rect 21612 27056 21614 27058
rect 21559 27047 21570 27051
rect 21554 27041 21570 27047
rect 21545 27031 21549 27041
rect 21513 26987 21519 27023
rect 21532 27020 21535 27031
rect 21528 27010 21535 27020
rect 21540 27020 21549 27031
rect 21540 27015 21550 27020
rect 21532 26990 21535 27010
rect 21538 27010 21542 27015
rect 21545 27010 21550 27015
rect 21559 27015 21566 27041
rect 21608 27040 21609 27056
rect 21610 27026 21614 27056
rect 21538 27001 21552 27010
rect 21538 26996 21542 27001
rect 21545 26996 21550 27001
rect 21524 26987 21535 26990
rect 21540 26993 21542 26996
rect 21540 26987 21544 26993
rect 21559 26987 21562 27015
rect 21564 26987 21566 27015
rect 21612 27004 21614 27026
rect 21599 26994 21602 26998
rect 21599 26988 21603 26994
rect 21608 26987 21614 27004
rect 21660 27055 21662 27058
rect 21660 27025 21669 27055
rect 21674 27048 21677 27055
rect 21684 27048 21686 27058
rect 21689 27048 21696 27058
rect 21684 27032 21700 27048
rect 21684 27025 21687 27032
rect 21660 26987 21662 27025
rect 21672 27002 21676 27012
rect 21684 27010 21686 27025
rect 21684 27002 21688 27010
rect 21670 26988 21678 26998
rect 21682 26996 21688 27002
rect 21689 26996 21696 27032
rect 21682 26988 21696 26996
rect 21680 26987 21689 26988
rect 21708 26987 21710 27058
rect 21780 27055 21782 27317
rect 21804 27312 21806 27317
rect 21828 27312 21830 27317
rect 21794 27304 21806 27312
rect 21822 27304 21834 27312
rect 21854 27304 21862 27312
rect 21882 27304 21898 27312
rect 21790 27296 21794 27304
rect 21737 27020 21740 27047
rect 21742 27025 21753 27047
rect 21755 27025 21758 27055
rect 21780 27025 21789 27055
rect 21804 27025 21806 27304
rect 21818 27296 21822 27304
rect 21809 27025 21816 27055
rect 21828 27047 21830 27304
rect 21862 27296 21870 27304
rect 21900 27055 21902 27317
rect 21924 27312 21926 27317
rect 21948 27312 21950 27317
rect 21914 27304 21926 27312
rect 21942 27304 21954 27312
rect 21974 27304 21982 27312
rect 22002 27304 22016 27312
rect 21910 27296 21914 27304
rect 21737 27017 21749 27020
rect 21780 26987 21782 27025
rect 21799 27017 21806 27025
rect 21826 27017 21833 27047
rect 21857 27020 21860 27047
rect 21862 27025 21873 27047
rect 21875 27025 21878 27055
rect 21900 27025 21909 27055
rect 21924 27025 21926 27304
rect 21938 27296 21942 27304
rect 21929 27025 21936 27055
rect 21948 27047 21950 27304
rect 21982 27296 21990 27304
rect 22016 27296 22018 27304
rect 22008 27096 22012 27106
rect 22020 27096 22022 27317
rect 22044 27312 22046 27317
rect 22068 27312 22070 27317
rect 22032 27304 22046 27312
rect 22060 27304 22072 27312
rect 22092 27304 22100 27312
rect 22030 27296 22032 27304
rect 22018 27066 22022 27096
rect 21857 27017 21869 27020
rect 21792 27002 21796 27012
rect 21804 27002 21806 27017
rect 21809 27007 21816 27017
rect 21802 26988 21816 27002
rect 21826 26991 21830 27017
rect 21803 26987 21816 26988
rect 21828 26987 21830 26991
rect 21900 26987 21902 27025
rect 21919 27017 21926 27025
rect 21946 27017 21953 27047
rect 21977 27020 21980 27047
rect 21982 27025 21993 27047
rect 21995 27025 21998 27055
rect 21977 27017 21989 27020
rect 21912 27002 21916 27012
rect 21924 27002 21926 27017
rect 21929 27007 21936 27017
rect 21922 26988 21936 27002
rect 21946 26991 21950 27017
rect 22020 27004 22022 27066
rect 22036 27055 22043 27065
rect 22036 27047 22039 27055
rect 22036 27020 22043 27047
rect 22032 27017 22043 27020
rect 22032 27010 22039 27017
rect 22044 27010 22046 27304
rect 22058 27296 22060 27304
rect 22068 27104 22070 27304
rect 22072 27296 22074 27304
rect 22100 27296 22108 27304
rect 22063 27096 22070 27104
rect 22116 27096 22118 27317
rect 22120 27304 22128 27312
rect 22148 27304 22162 27312
rect 22164 27304 22166 27317
rect 22188 27312 22190 27317
rect 22212 27312 22214 27317
rect 22701 27314 22717 27317
rect 22178 27304 22190 27312
rect 22206 27304 22218 27312
rect 22238 27304 22246 27312
rect 22266 27304 22282 27312
rect 22299 27304 22310 27312
rect 22328 27304 22338 27312
rect 22359 27304 22369 27312
rect 22388 27304 22397 27312
rect 22417 27304 22425 27312
rect 22445 27304 22453 27312
rect 22473 27304 22482 27312
rect 22501 27304 22510 27312
rect 22530 27304 22538 27312
rect 22558 27304 22566 27312
rect 22586 27304 22594 27312
rect 22614 27304 22622 27312
rect 22642 27304 22650 27312
rect 22670 27304 22678 27312
rect 22864 27309 22866 27317
rect 22726 27304 22734 27309
rect 22754 27304 22762 27309
rect 22128 27296 22136 27304
rect 22162 27296 22166 27304
rect 22176 27296 22178 27304
rect 22188 27296 22192 27304
rect 22204 27296 22206 27304
rect 22058 27095 22074 27096
rect 22049 27047 22053 27055
rect 22056 27051 22060 27061
rect 22063 27051 22066 27065
rect 22068 27051 22070 27095
rect 22112 27088 22118 27096
rect 22094 27058 22097 27088
rect 22116 27066 22119 27088
rect 22139 27066 22142 27096
rect 22164 27067 22166 27296
rect 22188 27067 22190 27296
rect 22212 27067 22214 27304
rect 22218 27296 22220 27304
rect 22246 27296 22254 27304
rect 22294 27296 22299 27304
rect 22322 27296 22328 27304
rect 22369 27296 22375 27304
rect 22397 27296 22404 27304
rect 22425 27296 22433 27304
rect 22453 27296 22461 27304
rect 22482 27296 22489 27304
rect 22510 27296 22517 27304
rect 22538 27296 22546 27304
rect 22566 27296 22574 27304
rect 22594 27296 22602 27304
rect 22622 27296 22630 27304
rect 22650 27296 22658 27304
rect 22678 27296 22686 27304
rect 22734 27293 22742 27304
rect 22762 27294 22770 27304
rect 22810 27301 22818 27309
rect 22838 27301 22846 27309
rect 22864 27301 22874 27309
rect 22894 27301 22904 27312
rect 22922 27301 22932 27312
rect 22950 27301 22960 27312
rect 22980 27304 22988 27312
rect 22818 27294 22826 27301
rect 22846 27294 22854 27301
rect 22754 27293 22770 27294
rect 22810 27293 22826 27294
rect 22838 27293 22854 27294
rect 22864 27294 22866 27301
rect 22874 27294 22882 27301
rect 22904 27296 22910 27301
rect 22932 27296 22938 27301
rect 22960 27296 22966 27301
rect 22988 27296 22996 27304
rect 22864 27293 22882 27294
rect 22894 27293 22902 27294
rect 22414 27279 22547 27287
rect 22552 27279 22605 27287
rect 22562 27261 22566 27270
rect 22630 27269 22637 27278
rect 22613 27257 22619 27262
rect 22638 27257 22647 27269
rect 22609 27252 22613 27257
rect 22638 27253 22654 27257
rect 22655 27253 22658 27257
rect 22322 27080 22328 27248
rect 22387 27238 22393 27246
rect 22424 27238 22435 27242
rect 22397 27230 22403 27238
rect 22378 27210 22393 27230
rect 22424 27227 22437 27238
rect 22462 27230 22469 27238
rect 22453 27227 22469 27230
rect 22500 27227 22510 27249
rect 22378 27200 22397 27210
rect 22404 27200 22423 27210
rect 22397 27198 22403 27200
rect 22444 27198 22447 27227
rect 22453 27208 22461 27227
rect 22527 27219 22533 27249
rect 22568 27219 22573 27249
rect 22609 27227 22610 27252
rect 22642 27227 22649 27253
rect 22449 27200 22462 27208
rect 22397 27192 22404 27198
rect 22397 27190 22411 27192
rect 22397 27185 22420 27190
rect 22386 27160 22393 27170
rect 22404 27168 22420 27185
rect 22430 27168 22437 27198
rect 22451 27195 22469 27198
rect 22444 27166 22451 27190
rect 22459 27168 22469 27195
rect 22642 27193 22647 27227
rect 22679 27221 22688 27222
rect 22685 27219 22688 27221
rect 22520 27190 22526 27193
rect 22404 27160 22458 27166
rect 22459 27160 22468 27168
rect 22485 27163 22501 27190
rect 22520 27163 22523 27190
rect 22526 27163 22527 27190
rect 22561 27185 22566 27193
rect 22561 27163 22577 27185
rect 22583 27163 22591 27185
rect 22485 27160 22492 27163
rect 22527 27160 22533 27163
rect 22394 27153 22403 27160
rect 22561 27155 22599 27163
rect 22630 27155 22637 27185
rect 22642 27163 22649 27193
rect 22864 27186 22866 27293
rect 22651 27163 22658 27185
rect 22663 27163 22667 27185
rect 22651 27155 22668 27163
rect 22752 27156 22764 27172
rect 22332 27100 22338 27111
rect 22394 27070 22401 27153
rect 22444 27122 22447 27133
rect 22526 27132 22533 27148
rect 22535 27133 22565 27140
rect 22642 27130 22647 27155
rect 22843 27148 22844 27164
rect 22859 27162 22867 27186
rect 22658 27133 22672 27140
rect 22444 27092 22451 27122
rect 22561 27100 22566 27130
rect 22602 27100 22609 27130
rect 22630 27100 22631 27122
rect 22642 27100 22649 27130
rect 22615 27092 22637 27100
rect 22663 27092 22670 27122
rect 22721 27106 22734 27122
rect 22739 27106 22743 27136
rect 22821 27110 22837 27126
rect 22830 27101 22837 27110
rect 22842 27106 22844 27128
rect 22859 27106 22868 27146
rect 22918 27106 22936 27108
rect 22897 27102 22906 27106
rect 22913 27102 22936 27106
rect 22813 27098 22817 27101
rect 22828 27098 22844 27101
rect 22918 27098 22936 27102
rect 22943 27098 22961 27108
rect 22444 27070 22447 27092
rect 22642 27083 22647 27092
rect 22102 27059 22110 27066
rect 22116 27059 22118 27066
rect 22119 27061 22124 27066
rect 22119 27059 22133 27061
rect 22102 27058 22133 27059
rect 22153 27058 22166 27067
rect 22173 27058 22193 27067
rect 22200 27058 22218 27067
rect 22378 27062 22430 27070
rect 22437 27062 22449 27070
rect 22493 27062 22529 27070
rect 22102 27056 22103 27058
rect 22104 27056 22108 27058
rect 22116 27056 22118 27058
rect 22063 27047 22070 27051
rect 22063 27021 22074 27047
rect 22112 27040 22113 27056
rect 22114 27026 22118 27056
rect 22063 27020 22070 27021
rect 21923 26987 21936 26988
rect 21948 26987 21950 26991
rect 22017 26987 22022 27004
rect 22036 26987 22039 27010
rect 22042 27007 22046 27010
rect 22049 27007 22054 27020
rect 22058 27017 22070 27020
rect 22042 26996 22056 27007
rect 22044 26987 22053 26996
rect 22063 26991 22070 27017
rect 22116 27004 22118 27026
rect 22063 26987 22066 26991
rect 22068 26987 22070 26991
rect 22103 26994 22106 26998
rect 22103 26988 22107 26994
rect 22112 26987 22118 27004
rect 22164 27055 22166 27058
rect 22164 27025 22173 27055
rect 22178 27048 22181 27055
rect 22188 27048 22190 27058
rect 22193 27048 22200 27058
rect 22188 27032 22204 27048
rect 22188 27025 22191 27032
rect 22164 26987 22166 27025
rect 22176 27002 22180 27012
rect 22188 27010 22190 27025
rect 22188 27002 22192 27010
rect 22174 26988 22182 26998
rect 22186 26996 22192 27002
rect 22193 26996 22200 27032
rect 22186 26988 22200 26996
rect 22184 26987 22193 26988
rect 22212 26987 22214 27058
rect 22241 27020 22244 27047
rect 22246 27025 22257 27047
rect 22259 27025 22262 27055
rect 22241 27017 22253 27020
rect 22320 27017 22325 27047
rect 22394 26987 22401 27062
rect 22444 27060 22447 27062
rect 22430 27052 22437 27060
rect 22430 27030 22446 27052
rect 22462 27030 22469 27060
rect 22520 27052 22526 27060
rect 22561 27052 22566 27060
rect 22642 27057 22649 27083
rect 22642 27052 22647 27057
rect 22503 27030 22515 27052
rect 22520 27030 22521 27052
rect 22526 27030 22527 27052
rect 22566 27030 22568 27052
rect 22579 27030 22594 27052
rect 22527 27027 22533 27030
rect 22499 27022 22533 27027
rect 22568 27022 22573 27030
rect 22630 27022 22637 27052
rect 22663 27026 22670 27052
rect 22672 27047 22680 27082
rect 22751 27027 22755 27043
rect 22756 27041 22767 27043
rect 22803 27041 22809 27098
rect 22822 27071 22823 27073
rect 22830 27071 22836 27098
rect 22936 27096 22941 27098
rect 22951 27096 22953 27098
rect 23004 27096 23006 27317
rect 23008 27304 23016 27312
rect 23036 27304 23048 27312
rect 23052 27304 23054 27317
rect 23076 27312 23078 27317
rect 23100 27312 23102 27317
rect 23064 27304 23078 27312
rect 23092 27304 23104 27312
rect 23124 27304 23132 27312
rect 23016 27296 23024 27304
rect 23048 27296 23054 27304
rect 23040 27096 23044 27106
rect 23052 27096 23054 27296
rect 23076 27296 23080 27304
rect 22879 27083 22882 27091
rect 22889 27081 22892 27083
rect 22819 27041 22826 27071
rect 22832 27041 22837 27063
rect 22842 27041 22848 27063
rect 22850 27041 22857 27071
rect 22859 27041 22868 27081
rect 22869 27041 22875 27063
rect 22877 27041 22884 27071
rect 22889 27041 22895 27081
rect 22906 27075 22913 27096
rect 22936 27075 22943 27096
rect 23000 27088 23006 27096
rect 22906 27073 22924 27075
rect 22905 27066 22924 27073
rect 22931 27066 22951 27075
rect 22958 27066 22973 27075
rect 22905 27063 22915 27066
rect 22936 27063 22941 27066
rect 22951 27063 22953 27066
rect 22766 27035 22767 27041
rect 22830 27033 22837 27041
rect 22859 27033 22867 27041
rect 22654 27022 22670 27026
rect 22444 26987 22447 27022
rect 22515 26999 22519 27015
rect 22520 26987 22523 26995
rect 22579 26991 22595 26993
rect 22642 26987 22647 27022
rect 22830 27018 22836 27033
rect 22729 27008 22737 27018
rect 22830 27013 22845 27018
rect 22739 27008 22748 27011
rect 22739 26992 22747 27008
rect 22748 26995 22755 27008
rect 22830 27003 22836 27013
rect 22860 26987 22867 27033
rect 22905 27013 22909 27063
rect 22918 27033 22931 27063
rect 22951 27051 22958 27063
rect 22982 27058 22985 27088
rect 23004 27066 23007 27088
rect 23027 27066 23030 27096
rect 23050 27066 23061 27096
rect 22990 27059 22998 27066
rect 23004 27059 23006 27066
rect 23007 27061 23012 27066
rect 23007 27059 23021 27061
rect 22990 27058 23021 27059
rect 22990 27056 22991 27058
rect 22992 27056 22996 27058
rect 23004 27056 23006 27058
rect 22951 27033 22961 27051
rect 23000 27040 23001 27056
rect 22921 27000 22925 27033
rect 22936 27020 22941 27033
rect 22936 26996 22942 27020
rect 22951 26987 22953 27033
rect 23002 27026 23006 27056
rect 23052 27053 23054 27066
rect 23004 27004 23006 27026
rect 23049 27013 23054 27053
rect 23068 27048 23075 27066
rect 23076 27048 23078 27296
rect 23081 27088 23088 27096
rect 23100 27088 23102 27304
rect 23104 27296 23108 27304
rect 23132 27296 23140 27304
rect 23148 27096 23150 27317
rect 23196 27312 23198 27317
rect 23220 27312 23222 27317
rect 23244 27312 23246 27317
rect 23152 27304 23160 27312
rect 23180 27304 23198 27312
rect 23212 27304 23224 27312
rect 23240 27304 23252 27312
rect 23160 27296 23168 27304
rect 23144 27088 23150 27096
rect 23081 27066 23085 27088
rect 23095 27061 23102 27088
rect 23088 27058 23106 27061
rect 23126 27058 23129 27088
rect 23148 27066 23151 27088
rect 23171 27066 23174 27096
rect 23134 27059 23142 27066
rect 23148 27059 23150 27066
rect 23151 27061 23156 27066
rect 23151 27059 23165 27061
rect 23134 27058 23165 27059
rect 23081 27048 23085 27058
rect 23088 27051 23092 27058
rect 23068 27020 23071 27048
rect 22991 26994 22994 26998
rect 22991 26988 22995 26994
rect 23000 26987 23006 27004
rect 23052 26987 23054 27013
rect 23064 27010 23071 27020
rect 23076 27032 23085 27048
rect 23086 27037 23092 27047
rect 23076 27020 23078 27032
rect 23081 27020 23085 27032
rect 23095 27021 23102 27058
rect 23134 27056 23135 27058
rect 23136 27056 23140 27058
rect 23148 27056 23150 27058
rect 23144 27040 23145 27056
rect 23146 27026 23150 27056
rect 23076 27018 23092 27020
rect 23076 27010 23078 27018
rect 23068 26996 23071 27010
rect 23074 26996 23080 27010
rect 23081 26996 23086 27018
rect 23055 26987 23071 26996
rect 23076 26987 23080 26996
rect 23095 26987 23098 27021
rect 23100 26987 23102 27021
rect 23148 27004 23150 27026
rect 23135 26994 23138 26998
rect 23135 26988 23139 26994
rect 23144 26987 23150 27004
rect 23196 26987 23198 27304
rect 23208 27296 23212 27304
rect 23220 27087 23222 27304
rect 23236 27296 23240 27304
rect 23244 27087 23246 27304
rect 23254 27146 23260 27279
rect 23254 27133 23262 27146
rect 23218 27079 23225 27087
rect 23200 27049 23205 27079
rect 23210 27049 23216 27058
rect 23220 27051 23222 27079
rect 23244 27058 23250 27087
rect 23254 27058 23260 27133
rect 23266 27079 23270 27081
rect 23264 27071 23270 27079
rect 23225 27053 23232 27058
rect 23225 27051 23241 27053
rect 23217 27049 23241 27051
rect 23220 27010 23222 27049
rect 23230 27039 23236 27049
rect 23244 27039 23246 27058
rect 23265 27049 23270 27051
rect 23276 27049 23282 27071
rect 23292 27059 23294 27317
rect 23316 27312 23318 27317
rect 23340 27312 23342 27317
rect 23308 27304 23318 27312
rect 23336 27304 23344 27312
rect 23368 27304 23384 27312
rect 23300 27296 23308 27304
rect 23285 27049 23294 27059
rect 23296 27049 23302 27079
rect 23316 27049 23318 27304
rect 23328 27296 23336 27304
rect 23321 27071 23328 27079
rect 23340 27071 23342 27304
rect 23350 27149 23356 27279
rect 23350 27133 23358 27149
rect 23340 27049 23346 27071
rect 23350 27049 23356 27133
rect 23376 27096 23380 27106
rect 23388 27096 23390 27317
rect 23412 27312 23414 27317
rect 23436 27312 23438 27317
rect 23400 27304 23414 27312
rect 23428 27304 23440 27312
rect 23460 27304 23468 27312
rect 23396 27296 23400 27304
rect 23386 27082 23390 27096
rect 23362 27079 23366 27081
rect 23360 27071 23366 27079
rect 23372 27079 23390 27082
rect 23372 27071 23397 27079
rect 23361 27049 23366 27051
rect 23372 27049 23378 27071
rect 23386 27066 23397 27071
rect 23240 27023 23246 27039
rect 23210 26991 23214 27000
rect 23220 26996 23224 27010
rect 23242 27009 23246 27023
rect 23218 26987 23225 26996
rect 23244 26987 23246 27009
rect 23292 26987 23294 27049
rect 23295 27041 23302 27049
rect 23314 27041 23321 27049
rect 23326 27041 23346 27049
rect 23388 27041 23390 27066
rect 23295 27023 23296 27041
rect 23316 26993 23318 27041
rect 23326 27039 23332 27041
rect 23340 27039 23342 27041
rect 23336 27023 23342 27039
rect 23338 27009 23342 27023
rect 23316 26987 23320 26993
rect 23340 26987 23342 27009
rect 23385 27023 23392 27041
rect 23404 27031 23411 27066
rect 23412 27031 23414 27304
rect 23424 27296 23428 27304
rect 23417 27071 23424 27079
rect 23436 27071 23438 27304
rect 23468 27296 23476 27304
rect 23484 27096 23486 27317
rect 23532 27312 23534 27317
rect 23556 27312 23558 27317
rect 23580 27312 23582 27317
rect 23488 27304 23496 27312
rect 23516 27304 23534 27312
rect 23548 27304 23560 27312
rect 23576 27304 23588 27312
rect 23496 27296 23504 27304
rect 23480 27088 23486 27096
rect 23417 27066 23421 27071
rect 23431 27051 23438 27071
rect 23462 27058 23465 27088
rect 23484 27066 23487 27088
rect 23507 27066 23510 27096
rect 23470 27059 23478 27066
rect 23484 27059 23486 27066
rect 23487 27061 23492 27066
rect 23487 27059 23501 27061
rect 23470 27058 23501 27059
rect 23470 27056 23471 27058
rect 23472 27056 23476 27058
rect 23484 27056 23486 27058
rect 23431 27047 23442 27051
rect 23426 27041 23442 27047
rect 23417 27031 23421 27041
rect 23385 26987 23391 27023
rect 23404 27020 23407 27031
rect 23400 27010 23407 27020
rect 23412 27020 23421 27031
rect 23412 27015 23422 27020
rect 23404 26990 23407 27010
rect 23410 27010 23414 27015
rect 23417 27010 23422 27015
rect 23431 27015 23438 27041
rect 23480 27040 23481 27056
rect 23482 27026 23486 27056
rect 23410 27001 23424 27010
rect 23410 26996 23414 27001
rect 23417 26996 23422 27001
rect 23396 26987 23407 26990
rect 23412 26993 23414 26996
rect 23412 26987 23416 26993
rect 23431 26987 23434 27015
rect 23436 26987 23438 27015
rect 23484 27004 23486 27026
rect 23471 26994 23474 26998
rect 23471 26988 23475 26994
rect 23480 26987 23486 27004
rect 23532 26987 23534 27304
rect 23544 27296 23548 27304
rect 23556 27087 23558 27304
rect 23572 27296 23576 27304
rect 23580 27087 23582 27304
rect 23590 27146 23596 27279
rect 23590 27133 23598 27146
rect 23554 27079 23561 27087
rect 23536 27049 23541 27079
rect 23546 27049 23552 27058
rect 23556 27051 23558 27079
rect 23580 27058 23586 27087
rect 23590 27058 23596 27133
rect 23602 27079 23606 27081
rect 23600 27071 23606 27079
rect 23561 27053 23568 27058
rect 23561 27051 23577 27053
rect 23553 27049 23577 27051
rect 23556 27010 23558 27049
rect 23566 27039 23572 27049
rect 23580 27039 23582 27058
rect 23601 27049 23606 27051
rect 23612 27049 23618 27071
rect 23628 27059 23630 27317
rect 23652 27312 23654 27317
rect 23676 27312 23678 27317
rect 23644 27304 23654 27312
rect 23672 27304 23680 27312
rect 23704 27304 23720 27312
rect 23636 27296 23644 27304
rect 23621 27049 23630 27059
rect 23632 27049 23638 27079
rect 23652 27049 23654 27304
rect 23664 27296 23672 27304
rect 23657 27071 23664 27079
rect 23676 27071 23678 27304
rect 23686 27149 23692 27279
rect 23686 27133 23694 27149
rect 23676 27049 23682 27071
rect 23686 27049 23692 27133
rect 23712 27096 23716 27106
rect 23724 27096 23726 27317
rect 23748 27312 23750 27317
rect 23772 27312 23774 27317
rect 23736 27304 23750 27312
rect 23764 27304 23776 27312
rect 23796 27304 23804 27312
rect 23732 27296 23736 27304
rect 23722 27082 23726 27096
rect 23698 27079 23702 27081
rect 23696 27071 23702 27079
rect 23708 27079 23726 27082
rect 23708 27071 23733 27079
rect 23697 27049 23702 27051
rect 23708 27049 23714 27071
rect 23722 27066 23733 27071
rect 23576 27023 23582 27039
rect 23546 26991 23550 27000
rect 23556 26996 23560 27010
rect 23578 27009 23582 27023
rect 23554 26987 23561 26996
rect 23580 26987 23582 27009
rect 23628 26987 23630 27049
rect 23631 27041 23638 27049
rect 23650 27041 23657 27049
rect 23662 27041 23682 27049
rect 23724 27041 23726 27066
rect 23631 27023 23632 27041
rect 23652 26993 23654 27041
rect 23662 27039 23668 27041
rect 23676 27039 23678 27041
rect 23672 27023 23678 27039
rect 23674 27009 23678 27023
rect 23652 26987 23656 26993
rect 23676 26987 23678 27009
rect 23721 27023 23728 27041
rect 23740 27031 23747 27066
rect 23748 27031 23750 27304
rect 23760 27296 23764 27304
rect 23753 27071 23760 27079
rect 23772 27071 23774 27304
rect 23804 27296 23812 27304
rect 23820 27096 23822 27317
rect 23824 27304 23832 27312
rect 23852 27304 23866 27312
rect 23868 27304 23870 27317
rect 23892 27312 23894 27317
rect 23916 27312 23918 27317
rect 23882 27304 23894 27312
rect 23910 27304 23922 27312
rect 23942 27304 23950 27312
rect 23832 27296 23840 27304
rect 23866 27296 23870 27304
rect 23880 27296 23882 27304
rect 23892 27296 23896 27304
rect 23908 27296 23910 27304
rect 23816 27088 23822 27096
rect 23753 27066 23757 27071
rect 23767 27051 23774 27071
rect 23798 27058 23801 27088
rect 23820 27066 23823 27088
rect 23843 27066 23846 27096
rect 23868 27067 23870 27296
rect 23892 27067 23894 27296
rect 23916 27067 23918 27304
rect 23922 27296 23924 27304
rect 23950 27296 23958 27304
rect 23806 27059 23814 27066
rect 23820 27059 23822 27066
rect 23823 27061 23828 27066
rect 23823 27059 23837 27061
rect 23806 27058 23837 27059
rect 23857 27058 23870 27067
rect 23877 27058 23897 27067
rect 23904 27058 23922 27067
rect 23806 27056 23807 27058
rect 23808 27056 23812 27058
rect 23820 27056 23822 27058
rect 23767 27047 23778 27051
rect 23762 27041 23778 27047
rect 23753 27031 23757 27041
rect 23721 26987 23727 27023
rect 23740 27020 23743 27031
rect 23736 27010 23743 27020
rect 23748 27020 23757 27031
rect 23748 27015 23758 27020
rect 23740 26990 23743 27010
rect 23746 27010 23750 27015
rect 23753 27010 23758 27015
rect 23767 27015 23774 27041
rect 23816 27040 23817 27056
rect 23818 27026 23822 27056
rect 23746 27001 23760 27010
rect 23746 26996 23750 27001
rect 23753 26996 23758 27001
rect 23732 26987 23743 26990
rect 23748 26993 23750 26996
rect 23748 26987 23752 26993
rect 23767 26987 23770 27015
rect 23772 26987 23774 27015
rect 23820 27004 23822 27026
rect 23807 26994 23810 26998
rect 23807 26988 23811 26994
rect 23816 26987 23822 27004
rect 23868 27055 23870 27058
rect 23868 27025 23877 27055
rect 23882 27048 23885 27055
rect 23892 27048 23894 27058
rect 23897 27048 23904 27058
rect 23892 27032 23908 27048
rect 23892 27025 23895 27032
rect 23868 26987 23870 27025
rect 23880 27002 23884 27012
rect 23892 27010 23894 27025
rect 23892 27002 23896 27010
rect 23878 26988 23886 26998
rect 23890 26996 23896 27002
rect 23897 26996 23904 27032
rect 23890 26988 23904 26996
rect 23888 26987 23897 26988
rect 23916 26987 23918 27058
rect 23945 27020 23948 27047
rect 23950 27025 23961 27047
rect 23963 27025 23966 27055
rect 23945 27017 23957 27020
rect 23988 26987 23990 27317
rect 24012 27312 24014 27317
rect 24036 27312 24038 27317
rect 24004 27304 24014 27312
rect 24032 27304 24042 27312
rect 23998 27296 24004 27304
rect 23992 27049 24010 27059
rect 24012 27047 24014 27304
rect 24026 27296 24032 27304
rect 24036 27059 24038 27304
rect 24017 27049 24038 27059
rect 24046 27049 24052 27279
rect 24058 27079 24062 27081
rect 24056 27071 24062 27079
rect 24057 27049 24062 27051
rect 24068 27049 24074 27071
rect 24084 27056 24086 27317
rect 24132 27312 24134 27317
rect 24228 27312 24230 27317
rect 24252 27312 24254 27317
rect 24098 27304 24108 27312
rect 24126 27304 24136 27312
rect 24158 27304 24166 27312
rect 24186 27304 24200 27312
rect 24216 27304 24230 27312
rect 24244 27304 24256 27312
rect 24276 27304 24284 27312
rect 24092 27296 24098 27304
rect 24120 27296 24126 27304
rect 24089 27083 24098 27084
rect 24108 27083 24115 27084
rect 24122 27083 24123 27279
rect 24132 27083 24134 27304
rect 24166 27296 24174 27304
rect 24200 27296 24202 27304
rect 24214 27296 24216 27304
rect 24228 27106 24230 27304
rect 24242 27296 24244 27304
rect 24227 27104 24230 27106
rect 24089 27082 24120 27083
rect 24122 27082 24150 27083
rect 24165 27082 24175 27104
rect 24218 27096 24220 27098
rect 24225 27096 24230 27104
rect 24010 27017 24017 27047
rect 24024 27039 24028 27049
rect 24036 27047 24038 27049
rect 24036 27039 24042 27047
rect 24082 27046 24086 27056
rect 24032 27023 24042 27039
rect 24034 27017 24042 27023
rect 24012 26991 24014 27017
rect 24034 27009 24038 27017
rect 24012 26987 24026 26991
rect 24036 26987 24038 27009
rect 24084 26987 24086 27046
rect 24092 27041 24094 27046
rect 24112 27041 24116 27056
rect 24120 27041 24122 27071
rect 24132 27041 24134 27082
rect 24202 27074 24216 27096
rect 24218 27074 24225 27096
rect 24227 27074 24230 27096
rect 24247 27074 24251 27104
rect 24137 27041 24138 27071
rect 24202 27066 24203 27074
rect 24218 27066 24220 27074
rect 24098 27036 24134 27041
rect 24168 27038 24182 27046
rect 24098 27032 24106 27036
rect 24112 27032 24116 27036
rect 24098 27031 24102 27032
rect 24108 27015 24112 27031
rect 24110 27012 24112 27015
rect 24118 27012 24124 27020
rect 24110 27001 24124 27012
rect 24132 27010 24134 27036
rect 24216 27010 24220 27020
rect 24228 27010 24230 27074
rect 24240 27051 24244 27061
rect 24252 27051 24254 27304
rect 24256 27296 24258 27304
rect 24284 27296 24292 27304
rect 24300 27096 24302 27317
rect 24304 27304 24312 27312
rect 24332 27304 24346 27312
rect 24348 27304 24350 27317
rect 24372 27312 24374 27317
rect 24396 27312 24398 27317
rect 24362 27304 24374 27312
rect 24390 27304 24402 27312
rect 24422 27304 24430 27312
rect 24312 27296 24320 27304
rect 24346 27296 24350 27304
rect 24360 27296 24362 27304
rect 24372 27296 24376 27304
rect 24388 27296 24390 27304
rect 24296 27088 24302 27096
rect 24278 27058 24281 27088
rect 24300 27066 24303 27088
rect 24323 27066 24326 27096
rect 24348 27067 24350 27296
rect 24372 27067 24374 27296
rect 24396 27067 24398 27304
rect 24402 27296 24404 27304
rect 24430 27296 24438 27304
rect 24286 27059 24294 27066
rect 24300 27059 24302 27066
rect 24303 27061 24308 27066
rect 24303 27059 24317 27061
rect 24286 27058 24317 27059
rect 24337 27058 24350 27067
rect 24357 27058 24377 27067
rect 24384 27058 24402 27067
rect 24286 27056 24287 27058
rect 24288 27056 24292 27058
rect 24300 27056 24302 27058
rect 24238 27037 24244 27038
rect 24250 27037 24254 27051
rect 24296 27040 24297 27056
rect 24248 27034 24254 27037
rect 24128 26996 24134 27010
rect 24226 27008 24240 27010
rect 24247 27008 24254 27034
rect 24298 27026 24302 27056
rect 24211 26996 24218 27002
rect 24226 26996 24230 27008
rect 24132 26987 24134 26996
rect 24221 26988 24230 26996
rect 24228 26987 24230 26988
rect 24252 26987 24254 27008
rect 24300 27004 24302 27026
rect 24287 26994 24290 26998
rect 24287 26988 24291 26994
rect 24296 26987 24302 27004
rect 24348 27055 24350 27058
rect 24348 27025 24357 27055
rect 24362 27048 24365 27055
rect 24372 27048 24374 27058
rect 24377 27048 24384 27058
rect 24372 27032 24388 27048
rect 24372 27025 24375 27032
rect 24348 26987 24350 27025
rect 24360 27002 24364 27012
rect 24372 27010 24374 27025
rect 24372 27002 24376 27010
rect 24358 26988 24366 26998
rect 24370 26996 24376 27002
rect 24377 26996 24384 27032
rect 24370 26988 24384 26996
rect 24368 26987 24377 26988
rect 24396 26987 24398 27058
rect 24425 27020 24428 27047
rect 24430 27025 24441 27047
rect 24443 27025 24446 27055
rect 24425 27017 24437 27020
rect 24468 26987 24470 27317
rect 24492 27312 24494 27317
rect 24516 27312 24518 27317
rect 24484 27304 24494 27312
rect 24512 27304 24522 27312
rect 24544 27304 24560 27312
rect 24478 27296 24484 27304
rect 24472 27049 24490 27059
rect 24492 27047 24494 27304
rect 24506 27296 24512 27304
rect 24516 27059 24518 27304
rect 24497 27049 24518 27059
rect 24526 27049 24532 27279
rect 24552 27096 24556 27106
rect 24564 27096 24566 27317
rect 24588 27312 24590 27317
rect 24612 27312 24614 27317
rect 24576 27304 24590 27312
rect 24604 27304 24616 27312
rect 24636 27304 24644 27312
rect 24572 27296 24576 27304
rect 24562 27082 24566 27096
rect 24538 27079 24542 27081
rect 24536 27071 24542 27079
rect 24548 27079 24566 27082
rect 24548 27071 24573 27079
rect 24537 27049 24542 27051
rect 24548 27049 24554 27071
rect 24562 27066 24573 27071
rect 24490 27017 24497 27047
rect 24504 27039 24508 27049
rect 24516 27047 24518 27049
rect 24516 27039 24522 27047
rect 24564 27041 24566 27066
rect 24512 27023 24522 27039
rect 24514 27017 24522 27023
rect 24561 27023 24568 27041
rect 24580 27031 24587 27066
rect 24588 27031 24590 27304
rect 24600 27296 24604 27304
rect 24593 27071 24600 27079
rect 24612 27071 24614 27304
rect 24644 27296 24652 27304
rect 24660 27096 24662 27317
rect 24664 27304 24672 27312
rect 24692 27304 24706 27312
rect 24708 27304 24710 27317
rect 24732 27312 24734 27317
rect 24756 27312 24758 27317
rect 24722 27304 24734 27312
rect 24750 27304 24762 27312
rect 24782 27304 24790 27312
rect 24810 27304 24826 27312
rect 24672 27296 24680 27304
rect 24706 27296 24710 27304
rect 24720 27296 24722 27304
rect 24732 27296 24736 27304
rect 24748 27296 24750 27304
rect 24656 27088 24662 27096
rect 24593 27066 24597 27071
rect 24607 27051 24614 27071
rect 24638 27058 24641 27088
rect 24660 27066 24663 27088
rect 24683 27066 24686 27096
rect 24708 27067 24710 27296
rect 24732 27067 24734 27296
rect 24756 27067 24758 27304
rect 24762 27296 24764 27304
rect 24790 27296 24798 27304
rect 24646 27059 24654 27066
rect 24660 27059 24662 27066
rect 24663 27061 24668 27066
rect 24663 27059 24677 27061
rect 24646 27058 24677 27059
rect 24697 27058 24710 27067
rect 24717 27058 24737 27067
rect 24744 27058 24762 27067
rect 24646 27056 24647 27058
rect 24648 27056 24652 27058
rect 24660 27056 24662 27058
rect 24607 27047 24618 27051
rect 24602 27041 24618 27047
rect 24593 27031 24597 27041
rect 24492 26991 24494 27017
rect 24514 27009 24518 27017
rect 24492 26987 24506 26991
rect 24516 26987 24518 27009
rect 24561 26987 24567 27023
rect 24580 27020 24583 27031
rect 24576 27010 24583 27020
rect 24588 27020 24597 27031
rect 24588 27015 24598 27020
rect 24580 26990 24583 27010
rect 24586 27010 24590 27015
rect 24593 27010 24598 27015
rect 24607 27015 24614 27041
rect 24656 27040 24657 27056
rect 24658 27026 24662 27056
rect 24586 27001 24600 27010
rect 24586 26996 24590 27001
rect 24593 26996 24598 27001
rect 24572 26987 24583 26990
rect 24588 26993 24590 26996
rect 24588 26987 24592 26993
rect 24607 26987 24610 27015
rect 24612 26987 24614 27015
rect 24660 27004 24662 27026
rect 24647 26994 24650 26998
rect 24647 26988 24651 26994
rect 24656 26987 24662 27004
rect 24708 27055 24710 27058
rect 24708 27025 24717 27055
rect 24722 27048 24725 27055
rect 24732 27048 24734 27058
rect 24737 27048 24744 27058
rect 24732 27032 24748 27048
rect 24732 27025 24735 27032
rect 24708 26987 24710 27025
rect 24720 27002 24724 27012
rect 24732 27010 24734 27025
rect 24732 27002 24736 27010
rect 24718 26988 24726 26998
rect 24730 26996 24736 27002
rect 24737 26996 24744 27032
rect 24730 26988 24744 26996
rect 24728 26987 24737 26988
rect 24756 26987 24758 27058
rect 24828 27055 24830 27317
rect 24852 27312 24854 27317
rect 24876 27312 24878 27317
rect 24842 27304 24854 27312
rect 24870 27304 24882 27312
rect 24902 27304 24910 27312
rect 24930 27304 24944 27312
rect 24838 27296 24842 27304
rect 24785 27020 24788 27047
rect 24790 27025 24801 27047
rect 24803 27025 24806 27055
rect 24828 27025 24837 27055
rect 24852 27025 24854 27304
rect 24866 27296 24870 27304
rect 24857 27025 24864 27055
rect 24876 27047 24878 27304
rect 24910 27296 24918 27304
rect 24944 27296 24946 27304
rect 24936 27096 24940 27106
rect 24948 27096 24950 27317
rect 24972 27312 24974 27317
rect 24996 27312 24998 27317
rect 24960 27304 24974 27312
rect 24988 27304 25000 27312
rect 25020 27304 25028 27312
rect 24958 27296 24960 27304
rect 24946 27066 24950 27096
rect 24785 27017 24797 27020
rect 24828 26987 24830 27025
rect 24847 27017 24854 27025
rect 24874 27017 24881 27047
rect 24905 27020 24908 27047
rect 24910 27025 24921 27047
rect 24923 27025 24926 27055
rect 24905 27017 24917 27020
rect 24840 27002 24844 27012
rect 24852 27002 24854 27017
rect 24857 27007 24864 27017
rect 24850 26988 24864 27002
rect 24874 26991 24878 27017
rect 24948 27004 24950 27066
rect 24964 27055 24971 27065
rect 24964 27047 24967 27055
rect 24964 27020 24971 27047
rect 24960 27017 24971 27020
rect 24960 27010 24967 27017
rect 24972 27010 24974 27304
rect 24986 27296 24988 27304
rect 24996 27104 24998 27304
rect 25000 27296 25002 27304
rect 25028 27296 25036 27304
rect 24991 27096 24998 27104
rect 25044 27096 25046 27317
rect 25048 27304 25056 27312
rect 25076 27304 25090 27312
rect 25092 27304 25094 27317
rect 25140 27312 25142 27317
rect 25260 27312 25262 27317
rect 25356 27312 25358 27317
rect 25380 27312 25382 27317
rect 25106 27304 25118 27312
rect 25134 27304 25146 27312
rect 25166 27304 25174 27312
rect 25194 27304 25210 27312
rect 25226 27304 25238 27312
rect 25254 27304 25266 27312
rect 25286 27304 25294 27312
rect 25314 27304 25330 27312
rect 25346 27304 25358 27312
rect 25374 27304 25386 27312
rect 25406 27304 25414 27312
rect 25056 27296 25064 27304
rect 25090 27296 25094 27304
rect 25104 27296 25106 27304
rect 25118 27296 25120 27304
rect 25132 27296 25134 27304
rect 24986 27095 25002 27096
rect 24977 27047 24981 27055
rect 24984 27051 24988 27061
rect 24991 27051 24994 27065
rect 24996 27051 24998 27095
rect 25040 27088 25046 27096
rect 25022 27058 25025 27088
rect 25044 27066 25047 27088
rect 25067 27066 25070 27096
rect 25030 27059 25038 27066
rect 25044 27059 25046 27066
rect 25047 27061 25052 27066
rect 25047 27059 25061 27061
rect 25030 27058 25061 27059
rect 25030 27056 25031 27058
rect 25032 27056 25036 27058
rect 25044 27056 25046 27058
rect 24991 27047 24998 27051
rect 24991 27021 25002 27047
rect 25040 27040 25041 27056
rect 25042 27026 25046 27056
rect 24991 27020 24998 27021
rect 24851 26987 24864 26988
rect 24876 26987 24878 26991
rect 24945 26987 24950 27004
rect 24964 26987 24967 27010
rect 24970 27007 24974 27010
rect 24977 27007 24982 27020
rect 24986 27017 24998 27020
rect 24970 26996 24984 27007
rect 24972 26987 24981 26996
rect 24991 26991 24998 27017
rect 25044 27004 25046 27026
rect 24991 26987 24994 26991
rect 24996 26987 24998 26991
rect 25031 26994 25034 26998
rect 25031 26988 25035 26994
rect 25040 26987 25046 27004
rect 25092 26987 25094 27296
rect 25130 27124 25131 27279
rect 25140 27124 25142 27304
rect 25146 27296 25148 27304
rect 25174 27296 25182 27304
rect 25222 27296 25226 27304
rect 25250 27296 25254 27304
rect 25145 27124 25146 27125
rect 25130 27118 25146 27124
rect 25130 27098 25131 27118
rect 25097 27082 25101 27096
rect 25121 27088 25123 27096
rect 25130 27090 25132 27098
rect 25128 27088 25132 27090
rect 25140 27088 25142 27118
rect 25238 27116 25254 27124
rect 25121 27082 25128 27088
rect 25130 27082 25146 27088
rect 25173 27082 25183 27104
rect 25217 27082 25224 27104
rect 25226 27082 25233 27112
rect 25238 27110 25243 27112
rect 25250 27110 25254 27112
rect 25235 27082 25241 27104
rect 25128 27058 25130 27082
rect 25120 27048 25124 27056
rect 25118 27036 25124 27048
rect 25116 27032 25124 27036
rect 25118 27022 25120 27032
rect 25118 27018 25132 27022
rect 25126 27010 25132 27018
rect 25140 27010 25142 27082
rect 25145 27058 25146 27082
rect 25243 27074 25250 27104
rect 25252 27082 25259 27104
rect 25210 27046 25218 27056
rect 25176 27038 25190 27046
rect 25220 27038 25234 27046
rect 25240 27038 25244 27056
rect 25220 27034 25228 27038
rect 25220 27032 25234 27034
rect 25238 27032 25244 27038
rect 25220 27028 25230 27032
rect 25226 27024 25230 27028
rect 25238 27024 25240 27032
rect 25136 26996 25142 27010
rect 25220 27002 25222 27014
rect 25236 27012 25240 27024
rect 25252 27020 25256 27024
rect 25246 27012 25256 27020
rect 25236 27008 25252 27012
rect 25260 27010 25262 27304
rect 25294 27296 25302 27304
rect 25342 27296 25346 27304
rect 25293 27082 25303 27104
rect 25296 27038 25310 27046
rect 25346 27025 25351 27055
rect 25356 27029 25358 27304
rect 25370 27296 25374 27304
rect 25380 27034 25382 27304
rect 25414 27296 25422 27304
rect 25356 27027 25377 27029
rect 25353 27025 25377 27027
rect 25356 27012 25358 27025
rect 25240 26996 25243 27008
rect 25256 26996 25262 27010
rect 25344 27002 25348 27012
rect 25356 27008 25372 27012
rect 25378 27008 25382 27034
rect 25409 27020 25412 27047
rect 25414 27025 25425 27047
rect 25427 27025 25430 27055
rect 25409 27017 25421 27020
rect 25356 27002 25358 27008
rect 25140 26987 25142 26996
rect 25260 26987 25262 26996
rect 25342 26988 25346 26998
rect 25354 26988 25358 27002
rect 25355 26987 25358 26988
rect 25380 26987 25382 27008
rect 25452 26987 25454 27317
rect 25476 27312 25478 27317
rect 25500 27312 25502 27317
rect 25468 27304 25478 27312
rect 25496 27304 25506 27312
rect 25528 27304 25544 27312
rect 25462 27296 25468 27304
rect 25456 27049 25474 27059
rect 25476 27047 25478 27304
rect 25490 27296 25496 27304
rect 25500 27059 25502 27304
rect 25481 27049 25502 27059
rect 25510 27049 25516 27279
rect 25536 27096 25540 27106
rect 25548 27096 25550 27317
rect 25572 27312 25574 27317
rect 25596 27312 25598 27317
rect 25560 27304 25574 27312
rect 25588 27304 25600 27312
rect 25620 27304 25628 27312
rect 25556 27296 25560 27304
rect 25546 27082 25550 27096
rect 25522 27079 25526 27081
rect 25520 27071 25526 27079
rect 25532 27079 25550 27082
rect 25532 27071 25557 27079
rect 25521 27049 25526 27051
rect 25532 27049 25538 27071
rect 25546 27066 25557 27071
rect 25474 27017 25481 27047
rect 25488 27039 25492 27049
rect 25500 27047 25502 27049
rect 25500 27039 25506 27047
rect 25548 27041 25550 27066
rect 25496 27023 25506 27039
rect 25498 27017 25506 27023
rect 25545 27023 25552 27041
rect 25564 27031 25571 27066
rect 25572 27031 25574 27304
rect 25584 27296 25588 27304
rect 25577 27071 25584 27079
rect 25596 27071 25598 27304
rect 25628 27296 25636 27304
rect 25644 27096 25646 27317
rect 26109 27314 26125 27317
rect 25648 27304 25656 27312
rect 25676 27304 25690 27312
rect 25707 27304 25719 27312
rect 25736 27304 25748 27312
rect 25767 27304 25777 27312
rect 25796 27304 25805 27312
rect 25825 27304 25833 27312
rect 25853 27304 25861 27312
rect 25881 27304 25890 27312
rect 25909 27304 25918 27312
rect 25938 27304 25946 27312
rect 25966 27304 25974 27312
rect 25994 27304 26002 27312
rect 26022 27304 26030 27312
rect 26050 27304 26058 27312
rect 26078 27304 26086 27312
rect 26272 27309 26274 27317
rect 26733 27314 26749 27317
rect 26134 27304 26142 27309
rect 26162 27304 26170 27309
rect 25656 27296 25664 27304
rect 25690 27296 25692 27304
rect 25704 27296 25707 27304
rect 25719 27296 25720 27304
rect 25732 27296 25736 27304
rect 25777 27296 25783 27304
rect 25805 27296 25812 27304
rect 25833 27296 25841 27304
rect 25861 27296 25869 27304
rect 25890 27296 25897 27304
rect 25918 27296 25925 27304
rect 25946 27296 25954 27304
rect 25974 27296 25982 27304
rect 26002 27296 26010 27304
rect 26030 27296 26038 27304
rect 26058 27296 26066 27304
rect 26086 27296 26094 27304
rect 26142 27293 26150 27304
rect 26170 27294 26178 27304
rect 26218 27301 26226 27309
rect 26246 27301 26254 27309
rect 26272 27301 26282 27309
rect 26302 27301 26314 27312
rect 26331 27301 26343 27312
rect 26360 27301 26372 27312
rect 26391 27304 26401 27312
rect 26420 27304 26429 27312
rect 26449 27304 26457 27312
rect 26477 27304 26485 27312
rect 26505 27304 26514 27312
rect 26533 27304 26542 27312
rect 26562 27304 26570 27312
rect 26590 27304 26598 27312
rect 26618 27304 26626 27312
rect 26646 27304 26654 27312
rect 26674 27304 26682 27312
rect 26702 27304 26710 27312
rect 26896 27309 26898 27317
rect 27060 27312 27062 27317
rect 27108 27312 27110 27317
rect 27180 27312 27182 27317
rect 27276 27312 27278 27317
rect 27324 27312 27326 27317
rect 26758 27304 26766 27309
rect 26786 27304 26794 27309
rect 26226 27294 26234 27301
rect 26254 27294 26262 27301
rect 26162 27293 26178 27294
rect 26218 27293 26234 27294
rect 26246 27293 26262 27294
rect 26272 27294 26274 27301
rect 26282 27294 26290 27301
rect 26314 27296 26318 27301
rect 26330 27296 26331 27301
rect 26343 27296 26346 27301
rect 26358 27296 26360 27301
rect 26372 27296 26374 27301
rect 26401 27296 26407 27304
rect 26429 27296 26436 27304
rect 26457 27296 26465 27304
rect 26485 27296 26493 27304
rect 26514 27296 26521 27304
rect 26542 27296 26549 27304
rect 26570 27296 26578 27304
rect 26598 27296 26606 27304
rect 26626 27296 26634 27304
rect 26654 27296 26662 27304
rect 26682 27296 26690 27304
rect 26710 27296 26718 27304
rect 26272 27293 26290 27294
rect 26302 27293 26310 27294
rect 26766 27293 26774 27304
rect 26794 27294 26802 27304
rect 26842 27301 26850 27309
rect 26870 27301 26878 27309
rect 26896 27301 26906 27309
rect 26926 27301 26942 27312
rect 26958 27301 26970 27312
rect 26986 27301 26998 27312
rect 27018 27304 27026 27312
rect 27046 27304 27062 27312
rect 27076 27304 27088 27312
rect 27104 27304 27116 27312
rect 27174 27304 27182 27312
rect 27202 27304 27208 27312
rect 27234 27304 27242 27312
rect 27262 27304 27278 27312
rect 27292 27304 27304 27312
rect 27320 27304 27332 27312
rect 27352 27304 27368 27312
rect 26850 27294 26858 27301
rect 26878 27294 26886 27301
rect 26786 27293 26802 27294
rect 26842 27293 26858 27294
rect 26870 27293 26886 27294
rect 26896 27294 26898 27301
rect 26906 27294 26914 27301
rect 26954 27296 26958 27301
rect 26982 27296 26986 27301
rect 27026 27296 27034 27304
rect 26896 27293 26914 27294
rect 26926 27293 26934 27294
rect 25822 27279 25955 27287
rect 25960 27279 26013 27287
rect 25970 27261 25974 27270
rect 26038 27269 26045 27278
rect 26021 27257 26027 27262
rect 26046 27257 26055 27269
rect 26017 27252 26021 27257
rect 26046 27253 26062 27257
rect 26063 27253 26066 27257
rect 25640 27088 25646 27096
rect 25577 27066 25581 27071
rect 25591 27051 25598 27071
rect 25622 27058 25625 27088
rect 25644 27066 25647 27088
rect 25667 27066 25670 27096
rect 25730 27088 25736 27248
rect 25795 27238 25801 27246
rect 25832 27238 25843 27242
rect 25805 27230 25811 27238
rect 25786 27210 25801 27230
rect 25832 27227 25845 27238
rect 25870 27230 25877 27238
rect 25861 27227 25877 27230
rect 25908 27227 25918 27249
rect 25786 27200 25805 27210
rect 25812 27200 25831 27210
rect 25805 27198 25811 27200
rect 25852 27198 25855 27227
rect 25861 27208 25869 27227
rect 25935 27219 25941 27249
rect 25976 27219 25981 27249
rect 26017 27227 26018 27252
rect 26050 27227 26057 27253
rect 25857 27200 25870 27208
rect 25805 27192 25812 27198
rect 25805 27190 25819 27192
rect 25805 27185 25828 27190
rect 25794 27160 25801 27170
rect 25812 27168 25828 27185
rect 25838 27168 25845 27198
rect 25859 27195 25877 27198
rect 25852 27166 25859 27190
rect 25867 27168 25877 27195
rect 26050 27193 26055 27227
rect 26087 27221 26096 27222
rect 26093 27219 26096 27221
rect 25928 27190 25934 27193
rect 25812 27160 25866 27166
rect 25867 27160 25876 27168
rect 25893 27163 25909 27190
rect 25928 27163 25931 27190
rect 25934 27163 25935 27190
rect 25969 27185 25974 27193
rect 25969 27163 25985 27185
rect 25991 27163 25999 27185
rect 25893 27160 25900 27163
rect 25935 27160 25941 27163
rect 25802 27153 25811 27160
rect 25969 27155 26007 27163
rect 26038 27155 26045 27185
rect 26050 27163 26057 27193
rect 26272 27186 26274 27293
rect 26446 27279 26579 27287
rect 26584 27279 26637 27287
rect 26594 27261 26598 27270
rect 26662 27269 26669 27278
rect 26645 27257 26651 27262
rect 26670 27257 26679 27269
rect 26641 27252 26645 27257
rect 26670 27253 26686 27257
rect 26687 27253 26690 27257
rect 26059 27163 26066 27185
rect 26071 27163 26075 27185
rect 26059 27155 26076 27163
rect 26160 27156 26172 27172
rect 25740 27118 25746 27130
rect 25728 27080 25736 27088
rect 25630 27059 25638 27066
rect 25644 27059 25646 27066
rect 25647 27061 25652 27066
rect 25647 27059 25661 27061
rect 25630 27058 25661 27059
rect 25728 27058 25733 27080
rect 25802 27070 25809 27153
rect 25852 27122 25855 27133
rect 25934 27132 25941 27148
rect 25943 27133 25973 27140
rect 26050 27130 26055 27155
rect 26251 27148 26252 27164
rect 26267 27162 26275 27186
rect 26066 27133 26080 27140
rect 25852 27092 25859 27122
rect 25969 27100 25974 27130
rect 26010 27100 26017 27130
rect 26038 27100 26039 27122
rect 26050 27100 26057 27130
rect 26023 27092 26045 27100
rect 26071 27092 26078 27122
rect 26129 27106 26142 27122
rect 26147 27106 26151 27136
rect 26229 27110 26245 27126
rect 26238 27101 26245 27110
rect 26250 27106 26252 27128
rect 26267 27106 26276 27146
rect 26353 27128 26360 27248
rect 26419 27238 26425 27246
rect 26456 27238 26467 27242
rect 26429 27230 26435 27238
rect 26410 27210 26425 27230
rect 26456 27227 26469 27238
rect 26494 27230 26501 27238
rect 26485 27227 26501 27230
rect 26532 27227 26542 27249
rect 26410 27200 26429 27210
rect 26436 27200 26455 27210
rect 26429 27198 26435 27200
rect 26476 27198 26479 27227
rect 26485 27208 26493 27227
rect 26559 27219 26565 27249
rect 26600 27219 26605 27249
rect 26641 27227 26642 27252
rect 26674 27227 26681 27253
rect 26481 27200 26494 27208
rect 26429 27192 26436 27198
rect 26429 27190 26443 27192
rect 26429 27185 26452 27190
rect 26418 27160 26425 27170
rect 26436 27168 26452 27185
rect 26462 27168 26469 27198
rect 26483 27195 26501 27198
rect 26476 27166 26483 27190
rect 26491 27168 26501 27195
rect 26674 27193 26679 27227
rect 26711 27221 26720 27222
rect 26717 27219 26720 27221
rect 26552 27190 26558 27193
rect 26436 27160 26490 27166
rect 26491 27160 26500 27168
rect 26517 27163 26533 27190
rect 26552 27163 26555 27190
rect 26558 27163 26559 27190
rect 26593 27185 26598 27193
rect 26593 27163 26609 27185
rect 26615 27163 26623 27185
rect 26517 27160 26524 27163
rect 26559 27160 26565 27163
rect 26426 27153 26435 27160
rect 26593 27155 26631 27163
rect 26662 27155 26669 27185
rect 26674 27163 26681 27193
rect 26896 27186 26898 27293
rect 26683 27163 26690 27185
rect 26695 27163 26699 27185
rect 26683 27155 26700 27163
rect 26784 27156 26796 27172
rect 26221 27098 26225 27101
rect 26236 27098 26252 27101
rect 26351 27098 26360 27128
rect 26364 27100 26369 27128
rect 25852 27070 25855 27092
rect 26050 27083 26055 27092
rect 25786 27062 25838 27070
rect 25845 27062 25857 27070
rect 25901 27062 25937 27070
rect 25630 27056 25631 27058
rect 25632 27056 25636 27058
rect 25644 27056 25646 27058
rect 25591 27047 25602 27051
rect 25586 27041 25602 27047
rect 25577 27031 25581 27041
rect 25476 26991 25478 27017
rect 25498 27009 25502 27017
rect 25476 26987 25490 26991
rect 25500 26987 25502 27009
rect 25545 26987 25551 27023
rect 25564 27020 25567 27031
rect 25560 27010 25567 27020
rect 25572 27020 25581 27031
rect 25572 27015 25582 27020
rect 25564 26990 25567 27010
rect 25570 27010 25574 27015
rect 25577 27010 25582 27015
rect 25591 27015 25598 27041
rect 25640 27040 25641 27056
rect 25642 27026 25646 27056
rect 25570 27001 25584 27010
rect 25570 26996 25574 27001
rect 25577 26996 25582 27001
rect 25556 26987 25567 26990
rect 25572 26993 25574 26996
rect 25572 26987 25576 26993
rect 25591 26987 25594 27015
rect 25596 26987 25598 27015
rect 25644 27004 25646 27026
rect 25631 26994 25634 26998
rect 25631 26988 25635 26994
rect 25640 26987 25646 27004
rect 25802 26987 25809 27062
rect 25852 27060 25855 27062
rect 25838 27052 25845 27060
rect 25838 27030 25854 27052
rect 25870 27030 25877 27060
rect 25928 27052 25934 27060
rect 25969 27052 25974 27060
rect 26050 27057 26057 27083
rect 26050 27052 26055 27057
rect 25911 27030 25923 27052
rect 25928 27030 25929 27052
rect 25934 27030 25935 27052
rect 25974 27030 25976 27052
rect 25987 27030 26002 27052
rect 25935 27027 25941 27030
rect 25907 27022 25941 27027
rect 25976 27022 25981 27030
rect 26038 27022 26045 27052
rect 26071 27026 26078 27052
rect 26080 27047 26088 27082
rect 26159 27027 26163 27043
rect 26164 27041 26175 27043
rect 26211 27041 26217 27098
rect 26230 27071 26231 27073
rect 26238 27071 26244 27098
rect 26287 27083 26290 27091
rect 26297 27081 26300 27083
rect 26227 27041 26234 27071
rect 26240 27041 26245 27063
rect 26250 27041 26256 27063
rect 26258 27041 26265 27071
rect 26267 27041 26276 27081
rect 26277 27041 26283 27063
rect 26285 27041 26292 27071
rect 26297 27041 26303 27081
rect 26334 27070 26356 27073
rect 26366 27070 26379 27073
rect 26426 27070 26433 27153
rect 26476 27122 26479 27133
rect 26558 27132 26565 27148
rect 26567 27133 26597 27140
rect 26674 27130 26679 27155
rect 26875 27148 26876 27164
rect 26891 27162 26899 27186
rect 26690 27133 26704 27140
rect 26476 27092 26483 27122
rect 26593 27100 26598 27130
rect 26634 27100 26641 27130
rect 26662 27100 26663 27122
rect 26674 27100 26681 27130
rect 26647 27092 26669 27100
rect 26695 27092 26702 27122
rect 26753 27106 26766 27122
rect 26771 27106 26775 27136
rect 26853 27110 26869 27126
rect 26862 27101 26869 27110
rect 26874 27106 26876 27128
rect 26891 27106 26900 27146
rect 26983 27107 26993 27119
rect 26845 27098 26849 27101
rect 26860 27098 26876 27101
rect 26989 27098 26993 27107
rect 26995 27107 27003 27279
rect 26995 27098 27005 27107
rect 26476 27070 26479 27092
rect 26674 27083 26679 27092
rect 26174 27035 26175 27041
rect 26238 27033 26245 27041
rect 26267 27033 26275 27041
rect 26351 27033 26357 27063
rect 26410 27062 26462 27070
rect 26469 27062 26481 27070
rect 26525 27062 26561 27070
rect 26062 27022 26078 27026
rect 25852 26987 25855 27022
rect 25923 26999 25927 27015
rect 25928 26987 25931 26995
rect 25987 26991 26003 26993
rect 26050 26987 26055 27022
rect 26238 27018 26244 27033
rect 26137 27008 26145 27018
rect 26238 27013 26253 27018
rect 26147 27008 26156 27011
rect 26147 26992 26155 27008
rect 26156 26995 26163 27008
rect 26238 27003 26244 27013
rect 26268 26987 26275 27033
rect 26426 26987 26433 27062
rect 26476 27060 26479 27062
rect 26462 27052 26469 27060
rect 26462 27030 26478 27052
rect 26494 27030 26501 27060
rect 26552 27052 26558 27060
rect 26593 27052 26598 27060
rect 26674 27057 26681 27083
rect 26674 27052 26679 27057
rect 26535 27030 26547 27052
rect 26552 27030 26553 27052
rect 26558 27030 26559 27052
rect 26598 27030 26600 27052
rect 26611 27030 26626 27052
rect 26559 27027 26565 27030
rect 26531 27022 26565 27027
rect 26600 27022 26605 27030
rect 26662 27022 26669 27052
rect 26695 27026 26702 27052
rect 26704 27047 26712 27082
rect 26783 27027 26787 27043
rect 26788 27041 26799 27043
rect 26835 27041 26841 27098
rect 26854 27071 26855 27073
rect 26862 27071 26868 27098
rect 26911 27083 26914 27091
rect 26921 27081 26924 27083
rect 26851 27041 26858 27071
rect 26864 27041 26869 27063
rect 26874 27041 26880 27063
rect 26882 27041 26889 27071
rect 26891 27041 26900 27081
rect 26901 27041 26907 27063
rect 26909 27041 26916 27071
rect 26921 27041 26927 27081
rect 26968 27073 26975 27078
rect 26995 27073 27000 27093
rect 26798 27035 26799 27041
rect 26862 27033 26869 27041
rect 26891 27033 26899 27041
rect 26686 27022 26702 27026
rect 26476 26987 26479 27022
rect 26547 26999 26551 27015
rect 26552 26987 26555 26995
rect 26611 26991 26627 26993
rect 26674 26987 26679 27022
rect 26862 27018 26868 27033
rect 26761 27008 26769 27018
rect 26862 27013 26877 27018
rect 26771 27008 26780 27011
rect 26771 26992 26779 27008
rect 26780 26995 26787 27008
rect 26862 27003 26868 27013
rect 26892 26987 26899 27033
rect 26968 27033 26976 27073
rect 26984 27063 26993 27064
rect 26977 27048 26984 27063
rect 26986 27033 26993 27063
rect 26995 27048 27003 27073
rect 27060 27059 27062 27304
rect 27074 27296 27076 27304
rect 27088 27296 27090 27304
rect 27102 27296 27104 27304
rect 27071 27083 27087 27091
rect 27053 27049 27062 27059
rect 27064 27049 27070 27079
rect 27071 27077 27082 27079
rect 27071 27049 27080 27070
rect 26954 27013 26963 27023
rect 26968 27013 26973 27033
rect 26964 26999 26973 27013
rect 26968 26990 26973 26999
rect 27060 27015 27062 27049
rect 27063 27040 27070 27049
rect 27082 27040 27087 27070
rect 27063 27015 27064 27040
rect 27096 27039 27100 27049
rect 27108 27039 27110 27304
rect 27116 27296 27118 27304
rect 27164 27296 27174 27304
rect 27130 27079 27134 27081
rect 27128 27071 27134 27079
rect 27129 27049 27134 27051
rect 27140 27049 27146 27071
rect 27060 26991 27064 27015
rect 27070 27004 27072 27014
rect 27082 27004 27089 27015
rect 27106 27009 27110 27039
rect 27060 26987 27062 26991
rect 27063 26987 27064 26991
rect 27080 26991 27089 27004
rect 27094 26991 27098 27004
rect 27080 26990 27094 26991
rect 27082 26989 27090 26990
rect 27108 26987 27110 27009
rect 27180 27013 27182 27304
rect 27192 27296 27202 27304
rect 27242 27296 27250 27304
rect 27185 27048 27192 27078
rect 27194 27048 27200 27071
rect 27202 27041 27209 27071
rect 27211 27048 27220 27279
rect 27276 27059 27278 27304
rect 27290 27296 27292 27304
rect 27304 27296 27306 27304
rect 27318 27296 27320 27304
rect 27287 27083 27303 27091
rect 27269 27049 27278 27059
rect 27280 27049 27286 27079
rect 27287 27077 27298 27079
rect 27287 27049 27296 27070
rect 27194 27013 27196 27023
rect 27202 27015 27206 27041
rect 27276 27015 27278 27049
rect 27279 27040 27286 27049
rect 27298 27040 27303 27070
rect 27279 27015 27280 27040
rect 27312 27039 27316 27049
rect 27324 27039 27326 27304
rect 27332 27296 27334 27304
rect 27360 27096 27364 27106
rect 27372 27096 27374 27317
rect 27396 27312 27398 27317
rect 27420 27312 27422 27317
rect 27384 27304 27398 27312
rect 27412 27304 27424 27312
rect 27444 27304 27452 27312
rect 27380 27296 27384 27304
rect 27370 27082 27374 27096
rect 27346 27079 27350 27081
rect 27344 27071 27350 27079
rect 27356 27079 27374 27082
rect 27356 27071 27381 27079
rect 27345 27049 27350 27051
rect 27356 27049 27362 27071
rect 27370 27066 27381 27071
rect 27372 27041 27374 27066
rect 27180 27001 27194 27013
rect 27204 27001 27206 27013
rect 27180 26993 27182 27001
rect 27180 26987 27184 26993
rect 27276 26991 27280 27015
rect 27286 27004 27288 27014
rect 27298 27004 27305 27015
rect 27322 27009 27326 27039
rect 27276 26987 27278 26991
rect 27279 26987 27280 26991
rect 27296 26991 27305 27004
rect 27310 26991 27314 27004
rect 27296 26990 27310 26991
rect 27298 26989 27306 26990
rect 27324 26987 27326 27009
rect 27369 27023 27376 27041
rect 27388 27031 27395 27066
rect 27396 27031 27398 27304
rect 27408 27296 27412 27304
rect 27401 27071 27408 27079
rect 27420 27071 27422 27304
rect 27452 27296 27460 27304
rect 27468 27096 27470 27317
rect 27516 27312 27518 27317
rect 27540 27312 27542 27317
rect 27564 27312 27566 27317
rect 28029 27314 28045 27317
rect 28749 27314 28765 27317
rect 29469 27314 29485 27317
rect 30189 27314 30205 27317
rect 27472 27304 27480 27312
rect 27500 27304 27518 27312
rect 27532 27304 27544 27312
rect 27560 27304 27572 27312
rect 27627 27304 27636 27312
rect 27656 27304 27664 27312
rect 27687 27304 27697 27312
rect 27716 27304 27725 27312
rect 27745 27304 27753 27312
rect 27773 27304 27781 27312
rect 27801 27304 27810 27312
rect 27829 27304 27838 27312
rect 27858 27304 27866 27312
rect 27886 27304 27894 27312
rect 27914 27304 27922 27312
rect 27942 27304 27950 27312
rect 27970 27304 27978 27312
rect 27998 27304 28006 27312
rect 28062 27304 28070 27308
rect 28090 27304 28098 27308
rect 27480 27296 27488 27304
rect 27464 27088 27470 27096
rect 27401 27066 27405 27071
rect 27415 27051 27422 27071
rect 27446 27058 27449 27088
rect 27468 27066 27471 27088
rect 27491 27066 27494 27096
rect 27454 27059 27462 27066
rect 27468 27059 27470 27066
rect 27471 27061 27476 27066
rect 27471 27059 27485 27061
rect 27454 27058 27485 27059
rect 27454 27056 27455 27058
rect 27456 27056 27460 27058
rect 27468 27056 27470 27058
rect 27415 27047 27426 27051
rect 27410 27041 27426 27047
rect 27401 27031 27405 27041
rect 27369 26987 27375 27023
rect 27388 27020 27391 27031
rect 27384 27010 27391 27020
rect 27396 27020 27405 27031
rect 27396 27015 27406 27020
rect 27388 26990 27391 27010
rect 27394 27010 27398 27015
rect 27401 27010 27406 27015
rect 27415 27015 27422 27041
rect 27464 27040 27465 27056
rect 27466 27026 27470 27056
rect 27394 27001 27408 27010
rect 27394 26996 27398 27001
rect 27401 26996 27406 27001
rect 27380 26987 27391 26990
rect 27396 26993 27398 26996
rect 27396 26987 27400 26993
rect 27415 26987 27418 27015
rect 27420 26987 27422 27015
rect 27468 27004 27470 27026
rect 27455 26994 27458 26998
rect 27455 26988 27459 26994
rect 27464 26987 27470 27004
rect 27516 26987 27518 27304
rect 27528 27296 27532 27304
rect 27540 27087 27542 27304
rect 27556 27296 27560 27304
rect 27564 27087 27566 27304
rect 27620 27296 27627 27304
rect 27648 27296 27656 27304
rect 27697 27296 27703 27304
rect 27725 27296 27732 27304
rect 27753 27296 27761 27304
rect 27781 27296 27789 27304
rect 27810 27296 27817 27304
rect 27838 27296 27845 27304
rect 27866 27296 27874 27304
rect 27894 27296 27902 27304
rect 27922 27296 27930 27304
rect 27950 27296 27958 27304
rect 27978 27296 27986 27304
rect 28006 27296 28014 27304
rect 28054 27294 28062 27304
rect 28082 27294 28090 27304
rect 28122 27301 28130 27308
rect 28150 27301 28158 27308
rect 28178 27301 28186 27308
rect 28206 27301 28214 27308
rect 28234 27301 28242 27308
rect 28262 27301 28270 27308
rect 28290 27301 28298 27308
rect 28318 27301 28330 27312
rect 28347 27301 28359 27312
rect 28376 27301 28388 27312
rect 28407 27304 28417 27312
rect 28436 27304 28445 27312
rect 28465 27304 28473 27312
rect 28493 27304 28501 27312
rect 28521 27304 28530 27312
rect 28549 27304 28558 27312
rect 28578 27304 28586 27312
rect 28606 27304 28614 27312
rect 28634 27304 28642 27312
rect 28662 27304 28670 27312
rect 28690 27304 28698 27312
rect 28718 27304 28726 27312
rect 28782 27304 28790 27308
rect 28810 27304 28818 27308
rect 28130 27294 28138 27301
rect 28158 27294 28166 27301
rect 28186 27294 28194 27301
rect 28214 27294 28222 27301
rect 28242 27294 28250 27301
rect 28270 27294 28278 27301
rect 28298 27294 28306 27301
rect 28330 27296 28334 27301
rect 28346 27296 28347 27301
rect 28359 27296 28362 27301
rect 28374 27296 28376 27301
rect 28388 27296 28390 27301
rect 28417 27296 28423 27304
rect 28445 27296 28452 27304
rect 28473 27296 28481 27304
rect 28501 27296 28509 27304
rect 28530 27296 28537 27304
rect 28558 27296 28565 27304
rect 28586 27296 28594 27304
rect 28614 27296 28622 27304
rect 28642 27296 28650 27304
rect 28670 27296 28678 27304
rect 28698 27296 28706 27304
rect 28726 27296 28734 27304
rect 28774 27294 28782 27304
rect 28802 27294 28810 27304
rect 28842 27301 28850 27308
rect 28870 27301 28878 27308
rect 28898 27301 28906 27308
rect 28926 27301 28934 27308
rect 28954 27301 28962 27308
rect 28982 27301 28990 27308
rect 29010 27301 29018 27308
rect 29038 27301 29050 27312
rect 29067 27301 29079 27312
rect 29096 27301 29108 27312
rect 29127 27304 29137 27312
rect 29156 27304 29165 27312
rect 29185 27304 29193 27312
rect 29213 27304 29221 27312
rect 29241 27304 29250 27312
rect 29269 27304 29278 27312
rect 29298 27304 29306 27312
rect 29326 27304 29334 27312
rect 29354 27304 29362 27312
rect 29382 27304 29390 27312
rect 29410 27304 29418 27312
rect 29438 27304 29446 27312
rect 29502 27304 29510 27308
rect 29530 27304 29538 27308
rect 28850 27294 28858 27301
rect 28878 27294 28886 27301
rect 28906 27294 28914 27301
rect 28934 27294 28942 27301
rect 28962 27294 28970 27301
rect 28990 27294 28998 27301
rect 29018 27294 29026 27301
rect 29050 27296 29054 27301
rect 29066 27296 29067 27301
rect 29079 27296 29082 27301
rect 29094 27296 29096 27301
rect 29108 27296 29110 27301
rect 29137 27296 29143 27304
rect 29165 27296 29172 27304
rect 29193 27296 29201 27304
rect 29221 27296 29229 27304
rect 29250 27296 29257 27304
rect 29278 27296 29285 27304
rect 29306 27296 29314 27304
rect 29334 27296 29342 27304
rect 29362 27296 29370 27304
rect 29390 27296 29398 27304
rect 29418 27296 29426 27304
rect 29446 27296 29454 27304
rect 29494 27294 29502 27304
rect 29522 27294 29530 27304
rect 29562 27301 29570 27308
rect 29590 27301 29598 27308
rect 29618 27301 29626 27308
rect 29646 27301 29654 27308
rect 29674 27301 29682 27308
rect 29702 27301 29710 27308
rect 29730 27301 29738 27308
rect 29758 27301 29770 27312
rect 29787 27301 29799 27312
rect 29816 27301 29828 27312
rect 29847 27304 29857 27312
rect 29876 27304 29885 27312
rect 29905 27304 29913 27312
rect 29933 27304 29941 27312
rect 29961 27304 29970 27312
rect 29989 27304 29998 27312
rect 30018 27304 30026 27312
rect 30046 27304 30054 27312
rect 30074 27304 30082 27312
rect 30102 27304 30110 27312
rect 30130 27304 30138 27312
rect 30158 27304 30166 27312
rect 30222 27304 30230 27308
rect 30250 27304 30258 27308
rect 29570 27294 29578 27301
rect 29598 27294 29606 27301
rect 29626 27294 29634 27301
rect 29654 27294 29662 27301
rect 29682 27294 29690 27301
rect 29710 27294 29718 27301
rect 29738 27294 29746 27301
rect 29770 27296 29774 27301
rect 29786 27296 29787 27301
rect 29799 27296 29802 27301
rect 29814 27296 29816 27301
rect 29828 27296 29830 27301
rect 29857 27296 29863 27304
rect 29885 27296 29892 27304
rect 29913 27296 29921 27304
rect 29941 27296 29949 27304
rect 29970 27296 29977 27304
rect 29998 27296 30005 27304
rect 30026 27296 30034 27304
rect 30054 27296 30062 27304
rect 30082 27296 30090 27304
rect 30110 27296 30118 27304
rect 30138 27296 30146 27304
rect 30166 27296 30174 27304
rect 30214 27294 30222 27304
rect 30242 27294 30250 27304
rect 30282 27301 30290 27308
rect 30310 27301 30318 27308
rect 30338 27301 30346 27308
rect 30366 27301 30374 27308
rect 30394 27301 30402 27308
rect 30422 27301 30430 27308
rect 30450 27301 30458 27308
rect 30478 27301 30490 27312
rect 30492 27301 30494 27317
rect 30540 27312 30542 27317
rect 30506 27301 30518 27312
rect 30534 27301 30546 27312
rect 30566 27304 30574 27312
rect 30594 27304 30608 27312
rect 30290 27294 30298 27301
rect 30318 27294 30326 27301
rect 30346 27294 30354 27301
rect 30374 27294 30382 27301
rect 30402 27294 30410 27301
rect 30430 27294 30438 27301
rect 30458 27294 30466 27301
rect 30490 27296 30494 27301
rect 30518 27296 30522 27301
rect 28046 27292 28062 27294
rect 28074 27292 28090 27294
rect 28102 27292 28110 27294
rect 28122 27292 28138 27294
rect 28150 27292 28166 27294
rect 28178 27292 28194 27294
rect 28206 27292 28222 27294
rect 28234 27292 28250 27294
rect 28262 27292 28278 27294
rect 28290 27292 28306 27294
rect 28318 27292 28326 27294
rect 28766 27292 28782 27294
rect 28794 27292 28810 27294
rect 28822 27292 28830 27294
rect 28842 27292 28858 27294
rect 28870 27292 28886 27294
rect 28898 27292 28914 27294
rect 28926 27292 28942 27294
rect 28954 27292 28970 27294
rect 28982 27292 28998 27294
rect 29010 27292 29026 27294
rect 29038 27292 29046 27294
rect 29486 27292 29502 27294
rect 29514 27292 29530 27294
rect 29542 27292 29550 27294
rect 29562 27292 29578 27294
rect 29590 27292 29606 27294
rect 29618 27292 29634 27294
rect 29646 27292 29662 27294
rect 29674 27292 29690 27294
rect 29702 27292 29718 27294
rect 29730 27292 29746 27294
rect 29758 27292 29766 27294
rect 30206 27292 30222 27294
rect 30234 27292 30250 27294
rect 30262 27292 30270 27294
rect 30282 27292 30298 27294
rect 30310 27292 30326 27294
rect 30338 27292 30354 27294
rect 30366 27292 30382 27294
rect 30394 27292 30410 27294
rect 30422 27292 30438 27294
rect 30450 27292 30466 27294
rect 30478 27292 30486 27294
rect 27742 27279 27875 27287
rect 27880 27279 27933 27287
rect 28462 27279 28595 27287
rect 28600 27279 28653 27287
rect 29182 27279 29315 27287
rect 29320 27279 29373 27287
rect 29902 27279 30035 27287
rect 30040 27279 30093 27287
rect 27574 27146 27580 27279
rect 27890 27261 27894 27270
rect 27958 27269 27965 27278
rect 27941 27257 27947 27262
rect 27966 27257 27975 27269
rect 28610 27261 28614 27270
rect 28678 27269 28685 27278
rect 28661 27257 28667 27262
rect 28686 27257 28695 27269
rect 29330 27261 29334 27270
rect 29398 27269 29405 27278
rect 29381 27257 29387 27262
rect 29406 27257 29415 27269
rect 30050 27261 30054 27270
rect 30118 27269 30125 27278
rect 30101 27257 30107 27262
rect 30126 27257 30135 27269
rect 27937 27252 27941 27257
rect 27966 27253 27982 27257
rect 27983 27253 27986 27257
rect 27574 27133 27582 27146
rect 27538 27079 27545 27087
rect 27520 27049 27525 27079
rect 27530 27049 27536 27058
rect 27540 27051 27542 27079
rect 27564 27058 27570 27087
rect 27574 27058 27580 27133
rect 27586 27079 27590 27081
rect 27650 27080 27656 27248
rect 27715 27238 27721 27246
rect 27752 27238 27763 27242
rect 27725 27230 27731 27238
rect 27706 27210 27721 27230
rect 27752 27227 27765 27238
rect 27790 27230 27797 27238
rect 27781 27227 27797 27230
rect 27828 27227 27838 27249
rect 27706 27200 27725 27210
rect 27732 27200 27751 27210
rect 27725 27198 27731 27200
rect 27772 27198 27775 27227
rect 27781 27208 27789 27227
rect 27855 27219 27861 27249
rect 27896 27219 27901 27249
rect 27937 27227 27938 27252
rect 27970 27227 27977 27253
rect 28657 27252 28661 27257
rect 28686 27253 28702 27257
rect 28703 27253 28706 27257
rect 28435 27238 28441 27246
rect 28472 27238 28483 27242
rect 28445 27230 28451 27238
rect 27777 27200 27790 27208
rect 27725 27192 27732 27198
rect 27725 27190 27739 27192
rect 27725 27185 27748 27190
rect 27714 27160 27721 27170
rect 27732 27168 27748 27185
rect 27758 27168 27765 27198
rect 27779 27195 27797 27198
rect 27772 27166 27779 27190
rect 27787 27168 27797 27195
rect 27970 27193 27975 27227
rect 28007 27221 28016 27222
rect 28013 27219 28016 27221
rect 28426 27210 28441 27230
rect 28472 27227 28485 27238
rect 28510 27230 28517 27238
rect 28501 27227 28517 27230
rect 28548 27227 28558 27249
rect 28426 27200 28445 27210
rect 28452 27200 28471 27210
rect 28445 27198 28451 27200
rect 28492 27198 28495 27227
rect 28501 27208 28509 27227
rect 28575 27219 28581 27249
rect 28616 27219 28621 27249
rect 28657 27227 28658 27252
rect 28690 27227 28697 27253
rect 29377 27252 29381 27257
rect 29406 27253 29422 27257
rect 29423 27253 29426 27257
rect 29155 27238 29161 27246
rect 29192 27238 29203 27242
rect 29165 27230 29171 27238
rect 28497 27200 28510 27208
rect 28266 27195 28267 27196
rect 28280 27195 28282 27196
rect 27848 27190 27854 27193
rect 27732 27160 27786 27166
rect 27787 27160 27796 27168
rect 27813 27163 27829 27190
rect 27848 27163 27851 27190
rect 27854 27163 27855 27190
rect 27889 27185 27894 27193
rect 27889 27163 27905 27185
rect 27911 27163 27919 27185
rect 27813 27160 27820 27163
rect 27855 27160 27861 27163
rect 27722 27153 27731 27160
rect 27889 27155 27927 27163
rect 27958 27155 27965 27185
rect 27970 27163 27977 27193
rect 27979 27163 27986 27185
rect 27991 27163 27995 27185
rect 27979 27155 27996 27163
rect 28079 27155 28092 27183
rect 28145 27175 28149 27183
rect 28158 27175 28159 27193
rect 28227 27185 28246 27193
rect 28266 27188 28282 27195
rect 28170 27183 28178 27185
rect 28199 27183 28206 27185
rect 28170 27175 28180 27183
rect 28199 27175 28207 27183
rect 28225 27175 28227 27177
rect 28232 27175 28234 27183
rect 28262 27175 28264 27183
rect 28266 27182 28282 27183
rect 28301 27175 28310 27183
rect 28360 27175 28366 27185
rect 28376 27175 28378 27193
rect 28445 27192 28452 27198
rect 28445 27190 28459 27192
rect 28445 27185 28468 27190
rect 27660 27125 27666 27130
rect 27584 27071 27590 27079
rect 27545 27053 27552 27058
rect 27545 27051 27561 27053
rect 27537 27049 27561 27051
rect 27540 27010 27542 27049
rect 27550 27039 27556 27049
rect 27564 27039 27566 27058
rect 27585 27049 27590 27051
rect 27596 27049 27602 27071
rect 27648 27041 27653 27071
rect 27722 27070 27729 27153
rect 27772 27122 27775 27133
rect 27854 27132 27861 27148
rect 27863 27133 27893 27140
rect 27970 27130 27975 27155
rect 28155 27153 28159 27175
rect 27986 27133 28000 27140
rect 27772 27092 27779 27122
rect 27889 27100 27894 27130
rect 27930 27100 27937 27130
rect 27958 27100 27959 27122
rect 27970 27100 27977 27130
rect 28059 27129 28062 27139
rect 28069 27122 28072 27129
rect 28136 27123 28145 27153
rect 28155 27145 28158 27153
rect 27943 27092 27965 27100
rect 27991 27092 27998 27122
rect 28181 27113 28188 27175
rect 28200 27153 28206 27175
rect 28225 27153 28232 27175
rect 28257 27153 28262 27175
rect 28301 27153 28308 27175
rect 28313 27153 28320 27175
rect 28370 27168 28386 27175
rect 28368 27161 28383 27168
rect 28209 27145 28212 27153
rect 28222 27145 28227 27153
rect 28255 27145 28257 27153
rect 28285 27145 28292 27153
rect 28313 27145 28317 27153
rect 28368 27145 28376 27161
rect 28434 27160 28441 27170
rect 28452 27168 28468 27185
rect 28478 27168 28485 27198
rect 28499 27195 28517 27198
rect 28492 27166 28499 27190
rect 28507 27168 28517 27195
rect 28690 27193 28695 27227
rect 28727 27221 28736 27222
rect 28733 27219 28736 27221
rect 29146 27210 29161 27230
rect 29192 27227 29205 27238
rect 29230 27230 29237 27238
rect 29221 27227 29237 27230
rect 29268 27227 29278 27249
rect 29146 27200 29165 27210
rect 29172 27200 29191 27210
rect 29165 27198 29171 27200
rect 29212 27198 29215 27227
rect 29221 27208 29229 27227
rect 29295 27219 29301 27249
rect 29336 27219 29341 27249
rect 29377 27227 29378 27252
rect 29410 27227 29417 27253
rect 30097 27252 30101 27257
rect 30126 27253 30142 27257
rect 30143 27253 30146 27257
rect 29875 27238 29881 27246
rect 29912 27238 29923 27242
rect 29885 27230 29891 27238
rect 29217 27200 29230 27208
rect 28986 27195 28987 27196
rect 29000 27195 29002 27196
rect 28568 27190 28574 27193
rect 28452 27160 28506 27166
rect 28507 27160 28516 27168
rect 28533 27163 28549 27190
rect 28568 27163 28571 27190
rect 28574 27163 28575 27190
rect 28609 27185 28614 27193
rect 28609 27163 28625 27185
rect 28631 27163 28639 27185
rect 28533 27160 28540 27163
rect 28575 27160 28581 27163
rect 28246 27125 28297 27133
rect 28145 27105 28284 27113
rect 27772 27070 27775 27092
rect 27970 27083 27975 27092
rect 27706 27062 27758 27070
rect 27765 27062 27777 27070
rect 27821 27062 27857 27070
rect 27560 27023 27566 27039
rect 27530 26991 27534 27000
rect 27540 26996 27544 27010
rect 27562 27009 27566 27023
rect 27538 26987 27545 26996
rect 27564 26987 27566 27009
rect 27722 26987 27729 27062
rect 27772 27060 27775 27062
rect 27758 27052 27765 27060
rect 27758 27030 27774 27052
rect 27790 27030 27797 27060
rect 27848 27052 27854 27060
rect 27889 27052 27894 27060
rect 27970 27057 27977 27083
rect 27970 27052 27975 27057
rect 27831 27030 27843 27052
rect 27848 27030 27849 27052
rect 27854 27030 27855 27052
rect 27894 27030 27896 27052
rect 27907 27030 27922 27052
rect 27855 27022 27861 27030
rect 27896 27022 27901 27030
rect 27958 27022 27965 27052
rect 27991 27026 27998 27052
rect 28000 27047 28008 27082
rect 28039 27060 28045 27070
rect 28049 27049 28055 27060
rect 28125 27049 28131 27052
rect 28049 27044 28050 27049
rect 28079 27030 28095 27043
rect 28079 27027 28082 27030
rect 28092 27027 28095 27030
rect 28125 27033 28140 27049
rect 27982 27022 27998 27026
rect 27772 26987 27775 27022
rect 27848 26987 27851 26995
rect 27970 26987 27975 27022
rect 28049 27013 28054 27027
rect 28125 27022 28131 27033
rect 28135 27022 28141 27031
rect 28151 27023 28158 27105
rect 28181 27093 28188 27105
rect 28180 27085 28200 27093
rect 28227 27085 28239 27093
rect 28249 27085 28263 27093
rect 28274 27085 28290 27093
rect 28181 27083 28188 27085
rect 28264 27083 28265 27085
rect 28173 27064 28180 27083
rect 28163 27053 28180 27064
rect 28200 27079 28206 27083
rect 28200 27069 28207 27079
rect 28237 27075 28239 27083
rect 28255 27075 28257 27077
rect 28262 27075 28265 27083
rect 28200 27053 28206 27069
rect 28211 27053 28217 27069
rect 28237 27053 28253 27075
rect 28255 27053 28262 27075
rect 28264 27053 28282 27075
rect 28301 27061 28302 27145
rect 28316 27135 28317 27145
rect 28373 27115 28376 27145
rect 28442 27153 28451 27160
rect 28609 27155 28647 27163
rect 28678 27155 28685 27185
rect 28690 27163 28697 27193
rect 28699 27163 28706 27185
rect 28711 27163 28715 27185
rect 28699 27155 28716 27163
rect 28799 27155 28812 27183
rect 28865 27175 28869 27183
rect 28878 27175 28879 27193
rect 28947 27185 28966 27193
rect 28986 27188 29002 27195
rect 28890 27183 28898 27185
rect 28919 27183 28926 27185
rect 28890 27175 28900 27183
rect 28919 27175 28927 27183
rect 28945 27175 28947 27177
rect 28952 27175 28954 27183
rect 28982 27175 28984 27183
rect 28986 27182 29002 27183
rect 29021 27175 29030 27183
rect 29080 27175 29086 27185
rect 29096 27175 29098 27193
rect 29165 27192 29172 27198
rect 29165 27190 29179 27192
rect 29165 27185 29188 27190
rect 28442 27070 28449 27153
rect 28492 27122 28495 27133
rect 28574 27132 28581 27148
rect 28583 27133 28613 27140
rect 28690 27130 28695 27155
rect 28875 27153 28879 27175
rect 28706 27133 28720 27140
rect 28492 27092 28499 27122
rect 28609 27100 28614 27130
rect 28650 27100 28657 27130
rect 28678 27100 28679 27122
rect 28690 27100 28697 27130
rect 28779 27129 28782 27139
rect 28789 27122 28792 27129
rect 28856 27123 28865 27153
rect 28875 27145 28878 27153
rect 28663 27092 28685 27100
rect 28711 27092 28718 27122
rect 28901 27113 28908 27175
rect 28920 27153 28926 27175
rect 28945 27153 28952 27175
rect 28977 27153 28982 27175
rect 29021 27153 29028 27175
rect 29033 27153 29040 27175
rect 29090 27168 29106 27175
rect 29088 27161 29103 27168
rect 28929 27145 28932 27153
rect 28942 27145 28947 27153
rect 28975 27145 28977 27153
rect 29005 27145 29012 27153
rect 29033 27145 29037 27153
rect 29088 27145 29096 27161
rect 29154 27160 29161 27170
rect 29172 27168 29188 27185
rect 29198 27168 29205 27198
rect 29219 27195 29237 27198
rect 29212 27166 29219 27190
rect 29227 27168 29237 27195
rect 29410 27193 29415 27227
rect 29447 27221 29456 27222
rect 29453 27219 29456 27221
rect 29866 27210 29881 27230
rect 29912 27227 29925 27238
rect 29950 27230 29957 27238
rect 29941 27227 29957 27230
rect 29988 27227 29998 27249
rect 29866 27200 29885 27210
rect 29892 27200 29911 27210
rect 29885 27198 29891 27200
rect 29932 27198 29935 27227
rect 29941 27208 29949 27227
rect 30015 27219 30021 27249
rect 30056 27219 30061 27249
rect 30097 27227 30098 27252
rect 30130 27227 30137 27253
rect 29937 27200 29950 27208
rect 29706 27195 29707 27196
rect 29720 27195 29722 27196
rect 29288 27190 29294 27193
rect 29172 27160 29226 27166
rect 29227 27160 29236 27168
rect 29253 27163 29269 27190
rect 29288 27163 29291 27190
rect 29294 27163 29295 27190
rect 29329 27185 29334 27193
rect 29329 27163 29345 27185
rect 29351 27163 29359 27185
rect 29253 27160 29260 27163
rect 29295 27160 29301 27163
rect 28966 27125 29017 27133
rect 28865 27105 29004 27113
rect 28492 27070 28495 27092
rect 28690 27083 28695 27092
rect 28426 27062 28478 27070
rect 28485 27062 28497 27070
rect 28541 27062 28577 27070
rect 28167 27023 28168 27033
rect 28181 27023 28188 27053
rect 28200 27025 28224 27033
rect 28225 27031 28226 27051
rect 28255 27045 28257 27053
rect 28272 27045 28303 27053
rect 28301 27039 28302 27045
rect 28240 27031 28276 27033
rect 28225 27025 28276 27031
rect 28146 27022 28162 27023
rect 28177 27022 28178 27023
rect 28057 27008 28059 27018
rect 28049 26987 28054 27003
rect 28067 26992 28069 27008
rect 28200 27007 28203 27025
rect 28212 27015 28222 27023
rect 28228 27015 28235 27017
rect 28266 27015 28269 27023
rect 28214 27013 28224 27015
rect 28208 27009 28214 27013
rect 28235 27007 28238 27015
rect 28253 27007 28266 27015
rect 28280 27013 28290 27015
rect 28301 27013 28306 27039
rect 28151 26987 28158 27007
rect 28181 26987 28188 27007
rect 28301 26987 28302 27013
rect 28442 26987 28449 27062
rect 28492 27060 28495 27062
rect 28478 27052 28485 27060
rect 28478 27030 28494 27052
rect 28510 27030 28517 27060
rect 28568 27052 28574 27060
rect 28609 27052 28614 27060
rect 28690 27057 28697 27083
rect 28690 27052 28695 27057
rect 28551 27030 28563 27052
rect 28568 27030 28569 27052
rect 28574 27030 28575 27052
rect 28614 27030 28616 27052
rect 28627 27030 28642 27052
rect 28575 27022 28581 27030
rect 28616 27022 28621 27030
rect 28678 27022 28685 27052
rect 28711 27026 28718 27052
rect 28720 27047 28728 27082
rect 28759 27060 28765 27070
rect 28769 27049 28775 27060
rect 28845 27049 28851 27052
rect 28769 27044 28770 27049
rect 28799 27030 28815 27043
rect 28799 27027 28802 27030
rect 28812 27027 28815 27030
rect 28845 27033 28860 27049
rect 28702 27022 28718 27026
rect 28492 26987 28495 27022
rect 28568 26987 28571 26995
rect 28690 26987 28695 27022
rect 28769 27013 28774 27027
rect 28845 27022 28851 27033
rect 28855 27022 28861 27031
rect 28871 27023 28878 27105
rect 28901 27093 28908 27105
rect 28900 27085 28920 27093
rect 28947 27085 28959 27093
rect 28969 27085 28983 27093
rect 28994 27085 29010 27093
rect 28901 27083 28908 27085
rect 28984 27083 28985 27085
rect 28893 27064 28900 27083
rect 28883 27053 28900 27064
rect 28920 27079 28926 27083
rect 28920 27069 28927 27079
rect 28957 27075 28959 27083
rect 28975 27075 28977 27077
rect 28982 27075 28985 27083
rect 28920 27053 28926 27069
rect 28931 27053 28937 27069
rect 28957 27053 28973 27075
rect 28975 27053 28982 27075
rect 28984 27053 29002 27075
rect 29021 27061 29022 27145
rect 29036 27135 29037 27145
rect 29093 27115 29096 27145
rect 29162 27153 29171 27160
rect 29329 27155 29367 27163
rect 29398 27155 29405 27185
rect 29410 27163 29417 27193
rect 29419 27163 29426 27185
rect 29431 27163 29435 27185
rect 29419 27155 29436 27163
rect 29519 27155 29532 27183
rect 29585 27175 29589 27183
rect 29598 27175 29599 27193
rect 29667 27185 29686 27193
rect 29706 27188 29722 27195
rect 29610 27183 29618 27185
rect 29639 27183 29646 27185
rect 29610 27175 29620 27183
rect 29639 27175 29647 27183
rect 29665 27175 29667 27177
rect 29672 27175 29674 27183
rect 29702 27175 29704 27183
rect 29706 27182 29722 27183
rect 29741 27175 29750 27183
rect 29800 27175 29806 27185
rect 29816 27175 29818 27193
rect 29885 27192 29892 27198
rect 29885 27190 29899 27192
rect 29885 27185 29908 27190
rect 29162 27070 29169 27153
rect 29212 27122 29215 27133
rect 29294 27132 29301 27148
rect 29303 27133 29333 27140
rect 29410 27130 29415 27155
rect 29595 27153 29599 27175
rect 29426 27133 29440 27140
rect 29212 27092 29219 27122
rect 29329 27100 29334 27130
rect 29370 27100 29377 27130
rect 29398 27100 29399 27122
rect 29410 27100 29417 27130
rect 29499 27129 29502 27139
rect 29509 27122 29512 27129
rect 29576 27123 29585 27153
rect 29595 27145 29598 27153
rect 29383 27092 29405 27100
rect 29431 27092 29438 27122
rect 29621 27113 29628 27175
rect 29640 27153 29646 27175
rect 29665 27153 29672 27175
rect 29697 27153 29702 27175
rect 29741 27153 29748 27175
rect 29753 27153 29760 27175
rect 29810 27168 29826 27175
rect 29808 27161 29823 27168
rect 29649 27145 29652 27153
rect 29662 27145 29667 27153
rect 29695 27145 29697 27153
rect 29725 27145 29732 27153
rect 29753 27145 29757 27153
rect 29808 27145 29816 27161
rect 29874 27160 29881 27170
rect 29892 27168 29908 27185
rect 29918 27168 29925 27198
rect 29939 27195 29957 27198
rect 29932 27166 29939 27190
rect 29947 27168 29957 27195
rect 30130 27193 30135 27227
rect 30167 27221 30176 27222
rect 30173 27219 30176 27221
rect 30426 27195 30427 27196
rect 30440 27195 30442 27196
rect 30008 27190 30014 27193
rect 29892 27160 29946 27166
rect 29947 27160 29956 27168
rect 29973 27163 29989 27190
rect 30008 27163 30011 27190
rect 30014 27163 30015 27190
rect 30049 27185 30054 27193
rect 30049 27163 30065 27185
rect 30071 27163 30079 27185
rect 29973 27160 29980 27163
rect 30015 27160 30021 27163
rect 29686 27125 29737 27133
rect 29585 27105 29724 27113
rect 29212 27070 29215 27092
rect 29410 27083 29415 27092
rect 29146 27062 29198 27070
rect 29205 27062 29217 27070
rect 29261 27062 29297 27070
rect 28887 27023 28888 27033
rect 28901 27023 28908 27053
rect 28920 27025 28944 27033
rect 28945 27031 28946 27051
rect 28975 27045 28977 27053
rect 28992 27045 29023 27053
rect 29021 27039 29022 27045
rect 28960 27031 28996 27033
rect 28945 27025 28996 27031
rect 28866 27022 28882 27023
rect 28897 27022 28898 27023
rect 28777 27008 28779 27018
rect 28769 26987 28774 27003
rect 28787 26992 28789 27008
rect 28920 27007 28923 27025
rect 28932 27015 28942 27023
rect 28948 27015 28955 27017
rect 28986 27015 28989 27023
rect 28934 27013 28944 27015
rect 28928 27009 28934 27013
rect 28955 27007 28958 27015
rect 28973 27007 28986 27015
rect 29000 27013 29010 27015
rect 29021 27013 29026 27039
rect 28871 26987 28878 27007
rect 28901 26987 28908 27007
rect 29021 26987 29022 27013
rect 29162 26987 29169 27062
rect 29212 27060 29215 27062
rect 29198 27052 29205 27060
rect 29198 27030 29214 27052
rect 29230 27030 29237 27060
rect 29288 27052 29294 27060
rect 29329 27052 29334 27060
rect 29410 27057 29417 27083
rect 29410 27052 29415 27057
rect 29271 27030 29283 27052
rect 29288 27030 29289 27052
rect 29294 27030 29295 27052
rect 29334 27030 29336 27052
rect 29347 27030 29362 27052
rect 29295 27022 29301 27030
rect 29336 27022 29341 27030
rect 29398 27022 29405 27052
rect 29431 27026 29438 27052
rect 29440 27047 29448 27082
rect 29479 27060 29485 27070
rect 29489 27049 29495 27060
rect 29565 27049 29571 27052
rect 29489 27044 29490 27049
rect 29519 27030 29535 27043
rect 29519 27027 29522 27030
rect 29532 27027 29535 27030
rect 29565 27033 29580 27049
rect 29422 27022 29438 27026
rect 29212 26987 29215 27022
rect 29288 26987 29291 26995
rect 29410 26987 29415 27022
rect 29489 27013 29494 27027
rect 29565 27022 29571 27033
rect 29575 27022 29581 27031
rect 29591 27023 29598 27105
rect 29621 27093 29628 27105
rect 29620 27085 29640 27093
rect 29667 27085 29679 27093
rect 29689 27085 29703 27093
rect 29714 27085 29730 27093
rect 29621 27083 29628 27085
rect 29704 27083 29705 27085
rect 29613 27064 29620 27083
rect 29603 27053 29620 27064
rect 29640 27079 29646 27083
rect 29640 27069 29647 27079
rect 29677 27075 29679 27083
rect 29695 27075 29697 27077
rect 29702 27075 29705 27083
rect 29640 27053 29646 27069
rect 29651 27053 29657 27069
rect 29677 27053 29693 27075
rect 29695 27053 29702 27075
rect 29704 27053 29722 27075
rect 29741 27061 29742 27145
rect 29756 27135 29757 27145
rect 29813 27115 29816 27145
rect 29882 27153 29891 27160
rect 30049 27155 30087 27163
rect 30118 27155 30125 27185
rect 30130 27163 30137 27193
rect 30139 27163 30146 27185
rect 30151 27163 30155 27185
rect 30139 27155 30156 27163
rect 30239 27155 30252 27183
rect 30305 27175 30309 27183
rect 30318 27175 30319 27193
rect 30387 27185 30406 27193
rect 30426 27188 30442 27195
rect 30330 27183 30338 27185
rect 30359 27183 30366 27185
rect 30330 27175 30340 27183
rect 30359 27175 30367 27183
rect 30385 27175 30387 27177
rect 30392 27175 30394 27183
rect 30422 27175 30424 27183
rect 30426 27182 30442 27183
rect 30461 27175 30470 27183
rect 29882 27070 29889 27153
rect 29932 27122 29935 27133
rect 30014 27132 30021 27148
rect 30023 27133 30053 27140
rect 30130 27130 30135 27155
rect 30315 27153 30319 27175
rect 30146 27133 30160 27140
rect 29932 27092 29939 27122
rect 30049 27100 30054 27130
rect 30090 27100 30097 27130
rect 30118 27100 30119 27122
rect 30130 27100 30137 27130
rect 30219 27129 30222 27139
rect 30229 27122 30232 27129
rect 30296 27123 30305 27153
rect 30315 27145 30318 27153
rect 30103 27092 30125 27100
rect 30151 27092 30158 27122
rect 30341 27113 30348 27175
rect 30360 27153 30366 27175
rect 30385 27153 30392 27175
rect 30417 27153 30422 27175
rect 30461 27153 30468 27175
rect 30473 27153 30480 27175
rect 30369 27145 30372 27153
rect 30382 27145 30387 27153
rect 30415 27145 30417 27153
rect 30445 27145 30452 27153
rect 30473 27145 30477 27153
rect 30406 27125 30457 27133
rect 30305 27105 30444 27113
rect 29932 27070 29935 27092
rect 30130 27083 30135 27092
rect 29866 27062 29918 27070
rect 29925 27062 29937 27070
rect 29981 27062 30017 27070
rect 29607 27023 29608 27033
rect 29621 27023 29628 27053
rect 29640 27025 29664 27033
rect 29665 27031 29666 27051
rect 29695 27045 29697 27053
rect 29712 27045 29743 27053
rect 29741 27039 29742 27045
rect 29680 27031 29716 27033
rect 29665 27025 29716 27031
rect 29586 27022 29602 27023
rect 29617 27022 29618 27023
rect 29497 27008 29499 27018
rect 29489 26987 29494 27003
rect 29507 26992 29509 27008
rect 29640 27007 29643 27025
rect 29652 27015 29662 27023
rect 29668 27015 29675 27017
rect 29706 27015 29709 27023
rect 29654 27013 29664 27015
rect 29648 27009 29654 27013
rect 29675 27007 29678 27015
rect 29693 27007 29706 27015
rect 29720 27013 29730 27015
rect 29741 27013 29746 27039
rect 29591 26987 29598 27007
rect 29621 26987 29628 27007
rect 29741 26987 29742 27013
rect 29882 26987 29889 27062
rect 29932 27060 29935 27062
rect 29918 27052 29925 27060
rect 29918 27030 29934 27052
rect 29950 27030 29957 27060
rect 30008 27052 30014 27060
rect 30049 27052 30054 27060
rect 30130 27057 30137 27083
rect 30130 27052 30135 27057
rect 29991 27030 30003 27052
rect 30008 27030 30009 27052
rect 30014 27030 30015 27052
rect 30054 27030 30056 27052
rect 30067 27030 30082 27052
rect 30015 27022 30021 27030
rect 30056 27022 30061 27030
rect 30118 27022 30125 27052
rect 30151 27026 30158 27052
rect 30160 27047 30168 27082
rect 30199 27060 30205 27070
rect 30209 27049 30215 27060
rect 30285 27049 30291 27052
rect 30209 27044 30210 27049
rect 30239 27030 30255 27043
rect 30239 27027 30242 27030
rect 30252 27027 30255 27030
rect 30285 27033 30300 27049
rect 30142 27022 30158 27026
rect 29932 26987 29935 27022
rect 30008 26987 30011 26995
rect 30130 26987 30135 27022
rect 30209 27013 30214 27027
rect 30285 27022 30291 27033
rect 30295 27022 30301 27031
rect 30311 27023 30318 27105
rect 30341 27093 30348 27105
rect 30340 27085 30360 27093
rect 30387 27085 30399 27093
rect 30409 27085 30423 27093
rect 30434 27085 30450 27093
rect 30341 27083 30348 27085
rect 30424 27083 30425 27085
rect 30333 27064 30340 27083
rect 30323 27053 30340 27064
rect 30360 27079 30366 27083
rect 30360 27069 30367 27079
rect 30397 27075 30399 27083
rect 30415 27075 30417 27077
rect 30422 27075 30425 27083
rect 30360 27053 30366 27069
rect 30371 27053 30377 27069
rect 30397 27053 30413 27075
rect 30415 27053 30422 27075
rect 30424 27053 30442 27075
rect 30461 27061 30462 27145
rect 30476 27135 30477 27145
rect 30482 27055 30489 27065
rect 30492 27061 30494 27296
rect 30492 27055 30500 27061
rect 30327 27023 30328 27033
rect 30341 27023 30348 27053
rect 30360 27025 30384 27033
rect 30385 27031 30386 27051
rect 30415 27045 30417 27053
rect 30432 27045 30463 27053
rect 30492 27045 30499 27055
rect 30500 27045 30509 27055
rect 30511 27045 30516 27063
rect 30461 27039 30462 27045
rect 30400 27031 30436 27033
rect 30385 27025 30436 27031
rect 30306 27022 30322 27023
rect 30337 27022 30338 27023
rect 30217 27008 30219 27018
rect 30209 26987 30214 27003
rect 30227 26992 30229 27008
rect 30360 27007 30363 27025
rect 30372 27015 30382 27023
rect 30388 27015 30395 27017
rect 30426 27015 30429 27023
rect 30374 27013 30384 27015
rect 30368 27009 30374 27013
rect 30395 27007 30398 27015
rect 30413 27007 30426 27015
rect 30440 27013 30450 27015
rect 30461 27013 30466 27039
rect 30492 27025 30498 27045
rect 30508 27035 30509 27045
rect 30506 27025 30509 27031
rect 30518 27026 30519 27035
rect 30521 27026 30528 27073
rect 30540 27031 30542 27301
rect 30546 27296 30550 27301
rect 30574 27296 30582 27304
rect 30608 27296 30610 27304
rect 30600 27096 30604 27106
rect 30612 27096 30614 27317
rect 30636 27312 30638 27317
rect 30660 27312 30662 27317
rect 30624 27304 30638 27312
rect 30652 27304 30664 27312
rect 30684 27304 30692 27312
rect 30622 27296 30624 27304
rect 30610 27066 30614 27096
rect 30518 27025 30537 27026
rect 30492 27023 30494 27025
rect 30311 26987 30318 27007
rect 30341 26987 30348 27007
rect 30461 26987 30462 27013
rect 30492 26999 30496 27023
rect 30511 26999 30512 27025
rect 30521 27021 30528 27025
rect 30516 27005 30532 27012
rect 30538 27005 30542 27031
rect 30569 27020 30572 27047
rect 30574 27025 30585 27047
rect 30587 27025 30590 27055
rect 30569 27017 30581 27020
rect 30492 26987 30494 26999
rect 30521 26988 30528 27005
rect 30540 26987 30542 27005
rect 30612 27004 30614 27066
rect 30628 27055 30635 27065
rect 30628 27047 30631 27055
rect 30628 27020 30635 27047
rect 30624 27017 30635 27020
rect 30624 27010 30631 27017
rect 30636 27010 30638 27304
rect 30650 27296 30652 27304
rect 30660 27104 30662 27304
rect 30664 27296 30666 27304
rect 30692 27296 30700 27304
rect 30655 27096 30662 27104
rect 30708 27096 30710 27317
rect 30712 27304 30720 27312
rect 30740 27304 30752 27312
rect 30756 27304 30758 27317
rect 30780 27312 30782 27317
rect 30804 27312 30806 27317
rect 30768 27304 30782 27312
rect 30796 27304 30808 27312
rect 30828 27304 30836 27312
rect 30720 27296 30728 27304
rect 30752 27296 30758 27304
rect 30744 27096 30748 27106
rect 30756 27096 30758 27296
rect 30780 27296 30784 27304
rect 30650 27095 30666 27096
rect 30641 27047 30645 27055
rect 30648 27051 30652 27061
rect 30655 27051 30658 27065
rect 30660 27051 30662 27095
rect 30704 27088 30710 27096
rect 30686 27058 30689 27088
rect 30708 27066 30711 27088
rect 30731 27066 30734 27096
rect 30754 27066 30765 27096
rect 30694 27059 30702 27066
rect 30708 27059 30710 27066
rect 30711 27061 30716 27066
rect 30711 27059 30725 27061
rect 30694 27058 30725 27059
rect 30694 27056 30695 27058
rect 30696 27056 30700 27058
rect 30708 27056 30710 27058
rect 30655 27047 30662 27051
rect 30655 27021 30666 27047
rect 30704 27040 30705 27056
rect 30706 27026 30710 27056
rect 30756 27053 30758 27066
rect 30655 27020 30662 27021
rect 30609 26987 30614 27004
rect 30628 26987 30631 27010
rect 30634 27007 30638 27010
rect 30641 27007 30646 27020
rect 30650 27017 30662 27020
rect 30634 26996 30648 27007
rect 30636 26987 30645 26996
rect 30655 26991 30662 27017
rect 30708 27004 30710 27026
rect 30753 27013 30758 27053
rect 30772 27048 30779 27066
rect 30780 27048 30782 27296
rect 30785 27088 30792 27096
rect 30804 27088 30806 27304
rect 30808 27296 30812 27304
rect 30836 27296 30844 27304
rect 30852 27096 30854 27317
rect 30856 27304 30864 27312
rect 30884 27304 30896 27312
rect 30900 27304 30902 27317
rect 30924 27312 30926 27317
rect 30948 27312 30950 27317
rect 30912 27304 30926 27312
rect 30940 27304 30952 27312
rect 30972 27304 30980 27312
rect 30864 27296 30872 27304
rect 30896 27296 30902 27304
rect 30888 27096 30892 27106
rect 30900 27096 30902 27296
rect 30924 27296 30928 27304
rect 30848 27088 30854 27096
rect 30785 27066 30789 27088
rect 30799 27061 30806 27088
rect 30792 27058 30810 27061
rect 30830 27058 30833 27088
rect 30852 27066 30855 27088
rect 30875 27066 30878 27096
rect 30898 27066 30909 27096
rect 30838 27059 30846 27066
rect 30852 27059 30854 27066
rect 30855 27061 30860 27066
rect 30855 27059 30869 27061
rect 30838 27058 30869 27059
rect 30785 27048 30789 27058
rect 30792 27051 30796 27058
rect 30772 27020 30775 27048
rect 30655 26987 30658 26991
rect 30660 26987 30662 26991
rect 30695 26994 30698 26998
rect 30695 26988 30699 26994
rect 30704 26987 30710 27004
rect 30756 26987 30758 27013
rect 30768 27010 30775 27020
rect 30780 27032 30789 27048
rect 30790 27037 30796 27047
rect 30780 27020 30782 27032
rect 30785 27020 30789 27032
rect 30799 27021 30806 27058
rect 30838 27056 30839 27058
rect 30840 27056 30844 27058
rect 30852 27056 30854 27058
rect 30848 27040 30849 27056
rect 30850 27026 30854 27056
rect 30900 27053 30902 27066
rect 30780 27018 30796 27020
rect 30780 27010 30782 27018
rect 30772 26996 30775 27010
rect 30778 26996 30784 27010
rect 30785 26996 30790 27018
rect 30759 26987 30775 26996
rect 30780 26987 30784 26996
rect 30799 26987 30802 27021
rect 30804 26987 30806 27021
rect 30852 27004 30854 27026
rect 30897 27013 30902 27053
rect 30916 27048 30923 27066
rect 30924 27048 30926 27296
rect 30929 27088 30936 27096
rect 30948 27088 30950 27304
rect 30952 27296 30956 27304
rect 30980 27296 30988 27304
rect 30996 27096 30998 27317
rect 31000 27304 31008 27312
rect 31028 27304 31040 27312
rect 31044 27304 31046 27317
rect 31068 27312 31070 27317
rect 31092 27312 31094 27317
rect 31056 27304 31070 27312
rect 31084 27304 31096 27312
rect 31116 27304 31124 27312
rect 31008 27296 31016 27304
rect 31040 27296 31046 27304
rect 31032 27096 31036 27106
rect 31044 27096 31046 27296
rect 31068 27296 31072 27304
rect 30992 27088 30998 27096
rect 30929 27066 30933 27088
rect 30943 27061 30950 27088
rect 30936 27058 30954 27061
rect 30974 27058 30977 27088
rect 30996 27066 30999 27088
rect 31019 27066 31022 27096
rect 31042 27066 31053 27096
rect 30982 27059 30990 27066
rect 30996 27059 30998 27066
rect 30999 27061 31004 27066
rect 30999 27059 31013 27061
rect 30982 27058 31013 27059
rect 30929 27048 30933 27058
rect 30936 27051 30940 27058
rect 30916 27020 30919 27048
rect 30839 26994 30842 26998
rect 30839 26988 30843 26994
rect 30848 26987 30854 27004
rect 30900 26987 30902 27013
rect 30912 27010 30919 27020
rect 30924 27032 30933 27048
rect 30934 27037 30940 27047
rect 30924 27020 30926 27032
rect 30929 27020 30933 27032
rect 30943 27021 30950 27058
rect 30982 27056 30983 27058
rect 30984 27056 30988 27058
rect 30996 27056 30998 27058
rect 30992 27040 30993 27056
rect 30994 27026 30998 27056
rect 31044 27053 31046 27066
rect 30924 27018 30940 27020
rect 30924 27010 30926 27018
rect 30916 26996 30919 27010
rect 30922 26996 30928 27010
rect 30929 26996 30934 27018
rect 30903 26987 30919 26996
rect 30924 26987 30928 26996
rect 30943 26987 30946 27021
rect 30948 26987 30950 27021
rect 30996 27004 30998 27026
rect 31041 27013 31046 27053
rect 31060 27048 31067 27066
rect 31068 27048 31070 27296
rect 31073 27088 31080 27096
rect 31092 27088 31094 27304
rect 31096 27296 31100 27304
rect 31124 27296 31132 27304
rect 31140 27096 31142 27317
rect 31144 27304 31152 27312
rect 31172 27304 31186 27312
rect 31188 27304 31190 27317
rect 31236 27312 31238 27317
rect 31725 27314 31741 27317
rect 31202 27304 31214 27312
rect 31230 27304 31242 27312
rect 31262 27304 31270 27312
rect 31290 27304 31306 27312
rect 31323 27304 31334 27312
rect 31352 27304 31362 27312
rect 31383 27304 31393 27312
rect 31412 27304 31421 27312
rect 31441 27304 31449 27312
rect 31469 27304 31477 27312
rect 31497 27304 31506 27312
rect 31525 27304 31534 27312
rect 31554 27304 31562 27312
rect 31582 27304 31590 27312
rect 31610 27304 31618 27312
rect 31638 27304 31646 27312
rect 31666 27304 31674 27312
rect 31694 27304 31702 27312
rect 31888 27309 31890 27317
rect 32076 27312 32078 27317
rect 32100 27312 32102 27317
rect 31750 27304 31758 27309
rect 31778 27304 31786 27309
rect 31152 27296 31160 27304
rect 31186 27296 31190 27304
rect 31200 27296 31202 27304
rect 31214 27296 31216 27304
rect 31228 27296 31230 27304
rect 31136 27088 31142 27096
rect 31073 27066 31077 27088
rect 31087 27061 31094 27088
rect 31080 27058 31098 27061
rect 31118 27058 31121 27088
rect 31140 27066 31143 27088
rect 31163 27066 31166 27096
rect 31126 27059 31134 27066
rect 31140 27059 31142 27066
rect 31143 27061 31148 27066
rect 31143 27059 31157 27061
rect 31126 27058 31157 27059
rect 31073 27048 31077 27058
rect 31080 27051 31084 27058
rect 31060 27020 31063 27048
rect 30983 26994 30986 26998
rect 30983 26988 30987 26994
rect 30992 26987 30998 27004
rect 31044 26987 31046 27013
rect 31056 27010 31063 27020
rect 31068 27032 31077 27048
rect 31078 27037 31084 27047
rect 31068 27020 31070 27032
rect 31073 27020 31077 27032
rect 31087 27021 31094 27058
rect 31126 27056 31127 27058
rect 31128 27056 31132 27058
rect 31140 27056 31142 27058
rect 31136 27040 31137 27056
rect 31138 27026 31142 27056
rect 31068 27018 31084 27020
rect 31068 27010 31070 27018
rect 31060 26996 31063 27010
rect 31066 26996 31072 27010
rect 31073 26996 31078 27018
rect 31047 26987 31063 26996
rect 31068 26987 31072 26996
rect 31087 26987 31090 27021
rect 31092 26987 31094 27021
rect 31140 27004 31142 27026
rect 31127 26994 31130 26998
rect 31127 26988 31131 26994
rect 31136 26987 31142 27004
rect 31188 26987 31190 27296
rect 31226 27124 31227 27279
rect 31236 27124 31238 27304
rect 31242 27296 31244 27304
rect 31270 27296 31278 27304
rect 31318 27296 31323 27304
rect 31346 27296 31352 27304
rect 31393 27296 31399 27304
rect 31421 27296 31428 27304
rect 31449 27296 31457 27304
rect 31477 27296 31485 27304
rect 31506 27296 31513 27304
rect 31534 27296 31541 27304
rect 31562 27296 31570 27304
rect 31590 27296 31598 27304
rect 31618 27296 31626 27304
rect 31646 27296 31654 27304
rect 31674 27296 31682 27304
rect 31702 27296 31710 27304
rect 31758 27293 31766 27304
rect 31786 27294 31794 27304
rect 31834 27301 31842 27309
rect 31862 27301 31870 27309
rect 31888 27301 31898 27309
rect 31918 27301 31934 27312
rect 31950 27301 31962 27312
rect 31978 27301 31990 27312
rect 32010 27304 32018 27312
rect 32038 27304 32048 27312
rect 32066 27304 32078 27312
rect 32094 27304 32104 27312
rect 32124 27304 32132 27312
rect 31842 27294 31850 27301
rect 31870 27294 31878 27301
rect 31778 27293 31794 27294
rect 31834 27293 31850 27294
rect 31862 27293 31878 27294
rect 31888 27294 31890 27301
rect 31898 27294 31906 27301
rect 31946 27296 31950 27301
rect 31974 27296 31978 27301
rect 32018 27296 32026 27304
rect 32048 27296 32054 27304
rect 32076 27296 32082 27304
rect 31888 27293 31906 27294
rect 31918 27293 31926 27294
rect 31438 27279 31571 27287
rect 31576 27279 31629 27287
rect 31586 27261 31590 27270
rect 31654 27269 31661 27278
rect 31637 27257 31643 27262
rect 31662 27257 31671 27269
rect 31633 27252 31637 27257
rect 31662 27253 31678 27257
rect 31679 27253 31682 27257
rect 31411 27238 31417 27246
rect 31448 27238 31459 27242
rect 31421 27230 31427 27238
rect 31402 27210 31417 27230
rect 31448 27227 31461 27238
rect 31486 27230 31493 27238
rect 31477 27227 31493 27230
rect 31524 27227 31534 27249
rect 31402 27200 31421 27210
rect 31428 27200 31447 27210
rect 31421 27198 31427 27200
rect 31468 27198 31471 27227
rect 31477 27208 31485 27227
rect 31551 27219 31557 27249
rect 31592 27219 31597 27249
rect 31633 27227 31634 27252
rect 31666 27227 31673 27253
rect 31473 27200 31486 27208
rect 31421 27192 31428 27198
rect 31421 27190 31435 27192
rect 31421 27185 31444 27190
rect 31346 27156 31355 27166
rect 31410 27160 31417 27170
rect 31428 27168 31444 27185
rect 31454 27168 31461 27198
rect 31475 27195 31493 27198
rect 31468 27166 31475 27190
rect 31483 27168 31493 27195
rect 31666 27193 31671 27227
rect 31703 27221 31712 27222
rect 31709 27219 31712 27221
rect 31544 27190 31550 27193
rect 31428 27160 31482 27166
rect 31483 27160 31492 27168
rect 31509 27163 31525 27190
rect 31544 27163 31547 27190
rect 31550 27163 31551 27190
rect 31585 27185 31590 27193
rect 31585 27163 31601 27185
rect 31607 27163 31615 27185
rect 31509 27160 31516 27163
rect 31551 27160 31557 27163
rect 31342 27130 31350 27132
rect 31241 27124 31242 27125
rect 31226 27118 31242 27124
rect 31226 27098 31227 27118
rect 31193 27082 31197 27096
rect 31217 27088 31219 27096
rect 31226 27090 31228 27098
rect 31224 27088 31228 27090
rect 31236 27088 31238 27118
rect 31342 27116 31349 27130
rect 31356 27116 31365 27156
rect 31418 27153 31427 27160
rect 31585 27155 31623 27163
rect 31654 27155 31661 27185
rect 31666 27163 31673 27193
rect 31888 27186 31890 27293
rect 31675 27163 31682 27185
rect 31687 27163 31691 27185
rect 31675 27155 31692 27163
rect 31776 27156 31788 27172
rect 31217 27082 31224 27088
rect 31226 27082 31242 27088
rect 31269 27082 31279 27104
rect 31224 27058 31226 27082
rect 31216 27048 31220 27056
rect 31214 27036 31220 27048
rect 31212 27032 31220 27036
rect 31214 27022 31216 27032
rect 31214 27018 31228 27022
rect 31222 27010 31228 27018
rect 31236 27010 31238 27082
rect 31241 27058 31242 27082
rect 31326 27074 31330 27114
rect 31342 27074 31349 27104
rect 31356 27100 31367 27116
rect 31418 27070 31425 27153
rect 31468 27122 31471 27133
rect 31550 27132 31557 27148
rect 31559 27133 31589 27140
rect 31666 27130 31671 27155
rect 31867 27148 31868 27164
rect 31883 27162 31891 27186
rect 31960 27164 31967 27178
rect 31682 27133 31696 27140
rect 31468 27092 31475 27122
rect 31585 27100 31590 27130
rect 31626 27100 31633 27130
rect 31654 27100 31655 27122
rect 31666 27100 31673 27130
rect 31639 27092 31661 27100
rect 31687 27092 31694 27122
rect 31745 27106 31758 27122
rect 31763 27106 31767 27136
rect 31845 27110 31861 27126
rect 31854 27101 31861 27110
rect 31866 27106 31868 27128
rect 31883 27106 31892 27146
rect 31960 27138 31969 27164
rect 31960 27128 31968 27138
rect 31960 27116 31976 27128
rect 31837 27098 31841 27101
rect 31852 27098 31868 27101
rect 31960 27098 31968 27116
rect 31468 27070 31471 27092
rect 31666 27083 31671 27092
rect 31402 27062 31454 27070
rect 31461 27062 31473 27070
rect 31517 27062 31553 27070
rect 31272 27038 31286 27046
rect 31232 26996 31238 27010
rect 31236 26987 31238 26996
rect 31418 26987 31425 27062
rect 31468 27060 31471 27062
rect 31454 27052 31461 27060
rect 31454 27030 31470 27052
rect 31486 27030 31493 27060
rect 31544 27052 31550 27060
rect 31585 27052 31590 27060
rect 31666 27057 31673 27083
rect 31666 27052 31671 27057
rect 31527 27030 31539 27052
rect 31544 27030 31545 27052
rect 31550 27030 31551 27052
rect 31590 27030 31592 27052
rect 31603 27030 31618 27052
rect 31551 27027 31557 27030
rect 31523 27022 31557 27027
rect 31592 27022 31597 27030
rect 31654 27022 31661 27052
rect 31687 27026 31694 27052
rect 31696 27047 31704 27082
rect 31775 27027 31779 27043
rect 31780 27041 31791 27043
rect 31827 27041 31833 27098
rect 31846 27071 31847 27073
rect 31854 27071 31860 27098
rect 31903 27083 31906 27091
rect 31913 27081 31916 27083
rect 31843 27041 31850 27071
rect 31856 27041 31861 27063
rect 31866 27041 31872 27063
rect 31874 27041 31881 27071
rect 31883 27041 31892 27081
rect 31893 27041 31899 27063
rect 31901 27041 31908 27071
rect 31913 27041 31919 27081
rect 31960 27073 31967 27075
rect 31790 27035 31791 27041
rect 31854 27033 31861 27041
rect 31883 27033 31891 27041
rect 31678 27022 31694 27026
rect 31468 26987 31471 27022
rect 31539 26999 31543 27015
rect 31544 26987 31547 26995
rect 31603 26991 31619 26993
rect 31666 26987 31671 27022
rect 31854 27018 31860 27033
rect 31753 27008 31761 27018
rect 31854 27013 31869 27018
rect 31763 27008 31772 27011
rect 31763 26992 31771 27008
rect 31772 26995 31779 27008
rect 31854 27003 31860 27013
rect 31884 26987 31891 27033
rect 31933 27027 31937 27057
rect 31942 27033 31949 27057
rect 31951 27033 31958 27063
rect 31960 27033 31968 27073
rect 31969 27033 31976 27057
rect 31978 27033 31985 27063
rect 32068 27057 32075 27067
rect 31945 27000 31953 27027
rect 31960 26987 31967 27033
rect 32009 27019 32012 27049
rect 32014 27027 32025 27049
rect 32027 27027 32030 27057
rect 32068 27049 32071 27057
rect 32036 27019 32040 27027
rect 32068 27020 32075 27049
rect 32064 27019 32075 27020
rect 32020 26987 32029 27019
rect 32064 27010 32071 27019
rect 32076 27010 32078 27296
rect 32081 27049 32085 27057
rect 32088 27051 32092 27061
rect 32095 27051 32098 27067
rect 32100 27051 32102 27304
rect 32104 27296 32110 27304
rect 32132 27296 32140 27304
rect 32148 27096 32150 27317
rect 32152 27304 32160 27312
rect 32160 27296 32168 27304
rect 32144 27088 32150 27096
rect 32126 27058 32129 27088
rect 32148 27066 32151 27088
rect 32171 27066 32174 27096
rect 32134 27059 32142 27066
rect 32148 27059 32150 27066
rect 32151 27061 32156 27066
rect 32151 27059 32165 27061
rect 32134 27058 32165 27059
rect 32134 27056 32135 27058
rect 32136 27056 32140 27058
rect 32148 27056 32150 27058
rect 32095 27049 32102 27051
rect 32095 27021 32106 27049
rect 32144 27040 32145 27056
rect 32146 27026 32150 27056
rect 32095 27020 32102 27021
rect 32068 26987 32071 27010
rect 32074 26996 32078 27010
rect 32081 26996 32086 27020
rect 32090 27019 32102 27020
rect 32076 26987 32078 26996
rect 32095 26987 32098 27019
rect 32100 26987 32102 27019
rect 32148 27004 32150 27026
rect 32135 26994 32138 26998
rect 32135 26988 32139 26994
rect 32144 26987 32150 27004
rect -19052 26979 32184 26987
rect -19028 26976 -19022 26979
rect -18958 26976 -18948 26977
rect -18968 26919 -18964 26969
rect -18848 26967 -18839 26969
rect -18728 26967 -18719 26969
rect -18608 26967 -18599 26969
rect -18488 26967 -18479 26969
rect -18368 26967 -18359 26969
rect -18248 26967 -18239 26969
rect -18128 26967 -18119 26969
rect -18008 26967 -17999 26969
rect -18963 26919 -18952 26959
rect -18950 26911 -18947 26959
rect -18941 26842 -18937 26967
rect -18848 26919 -18837 26967
rect -18728 26919 -18717 26967
rect -18608 26919 -18597 26967
rect -18488 26919 -18477 26967
rect -18368 26919 -18357 26967
rect -18248 26919 -18237 26967
rect -18128 26919 -18117 26967
rect -18008 26919 -17997 26967
rect -17916 26921 -17914 26979
rect -17913 26969 -17912 26979
rect -17913 26921 -17906 26969
rect -17893 26961 -17879 26969
rect -17916 26915 -17906 26921
rect -17916 26658 -17914 26915
rect -17905 26911 -17902 26915
rect -17894 26911 -17889 26959
rect -17895 26841 -17889 26851
rect -17879 26841 -17876 26851
rect -17868 26841 -17866 26979
rect -17820 26917 -17818 26979
rect -17817 26953 -17801 26964
rect -17817 26917 -17811 26953
rect -17820 26916 -17811 26917
rect -17791 26916 -17789 26964
rect -17820 26893 -17816 26916
rect -17885 26793 -17879 26841
rect -17869 26793 -17866 26841
rect -17848 26833 -17842 26841
rect -17868 26658 -17866 26793
rect -17836 26793 -17830 26833
rect -17836 26667 -17832 26793
rect -19041 26650 -19031 26658
rect -18978 26650 -18968 26658
rect -18950 26650 -18938 26658
rect -18918 26650 -18910 26658
rect -18890 26650 -18874 26658
rect -18858 26650 -18846 26658
rect -18830 26650 -18818 26658
rect -18798 26650 -18790 26658
rect -18770 26650 -18754 26658
rect -18738 26650 -18726 26658
rect -18710 26650 -18698 26658
rect -18678 26650 -18670 26658
rect -18650 26650 -18634 26658
rect -18618 26650 -18606 26658
rect -18590 26650 -18578 26658
rect -18558 26650 -18550 26658
rect -18530 26650 -18514 26658
rect -18498 26650 -18486 26658
rect -18470 26650 -18458 26658
rect -18438 26650 -18430 26658
rect -18410 26650 -18394 26658
rect -18378 26650 -18366 26658
rect -18350 26650 -18338 26658
rect -18318 26650 -18310 26658
rect -18290 26650 -18274 26658
rect -18258 26650 -18246 26658
rect -18230 26650 -18218 26658
rect -18198 26650 -18190 26658
rect -18170 26650 -18154 26658
rect -18138 26650 -18126 26658
rect -18110 26650 -18098 26658
rect -18078 26650 -18070 26658
rect -18050 26650 -18034 26658
rect -18018 26650 -18006 26658
rect -17990 26650 -17978 26658
rect -17958 26650 -17950 26658
rect -17930 26650 -17914 26658
rect -17900 26650 -17888 26658
rect -17872 26650 -17860 26658
rect -19031 26642 -19025 26650
rect -18984 26642 -18978 26650
rect -18955 26642 -18950 26650
rect -18910 26642 -18902 26650
rect -18862 26642 -18858 26650
rect -18834 26642 -18830 26650
rect -18790 26642 -18782 26650
rect -18742 26642 -18738 26650
rect -18714 26642 -18710 26650
rect -18670 26642 -18662 26650
rect -18622 26642 -18618 26650
rect -18594 26642 -18590 26650
rect -18550 26642 -18542 26650
rect -18502 26642 -18498 26650
rect -18474 26642 -18470 26650
rect -18430 26642 -18422 26650
rect -18382 26642 -18378 26650
rect -18354 26642 -18350 26650
rect -18310 26642 -18302 26650
rect -18262 26642 -18258 26650
rect -18234 26642 -18230 26650
rect -18190 26642 -18182 26650
rect -18142 26642 -18138 26650
rect -18114 26642 -18110 26650
rect -18070 26642 -18062 26650
rect -18022 26642 -18018 26650
rect -17994 26642 -17990 26650
rect -17950 26642 -17942 26650
rect -17916 26639 -17914 26650
rect -17902 26642 -17900 26650
rect -17888 26642 -17886 26650
rect -17874 26642 -17872 26650
rect -17868 26639 -17866 26650
rect -17860 26642 -17858 26650
rect -17820 26639 -17818 26893
rect -17772 26658 -17770 26979
rect -17652 26966 -17650 26979
rect -17741 26916 -17729 26956
rect -17679 26932 -17674 26956
rect -17663 26955 -17660 26965
rect -17654 26955 -17653 26956
rect -17652 26955 -17643 26966
rect -17654 26939 -17650 26955
rect -17612 26948 -17603 26979
rect -17576 26947 -17568 26956
rect -17577 26942 -17568 26947
rect -17680 26916 -17664 26932
rect -17679 26908 -17674 26916
rect -17654 26908 -17653 26939
rect -17677 26789 -17673 26847
rect -17652 26658 -17650 26939
rect -17626 26934 -17624 26939
rect -17614 26934 -17612 26939
rect -17612 26929 -17604 26934
rect -17602 26924 -17594 26929
rect -17580 26921 -17578 26934
rect -17570 26932 -17561 26942
rect -17551 26932 -17544 26979
rect -17543 26955 -17540 26965
rect -17532 26955 -17530 26979
rect -17560 26931 -17551 26932
rect -17536 26929 -17534 26942
rect -17533 26939 -17530 26955
rect -17492 26948 -17483 26979
rect -17436 26971 -17434 26979
rect -17437 26961 -17432 26971
rect -17416 26961 -17410 26979
rect -17436 26957 -17432 26961
rect -17645 26789 -17643 26919
rect -17605 26883 -17599 26909
rect -17580 26908 -17578 26911
rect -17569 26847 -17560 26911
rect -17624 26819 -17619 26847
rect -17569 26837 -17559 26847
rect -17551 26837 -17544 26916
rect -17532 26885 -17530 26939
rect -17506 26934 -17504 26939
rect -17494 26934 -17492 26939
rect -17492 26929 -17484 26934
rect -17438 26931 -17431 26957
rect -17482 26924 -17474 26929
rect -17525 26911 -17516 26919
rect -17525 26885 -17523 26901
rect -17532 26861 -17523 26885
rect -17485 26883 -17479 26909
rect -17460 26908 -17458 26911
rect -17606 26829 -17602 26837
rect -17590 26829 -17580 26837
rect -17623 26789 -17619 26819
rect -17618 26789 -17607 26829
rect -17605 26789 -17602 26829
rect -17578 26827 -17571 26837
rect -17579 26789 -17570 26827
rect -17569 26789 -17563 26829
rect -17623 26781 -17620 26789
rect -17596 26667 -17592 26789
rect -17561 26781 -17554 26829
rect -17552 26781 -17543 26837
rect -17532 26829 -17530 26861
rect -17542 26789 -17536 26829
rect -17534 26781 -17527 26829
rect -17525 26789 -17516 26839
rect -17504 26819 -17499 26847
rect -17456 26839 -17451 26841
rect -17486 26829 -17482 26837
rect -17503 26789 -17499 26819
rect -17498 26789 -17487 26829
rect -17485 26789 -17482 26829
rect -17503 26781 -17500 26789
rect -17532 26658 -17530 26781
rect -17476 26667 -17472 26789
rect -17456 26667 -17450 26839
rect -17436 26829 -17434 26931
rect -17412 26901 -17410 26961
rect -17364 26917 -17362 26979
rect -17361 26953 -17345 26964
rect -17361 26917 -17355 26953
rect -17364 26916 -17355 26917
rect -17335 26916 -17333 26964
rect -17412 26885 -17404 26901
rect -17364 26893 -17360 26916
rect -17412 26861 -17403 26885
rect -17423 26841 -17420 26851
rect -17412 26841 -17410 26861
rect -17431 26839 -17424 26841
rect -17431 26829 -17423 26839
rect -17413 26829 -17410 26841
rect -17449 26793 -17440 26829
rect -17438 26793 -17433 26829
rect -17429 26793 -17423 26829
rect -17422 26793 -17406 26829
rect -17438 26785 -17431 26793
rect -17412 26785 -17406 26793
rect -17436 26658 -17434 26785
rect -17412 26658 -17410 26785
rect -17402 26667 -17396 26839
rect -17392 26833 -17386 26841
rect -17380 26793 -17374 26833
rect -17380 26667 -17376 26793
rect -17806 26650 -17796 26658
rect -17778 26650 -17768 26658
rect -17746 26650 -17738 26658
rect -17682 26650 -17674 26658
rect -17654 26650 -17646 26658
rect -17622 26650 -17614 26658
rect -17594 26650 -17578 26658
rect -17562 26650 -17550 26658
rect -17534 26650 -17522 26658
rect -17502 26650 -17494 26658
rect -17474 26650 -17460 26658
rect -17444 26650 -17432 26658
rect -17416 26650 -17404 26658
rect -17812 26642 -17806 26650
rect -17784 26642 -17778 26650
rect -17772 26639 -17770 26650
rect -17738 26642 -17730 26650
rect -17690 26642 -17682 26650
rect -17662 26642 -17654 26650
rect -17652 26639 -17650 26650
rect -17614 26642 -17606 26650
rect -17566 26642 -17562 26650
rect -17538 26642 -17534 26650
rect -17532 26639 -17530 26650
rect -17494 26642 -17486 26650
rect -17460 26642 -17458 26650
rect -17446 26642 -17444 26650
rect -17436 26639 -17434 26650
rect -17432 26642 -17430 26650
rect -17418 26642 -17416 26650
rect -17412 26639 -17410 26650
rect -17404 26642 -17402 26650
rect -17364 26639 -17362 26893
rect -17316 26658 -17314 26979
rect -17222 26977 -17215 26979
rect -17222 26966 -17213 26977
rect -17222 26961 -17205 26966
rect -17285 26916 -17273 26956
rect -17222 26900 -17215 26961
rect -17200 26908 -17197 26956
rect -17220 26851 -17218 26900
rect -17221 26667 -17214 26851
rect -17207 26841 -17204 26851
rect -17196 26841 -17194 26979
rect -17124 26969 -17119 26979
rect -17124 26953 -17121 26969
rect -17120 26967 -17119 26969
rect -17028 26969 -17024 26979
rect -17120 26953 -17112 26967
rect -17028 26956 -17018 26969
rect -17197 26793 -17194 26841
rect -17176 26833 -17170 26841
rect -17220 26658 -17218 26667
rect -17196 26658 -17194 26793
rect -17164 26793 -17158 26833
rect -17164 26667 -17160 26793
rect -17124 26658 -17122 26953
rect -17119 26919 -17112 26953
rect -17030 26942 -17026 26956
rect -17093 26667 -17084 26843
rect -17028 26658 -17026 26942
rect -17017 26942 -17016 26956
rect -17009 26942 -17002 26959
rect -16991 26955 -16988 26965
rect -16980 26955 -16978 26979
rect -17017 26932 -17002 26942
rect -16981 26939 -16978 26955
rect -16940 26948 -16931 26979
rect -16884 26971 -16882 26979
rect -16885 26961 -16880 26971
rect -16864 26961 -16858 26979
rect -16884 26957 -16880 26961
rect -17017 26916 -17001 26932
rect -17017 26911 -17002 26916
rect -17017 26847 -17008 26911
rect -17017 26837 -17001 26847
rect -17000 26667 -16991 26837
rect -16980 26658 -16978 26939
rect -16954 26934 -16952 26939
rect -16942 26934 -16940 26939
rect -16940 26929 -16932 26934
rect -16886 26931 -16879 26957
rect -16930 26924 -16922 26929
rect -16933 26883 -16927 26909
rect -16908 26908 -16906 26911
rect -16952 26819 -16947 26847
rect -16904 26839 -16899 26841
rect -16934 26829 -16930 26837
rect -16951 26789 -16947 26819
rect -16946 26789 -16935 26829
rect -16933 26789 -16930 26829
rect -16951 26781 -16948 26789
rect -16924 26667 -16920 26789
rect -16904 26667 -16898 26839
rect -16884 26829 -16882 26931
rect -16860 26901 -16858 26961
rect -16822 26915 -16819 26925
rect -16812 26917 -16810 26979
rect -16799 26977 -16794 26979
rect -16790 26953 -16783 26979
rect -16860 26885 -16852 26901
rect -16812 26893 -16808 26917
rect -16860 26861 -16851 26885
rect -16871 26841 -16868 26851
rect -16860 26841 -16858 26861
rect -16879 26839 -16872 26841
rect -16879 26829 -16871 26839
rect -16861 26829 -16858 26841
rect -16897 26793 -16888 26829
rect -16886 26793 -16881 26829
rect -16877 26793 -16871 26829
rect -16870 26793 -16854 26829
rect -16886 26785 -16879 26793
rect -16860 26785 -16854 26793
rect -16884 26658 -16882 26785
rect -16860 26658 -16858 26785
rect -16850 26667 -16844 26839
rect -16840 26833 -16834 26841
rect -16828 26793 -16822 26833
rect -16828 26667 -16824 26793
rect -17350 26650 -17340 26658
rect -17322 26650 -17312 26658
rect -17290 26650 -17282 26658
rect -17228 26650 -17218 26658
rect -17200 26650 -17190 26658
rect -17130 26650 -17122 26658
rect -17102 26650 -17096 26658
rect -17070 26650 -17062 26658
rect -17042 26650 -17026 26658
rect -17010 26650 -16998 26658
rect -16982 26650 -16970 26658
rect -16950 26650 -16942 26658
rect -16922 26650 -16908 26658
rect -16892 26650 -16880 26658
rect -16864 26650 -16852 26658
rect -17356 26642 -17350 26650
rect -17328 26642 -17322 26650
rect -17316 26639 -17314 26650
rect -17282 26642 -17274 26650
rect -17234 26642 -17228 26650
rect -17220 26639 -17218 26650
rect -17206 26642 -17200 26650
rect -17196 26639 -17194 26650
rect -17140 26642 -17130 26650
rect -17124 26639 -17122 26650
rect -17112 26642 -17102 26650
rect -17062 26642 -17054 26650
rect -17028 26639 -17026 26650
rect -17014 26642 -17010 26650
rect -16986 26642 -16982 26650
rect -16980 26639 -16978 26650
rect -16942 26642 -16934 26650
rect -16908 26642 -16906 26650
rect -16894 26642 -16892 26650
rect -16884 26639 -16882 26650
rect -16880 26642 -16878 26650
rect -16866 26642 -16864 26650
rect -16860 26639 -16858 26650
rect -16852 26642 -16850 26650
rect -16812 26639 -16810 26893
rect -16808 26667 -16802 26841
rect -16788 26833 -16786 26953
rect -16775 26841 -16772 26851
rect -16764 26841 -16762 26979
rect -16726 26915 -16723 26925
rect -16716 26917 -16714 26979
rect -16703 26977 -16698 26979
rect -16694 26953 -16687 26979
rect -16716 26893 -16712 26917
rect -16783 26833 -16775 26841
rect -16765 26833 -16762 26841
rect -16801 26793 -16792 26833
rect -16790 26793 -16785 26833
rect -16781 26793 -16775 26833
rect -16774 26793 -16758 26833
rect -16790 26785 -16783 26793
rect -16764 26785 -16758 26793
rect -16788 26658 -16786 26785
rect -16764 26658 -16762 26785
rect -16754 26667 -16748 26841
rect -16744 26833 -16738 26841
rect -16732 26793 -16726 26833
rect -16732 26667 -16728 26793
rect -16796 26650 -16786 26658
rect -16768 26650 -16760 26658
rect -16804 26642 -16796 26650
rect -16788 26639 -16786 26650
rect -16776 26642 -16768 26650
rect -16764 26639 -16762 26650
rect -16716 26639 -16714 26893
rect -16712 26667 -16706 26841
rect -16692 26833 -16690 26953
rect -16679 26841 -16676 26851
rect -16668 26841 -16666 26979
rect -16604 26969 -16601 26979
rect -16596 26953 -16587 26979
rect -16633 26931 -16627 26941
rect -16604 26931 -16601 26953
rect -16623 26903 -16611 26931
rect -16618 26883 -16611 26903
rect -16596 26893 -16594 26953
rect -16603 26883 -16594 26893
rect -16687 26833 -16679 26841
rect -16669 26833 -16666 26841
rect -16705 26793 -16696 26833
rect -16694 26793 -16689 26833
rect -16685 26793 -16679 26833
rect -16678 26793 -16662 26833
rect -16694 26785 -16687 26793
rect -16668 26785 -16662 26793
rect -16692 26658 -16690 26785
rect -16668 26658 -16666 26785
rect -16658 26667 -16652 26841
rect -16648 26833 -16642 26841
rect -16604 26833 -16594 26883
rect -16591 26931 -16587 26953
rect -16528 26933 -16523 26979
rect -16591 26883 -16584 26931
rect -16558 26923 -16548 26931
rect -16547 26883 -16533 26923
rect -16528 26883 -16520 26933
rect -16500 26931 -16492 26979
rect -16490 26949 -16488 26953
rect -16482 26949 -16481 26979
rect -16415 26977 -16414 26979
rect -16404 26977 -16390 26979
rect -16405 26966 -16389 26977
rect -16380 26966 -16376 26979
rect -16405 26961 -16402 26966
rect -16483 26935 -16464 26941
rect -16483 26934 -16482 26935
rect -16491 26933 -16482 26934
rect -16482 26931 -16481 26933
rect -16500 26928 -16482 26931
rect -16500 26923 -16491 26928
rect -16500 26883 -16492 26923
rect -16591 26833 -16587 26883
rect -16540 26875 -16533 26883
rect -16509 26875 -16502 26883
rect -16500 26875 -16498 26883
rect -16482 26875 -16475 26923
rect -16473 26883 -16472 26923
rect -16464 26883 -16457 26931
rect -16438 26915 -16436 26925
rect -16428 26901 -16426 26915
rect -16452 26875 -16447 26883
rect -16528 26868 -16523 26875
rect -16528 26858 -16521 26868
rect -16514 26866 -16508 26868
rect -16515 26858 -16508 26866
rect -16500 26867 -16492 26875
rect -16482 26867 -16481 26875
rect -16500 26858 -16498 26867
rect -16636 26793 -16630 26833
rect -16604 26807 -16597 26833
rect -16596 26807 -16594 26833
rect -16528 26832 -16523 26858
rect -16520 26856 -16508 26858
rect -16504 26856 -16498 26858
rect -16520 26842 -16511 26856
rect -16505 26842 -16498 26856
rect -16604 26800 -16579 26807
rect -16570 26806 -16566 26818
rect -16528 26806 -16523 26816
rect -16500 26806 -16498 26842
rect -16424 26834 -16412 26841
rect -16497 26806 -16493 26809
rect -16465 26808 -16464 26809
rect -16461 26806 -16457 26808
rect -16636 26667 -16632 26793
rect -16596 26791 -16579 26800
rect -16700 26650 -16690 26658
rect -16672 26650 -16664 26658
rect -16612 26650 -16607 26658
rect -16596 26650 -16594 26791
rect -16558 26785 -16554 26806
rect -16528 26799 -16520 26806
rect -16528 26792 -16503 26799
rect -16558 26758 -16556 26785
rect -16527 26667 -16520 26792
rect -16519 26783 -16503 26792
rect -16500 26798 -16493 26806
rect -16470 26803 -16457 26806
rect -16500 26784 -16498 26798
rect -16482 26784 -16475 26798
rect -16500 26783 -16493 26784
rect -16500 26658 -16498 26783
rect -16482 26758 -16474 26784
rect -16473 26758 -16466 26798
rect -16464 26758 -16457 26803
rect -16424 26798 -16421 26834
rect -16404 26798 -16402 26961
rect -16384 26875 -16381 26923
rect -16391 26841 -16388 26851
rect -16380 26841 -16378 26966
rect -16342 26915 -16339 26925
rect -16332 26917 -16330 26979
rect -16319 26977 -16314 26979
rect -16310 26953 -16303 26979
rect -16332 26893 -16328 26917
rect -16381 26798 -16378 26841
rect -16360 26833 -16354 26841
rect -16424 26793 -16408 26798
rect -16406 26793 -16399 26798
rect -16397 26793 -16378 26798
rect -16482 26750 -16475 26758
rect -16451 26667 -16447 26758
rect -16404 26658 -16402 26793
rect -16384 26780 -16381 26793
rect -16380 26658 -16378 26793
rect -16348 26793 -16342 26833
rect -16348 26667 -16344 26793
rect -16584 26650 -16579 26658
rect -16531 26650 -16523 26658
rect -16503 26650 -16495 26658
rect -16475 26650 -16467 26658
rect -16412 26650 -16402 26658
rect -16384 26650 -16375 26658
rect -16708 26642 -16700 26650
rect -16692 26639 -16690 26650
rect -16680 26642 -16672 26650
rect -16668 26639 -16666 26650
rect -16607 26642 -16594 26650
rect -16579 26642 -16568 26650
rect -16523 26642 -16515 26650
rect -16596 26639 -16594 26642
rect -16500 26639 -16498 26650
rect -16495 26642 -16487 26650
rect -16467 26642 -16459 26650
rect -16419 26642 -16412 26650
rect -16404 26639 -16402 26650
rect -16391 26642 -16384 26650
rect -16380 26639 -16378 26650
rect -16332 26639 -16330 26893
rect -16328 26667 -16322 26841
rect -16308 26833 -16306 26953
rect -16295 26841 -16292 26851
rect -16284 26841 -16282 26979
rect -16246 26915 -16243 26925
rect -16236 26917 -16234 26979
rect -16223 26977 -16218 26979
rect -16214 26953 -16207 26979
rect -16236 26893 -16232 26917
rect -16303 26833 -16295 26841
rect -16285 26833 -16282 26841
rect -16321 26793 -16312 26833
rect -16310 26793 -16305 26833
rect -16301 26793 -16295 26833
rect -16294 26793 -16278 26833
rect -16310 26785 -16303 26793
rect -16284 26785 -16278 26793
rect -16308 26658 -16306 26785
rect -16284 26658 -16282 26785
rect -16274 26667 -16268 26841
rect -16264 26833 -16258 26841
rect -16252 26793 -16246 26833
rect -16252 26667 -16248 26793
rect -16316 26650 -16306 26658
rect -16288 26650 -16280 26658
rect -16324 26642 -16316 26650
rect -16308 26639 -16306 26650
rect -16296 26642 -16288 26650
rect -16284 26639 -16282 26650
rect -16236 26639 -16234 26893
rect -16232 26667 -16226 26841
rect -16212 26833 -16210 26953
rect -16199 26841 -16196 26851
rect -16188 26841 -16186 26979
rect -16142 26893 -16123 26902
rect -16030 26882 -16023 26979
rect -15980 26976 -15977 26979
rect -15904 26968 -15901 26979
rect -15863 26970 -15860 26979
rect -15845 26978 -15759 26979
rect -15810 26960 -15807 26961
rect -16000 26952 -15994 26960
rect -15987 26952 -15973 26960
rect -15913 26952 -15904 26953
rect -15844 26952 -15842 26960
rect -15835 26952 -15801 26960
rect -15980 26950 -15977 26952
rect -15904 26950 -15901 26952
rect -15994 26902 -15987 26950
rect -15984 26902 -15983 26942
rect -15999 26894 -15990 26902
rect -15980 26894 -15973 26942
rect -15962 26902 -15955 26950
rect -15911 26947 -15897 26950
rect -15904 26942 -15897 26947
rect -15923 26902 -15920 26942
rect -15968 26894 -15923 26902
rect -15918 26894 -15911 26942
rect -15903 26894 -15897 26942
rect -15846 26902 -15844 26942
rect -15842 26902 -15835 26950
rect -15815 26947 -15794 26950
rect -15801 26942 -15794 26947
rect -15748 26942 -15744 26978
rect -15827 26902 -15826 26942
rect -15877 26894 -15870 26902
rect -15824 26894 -15817 26942
rect -15813 26902 -15809 26942
rect -15801 26902 -15797 26942
rect -15770 26902 -15769 26942
rect -15794 26894 -15787 26902
rect -15761 26894 -15754 26942
rect -15980 26882 -15977 26894
rect -15904 26892 -15897 26894
rect -15904 26882 -15901 26892
rect -16040 26874 -15968 26882
rect -15923 26874 -15846 26882
rect -16030 26872 -16023 26874
rect -16020 26856 -16016 26862
rect -16207 26833 -16199 26841
rect -16189 26833 -16186 26841
rect -16225 26793 -16216 26833
rect -16214 26793 -16209 26833
rect -16205 26793 -16199 26833
rect -16198 26793 -16182 26833
rect -16214 26785 -16207 26793
rect -16188 26785 -16182 26793
rect -16212 26658 -16210 26785
rect -16188 26658 -16186 26785
rect -16178 26667 -16172 26841
rect -16168 26833 -16162 26841
rect -16156 26793 -16150 26833
rect -16156 26667 -16152 26793
rect -16132 26667 -16130 26843
rect -16104 26824 -16099 26833
rect -16129 26785 -16116 26824
rect -16106 26785 -16104 26824
rect -16102 26785 -16099 26824
rect -16096 26785 -16086 26824
rect -16030 26816 -16023 26856
rect -15980 26841 -15977 26874
rect -15976 26864 -15973 26874
rect -15966 26854 -15963 26864
rect -15966 26848 -15950 26854
rect -15922 26848 -15910 26854
rect -16008 26824 -16004 26834
rect -15994 26826 -15972 26834
rect -15994 26825 -15978 26826
rect -15904 26824 -15901 26874
rect -15878 26854 -15756 26859
rect -15852 26839 -15834 26846
rect -15897 26826 -15877 26834
rect -15748 26826 -15744 26894
rect -15998 26820 -15980 26824
rect -16111 26777 -16106 26785
rect -16038 26768 -16031 26816
rect -15998 26776 -15992 26820
rect -15962 26776 -15955 26824
rect -15904 26816 -15896 26824
rect -15842 26816 -15835 26824
rect -15922 26776 -15920 26816
rect -16020 26768 -16004 26775
rect -15998 26768 -15994 26776
rect -15918 26768 -15911 26816
rect -15903 26768 -15896 26816
rect -15860 26777 -15852 26816
rect -15860 26776 -15844 26777
rect -16030 26705 -16023 26768
rect -15904 26765 -15896 26768
rect -15877 26765 -15870 26776
rect -15852 26768 -15844 26776
rect -15824 26768 -15817 26816
rect -15815 26776 -15811 26816
rect -15801 26776 -15799 26824
rect -15794 26768 -15787 26816
rect -15782 26778 -15776 26816
rect -15748 26778 -15741 26826
rect -15739 26778 -15735 26816
rect -15761 26768 -15754 26778
rect -15678 26771 -15674 26818
rect -15605 26815 -15602 26841
rect -15594 26815 -15588 26979
rect -15564 26824 -15557 26979
rect -15430 26915 -15427 26925
rect -15420 26917 -15418 26979
rect -15407 26977 -15402 26979
rect -15398 26953 -15391 26979
rect -15420 26893 -15416 26917
rect -15660 26783 -15659 26813
rect -15613 26805 -15611 26815
rect -15594 26805 -15587 26815
rect -15574 26805 -15567 26824
rect -15551 26823 -15539 26824
rect -15552 26807 -15539 26823
rect -15603 26789 -15601 26805
rect -15584 26789 -15567 26805
rect -15678 26770 -15661 26771
rect -15792 26767 -15789 26768
rect -15748 26767 -15744 26768
rect -16016 26747 -15980 26755
rect -15904 26753 -15901 26765
rect -15594 26763 -15588 26789
rect -15582 26776 -15567 26789
rect -15547 26776 -15540 26807
rect -15512 26793 -15511 26841
rect -15487 26826 -15481 26841
rect -15448 26833 -15442 26841
rect -15487 26816 -15480 26826
rect -15506 26793 -15496 26816
rect -15494 26793 -15490 26816
rect -15488 26793 -15487 26816
rect -15485 26793 -15480 26816
rect -15479 26793 -15469 26816
rect -15494 26785 -15488 26793
rect -15467 26785 -15463 26816
rect -15928 26747 -15880 26753
rect -15822 26747 -15811 26755
rect -15981 26737 -15980 26747
rect -15956 26745 -15955 26747
rect -15962 26737 -15955 26745
rect -15904 26743 -15901 26747
rect -16030 26697 -16014 26705
rect -16040 26685 -16032 26695
rect -16030 26689 -16021 26697
rect -16006 26687 -16004 26715
rect -15981 26689 -15973 26737
rect -15956 26697 -15955 26737
rect -15935 26689 -15928 26737
rect -15918 26727 -15902 26737
rect -15842 26735 -15835 26745
rect -15792 26735 -15786 26755
rect -15778 26737 -15769 26745
rect -15766 26737 -15759 26755
rect -15714 26747 -15697 26755
rect -15687 26747 -15674 26755
rect -15676 26746 -15674 26747
rect -15842 26719 -15826 26735
rect -15864 26693 -15858 26699
rect -15766 26697 -15757 26737
rect -15704 26697 -15693 26737
rect -15675 26697 -15674 26746
rect -15621 26737 -15615 26755
rect -15609 26747 -15601 26759
rect -15564 26755 -15557 26776
rect -15598 26751 -15574 26755
rect -15567 26751 -15556 26755
rect -15598 26747 -15585 26751
rect -15609 26745 -15599 26747
rect -15594 26745 -15588 26747
rect -15564 26745 -15557 26751
rect -15546 26745 -15539 26747
rect -15605 26742 -15594 26745
rect -15587 26742 -15580 26745
rect -15605 26737 -15596 26742
rect -15575 26737 -15566 26745
rect -15547 26737 -15539 26745
rect -15533 26737 -15529 26751
rect -15628 26697 -15625 26737
rect -15623 26697 -15616 26737
rect -15612 26697 -15608 26737
rect -15605 26697 -15598 26737
rect -15593 26697 -15586 26737
rect -15582 26697 -15577 26737
rect -15574 26697 -15567 26737
rect -15565 26697 -15556 26737
rect -15555 26697 -15549 26737
rect -15547 26697 -15540 26737
rect -15868 26689 -15864 26693
rect -15802 26685 -15796 26695
rect -15766 26689 -15759 26697
rect -15628 26689 -15608 26697
rect -15594 26689 -15587 26697
rect -15565 26689 -15557 26697
rect -15536 26689 -15529 26737
rect -15512 26689 -15510 26747
rect -16030 26677 -16022 26685
rect -15792 26677 -15786 26685
rect -15562 26677 -15559 26689
rect -16030 26669 -15914 26677
rect -15792 26669 -15785 26677
rect -15769 26669 -15751 26677
rect -15735 26669 -15720 26677
rect -15562 26669 -15555 26677
rect -15539 26669 -15512 26677
rect -15496 26669 -15493 26677
rect -15458 26667 -15453 26826
rect -15436 26793 -15430 26833
rect -15436 26667 -15432 26793
rect -16220 26650 -16210 26658
rect -16192 26650 -16184 26658
rect -16122 26650 -16116 26658
rect -16094 26650 -16088 26658
rect -16062 26650 -16054 26658
rect -16034 26650 -16026 26658
rect -16006 26650 -15998 26658
rect -15978 26650 -15970 26658
rect -15967 26656 -15954 26658
rect -15950 26650 -15942 26658
rect -15922 26650 -15914 26658
rect -15909 26656 -15898 26658
rect -15894 26650 -15886 26658
rect -15866 26650 -15858 26658
rect -15838 26650 -15830 26658
rect -15810 26650 -15802 26658
rect -15782 26650 -15774 26658
rect -15754 26656 -15736 26658
rect -15754 26650 -15746 26656
rect -15698 26650 -15692 26661
rect -15670 26650 -15664 26661
rect -15628 26653 -15620 26661
rect -15616 26653 -15608 26661
rect -15600 26653 -15592 26661
rect -15588 26653 -15580 26661
rect -15572 26653 -15564 26661
rect -15560 26653 -15552 26661
rect -15544 26653 -15536 26661
rect -15532 26653 -15516 26658
rect -15500 26653 -15488 26658
rect -15472 26653 -15460 26658
rect -15616 26652 -15600 26653
rect -15588 26652 -15572 26653
rect -15560 26652 -15544 26653
rect -15532 26652 -15524 26653
rect -16228 26642 -16220 26650
rect -16212 26639 -16210 26650
rect -16200 26642 -16192 26650
rect -16188 26639 -16186 26650
rect -16132 26642 -16122 26650
rect -16104 26642 -16094 26650
rect -16054 26642 -16046 26650
rect -16026 26642 -16018 26650
rect -15998 26642 -15990 26650
rect -15970 26642 -15962 26650
rect -15942 26642 -15934 26650
rect -15914 26642 -15906 26650
rect -15886 26642 -15878 26650
rect -15858 26642 -15850 26650
rect -15830 26642 -15822 26650
rect -15802 26642 -15794 26650
rect -15774 26642 -15766 26650
rect -15746 26642 -15738 26650
rect -15692 26645 -15682 26650
rect -15664 26645 -15654 26650
rect -15608 26645 -15600 26652
rect -15580 26645 -15572 26652
rect -15552 26645 -15544 26652
rect -15504 26642 -15500 26653
rect -15476 26642 -15472 26653
rect -16056 26639 -16020 26642
rect -15670 26639 -15636 26641
rect -15420 26639 -15418 26893
rect -15416 26667 -15410 26841
rect -15396 26833 -15394 26953
rect -15383 26841 -15380 26851
rect -15372 26841 -15370 26979
rect -15300 26969 -15295 26979
rect -15300 26953 -15297 26969
rect -15296 26967 -15295 26969
rect -15176 26967 -15167 26969
rect -15296 26953 -15288 26967
rect -15391 26833 -15383 26841
rect -15373 26833 -15370 26841
rect -15409 26793 -15400 26833
rect -15398 26793 -15393 26833
rect -15389 26793 -15383 26833
rect -15382 26793 -15366 26833
rect -15398 26785 -15391 26793
rect -15372 26785 -15366 26793
rect -15396 26658 -15394 26785
rect -15372 26658 -15370 26785
rect -15362 26667 -15356 26841
rect -15352 26833 -15346 26841
rect -15340 26793 -15334 26833
rect -15340 26667 -15336 26793
rect -15300 26658 -15298 26953
rect -15295 26919 -15288 26953
rect -15176 26919 -15165 26967
rect -15269 26667 -15260 26843
rect -15404 26650 -15394 26658
rect -15376 26650 -15368 26658
rect -15306 26650 -15298 26658
rect -15278 26650 -15272 26658
rect -15246 26650 -15238 26658
rect -15218 26650 -15202 26658
rect -15186 26650 -15174 26658
rect -15158 26650 -15146 26658
rect -15126 26650 -15118 26658
rect -15098 26650 -15086 26658
rect -15084 26650 -15082 26979
rect -15076 26964 -15074 26969
rect -15081 26916 -15074 26964
rect -15073 26916 -15057 26959
rect -15058 26911 -15057 26916
rect -15036 26658 -15034 26979
rect -14942 26977 -14935 26979
rect -14942 26966 -14933 26977
rect -14942 26961 -14925 26966
rect -15005 26916 -14993 26956
rect -14942 26900 -14935 26961
rect -14920 26908 -14917 26956
rect -14940 26851 -14938 26900
rect -14941 26667 -14934 26851
rect -14927 26841 -14924 26851
rect -14916 26841 -14914 26979
rect -14868 26917 -14866 26979
rect -14865 26953 -14849 26964
rect -14865 26917 -14859 26953
rect -14868 26916 -14859 26917
rect -14839 26916 -14837 26964
rect -14868 26893 -14864 26916
rect -14917 26793 -14914 26841
rect -14896 26833 -14890 26841
rect -14940 26658 -14938 26667
rect -14916 26658 -14914 26793
rect -14884 26793 -14878 26833
rect -14884 26667 -14880 26793
rect -15070 26650 -15058 26658
rect -15042 26650 -15030 26658
rect -15010 26650 -15002 26658
rect -14948 26650 -14938 26658
rect -14920 26650 -14910 26658
rect -15412 26642 -15404 26650
rect -15396 26639 -15394 26650
rect -15384 26642 -15376 26650
rect -15372 26639 -15370 26650
rect -15316 26642 -15306 26650
rect -15300 26639 -15298 26650
rect -15288 26642 -15278 26650
rect -15238 26642 -15230 26650
rect -15190 26642 -15186 26650
rect -15162 26642 -15158 26650
rect -15118 26642 -15110 26650
rect -15086 26642 -15082 26650
rect -15058 26642 -15054 26650
rect -15084 26639 -15082 26642
rect -15036 26639 -15034 26650
rect -15030 26642 -15026 26650
rect -15002 26642 -14994 26650
rect -14954 26642 -14948 26650
rect -14940 26639 -14938 26650
rect -14926 26642 -14920 26650
rect -14916 26639 -14914 26650
rect -14868 26639 -14866 26893
rect -14820 26658 -14818 26979
rect -14726 26977 -14719 26979
rect -14726 26966 -14717 26977
rect -14726 26961 -14709 26966
rect -14789 26916 -14777 26956
rect -14726 26900 -14719 26961
rect -14704 26908 -14701 26956
rect -14724 26851 -14722 26900
rect -14725 26667 -14718 26851
rect -14711 26841 -14708 26851
rect -14700 26841 -14698 26979
rect -14664 26956 -14659 26966
rect -14652 26956 -14649 26979
rect -14654 26953 -14640 26956
rect -14654 26942 -14649 26953
rect -14652 26917 -14649 26942
rect -14623 26932 -14616 26979
rect -14615 26955 -14612 26965
rect -14604 26955 -14602 26979
rect -14605 26939 -14602 26955
rect -14564 26948 -14555 26979
rect -14508 26971 -14506 26979
rect -14509 26961 -14504 26971
rect -14488 26961 -14482 26979
rect -14508 26957 -14504 26961
rect -14652 26893 -14648 26917
rect -14701 26793 -14698 26841
rect -14680 26833 -14674 26841
rect -14652 26837 -14650 26893
rect -14635 26847 -14632 26893
rect -14635 26837 -14625 26847
rect -14623 26837 -14616 26916
rect -14662 26833 -14643 26837
rect -14724 26658 -14722 26667
rect -14700 26658 -14698 26793
rect -14668 26793 -14662 26833
rect -14652 26827 -14643 26833
rect -14668 26667 -14664 26793
rect -14652 26789 -14642 26827
rect -14641 26789 -14635 26833
rect -14854 26650 -14844 26658
rect -14826 26650 -14816 26658
rect -14794 26650 -14786 26658
rect -14732 26650 -14722 26658
rect -14704 26650 -14694 26658
rect -14860 26642 -14854 26650
rect -14832 26642 -14826 26650
rect -14820 26639 -14818 26650
rect -14786 26642 -14778 26650
rect -14738 26642 -14732 26650
rect -14724 26639 -14722 26650
rect -14710 26642 -14704 26650
rect -14700 26639 -14698 26650
rect -14652 26639 -14650 26789
rect -14633 26785 -14626 26833
rect -14624 26785 -14615 26837
rect -14604 26833 -14602 26939
rect -14578 26934 -14576 26939
rect -14566 26934 -14564 26939
rect -14564 26929 -14556 26934
rect -14510 26931 -14503 26957
rect -14554 26924 -14546 26929
rect -14557 26883 -14551 26909
rect -14532 26908 -14530 26911
rect -14614 26789 -14608 26833
rect -14606 26785 -14599 26833
rect -14597 26789 -14588 26843
rect -14576 26819 -14571 26847
rect -14528 26839 -14523 26841
rect -14558 26829 -14554 26837
rect -14575 26789 -14571 26819
rect -14570 26789 -14559 26829
rect -14557 26789 -14554 26829
rect -14623 26781 -14616 26785
rect -14604 26658 -14602 26785
rect -14575 26781 -14572 26789
rect -14548 26667 -14544 26789
rect -14528 26667 -14522 26839
rect -14508 26829 -14506 26931
rect -14484 26901 -14482 26961
rect -14448 26956 -14443 26966
rect -14436 26956 -14433 26979
rect -14438 26953 -14424 26956
rect -14438 26942 -14433 26953
rect -14436 26917 -14433 26942
rect -14407 26932 -14400 26979
rect -14399 26955 -14396 26965
rect -14388 26955 -14386 26979
rect -14389 26939 -14386 26955
rect -14348 26948 -14339 26979
rect -14312 26947 -14304 26956
rect -14313 26942 -14304 26947
rect -14484 26885 -14476 26901
rect -14436 26893 -14432 26917
rect -14484 26861 -14475 26885
rect -14495 26841 -14492 26851
rect -14484 26841 -14482 26861
rect -14503 26839 -14496 26841
rect -14503 26829 -14495 26839
rect -14485 26829 -14482 26841
rect -14521 26793 -14512 26829
rect -14510 26793 -14505 26829
rect -14501 26793 -14495 26829
rect -14494 26793 -14478 26829
rect -14510 26785 -14503 26793
rect -14484 26785 -14478 26793
rect -14508 26658 -14506 26785
rect -14484 26658 -14482 26785
rect -14474 26667 -14468 26839
rect -14464 26833 -14458 26841
rect -14436 26837 -14434 26893
rect -14419 26847 -14416 26893
rect -14419 26837 -14409 26847
rect -14407 26837 -14400 26916
rect -14446 26833 -14427 26837
rect -14452 26793 -14446 26833
rect -14436 26827 -14427 26833
rect -14452 26667 -14448 26793
rect -14436 26789 -14426 26827
rect -14425 26789 -14419 26833
rect -14634 26650 -14628 26658
rect -14606 26650 -14600 26658
rect -14574 26650 -14566 26658
rect -14546 26650 -14532 26658
rect -14516 26650 -14504 26658
rect -14488 26650 -14476 26658
rect -14644 26642 -14634 26650
rect -14616 26642 -14606 26650
rect -14604 26639 -14602 26650
rect -14566 26642 -14558 26650
rect -14532 26642 -14530 26650
rect -14518 26642 -14516 26650
rect -14508 26639 -14506 26650
rect -14504 26642 -14502 26650
rect -14490 26642 -14488 26650
rect -14484 26639 -14482 26650
rect -14476 26642 -14474 26650
rect -14436 26639 -14434 26789
rect -14417 26785 -14410 26833
rect -14408 26785 -14399 26837
rect -14388 26833 -14386 26939
rect -14362 26934 -14360 26939
rect -14350 26934 -14348 26939
rect -14348 26929 -14340 26934
rect -14338 26924 -14330 26929
rect -14316 26921 -14314 26934
rect -14306 26932 -14297 26942
rect -14287 26932 -14280 26979
rect -14279 26955 -14276 26965
rect -14268 26955 -14266 26979
rect -14296 26931 -14287 26932
rect -14272 26929 -14270 26942
rect -14269 26939 -14266 26955
rect -14228 26948 -14219 26979
rect -14172 26971 -14170 26979
rect -14152 26977 -14148 26979
rect -14172 26957 -14168 26971
rect -14152 26967 -14142 26977
rect -14167 26957 -14160 26967
rect -14172 26947 -14160 26957
rect -14341 26883 -14335 26909
rect -14316 26908 -14314 26911
rect -14305 26847 -14296 26911
rect -14398 26789 -14392 26833
rect -14390 26785 -14383 26833
rect -14381 26789 -14372 26843
rect -14360 26819 -14355 26847
rect -14305 26837 -14295 26847
rect -14287 26837 -14280 26916
rect -14268 26885 -14266 26939
rect -14242 26934 -14240 26939
rect -14230 26934 -14228 26939
rect -14228 26929 -14220 26934
rect -14218 26924 -14210 26929
rect -14261 26911 -14252 26919
rect -14261 26885 -14259 26901
rect -14268 26861 -14259 26885
rect -14221 26883 -14215 26909
rect -14342 26829 -14338 26837
rect -14326 26829 -14316 26837
rect -14359 26789 -14355 26819
rect -14354 26789 -14343 26829
rect -14341 26789 -14338 26829
rect -14314 26827 -14307 26837
rect -14315 26789 -14306 26827
rect -14305 26789 -14299 26829
rect -14407 26781 -14400 26785
rect -14388 26658 -14386 26785
rect -14359 26781 -14356 26789
rect -14332 26667 -14328 26789
rect -14297 26781 -14290 26829
rect -14288 26781 -14279 26837
rect -14268 26829 -14266 26861
rect -14278 26789 -14272 26829
rect -14270 26781 -14263 26829
rect -14261 26789 -14252 26839
rect -14240 26819 -14235 26847
rect -14222 26829 -14218 26837
rect -14239 26789 -14235 26819
rect -14234 26789 -14223 26829
rect -14221 26789 -14218 26829
rect -14239 26781 -14236 26789
rect -14268 26658 -14266 26781
rect -14212 26667 -14208 26789
rect -14172 26658 -14170 26947
rect -14168 26931 -14160 26947
rect -14167 26919 -14160 26931
rect -14141 26911 -14132 26967
rect -14076 26921 -14074 26979
rect -14073 26969 -14072 26979
rect -14073 26921 -14066 26969
rect -14053 26961 -14039 26969
rect -14076 26915 -14066 26921
rect -14141 26861 -14139 26901
rect -14141 26667 -14132 26839
rect -14076 26658 -14074 26915
rect -14065 26911 -14062 26915
rect -14054 26911 -14049 26959
rect -14055 26841 -14049 26851
rect -14039 26841 -14036 26851
rect -14028 26841 -14026 26979
rect -13990 26915 -13987 26925
rect -13980 26917 -13978 26979
rect -13967 26977 -13962 26979
rect -13958 26953 -13951 26979
rect -13980 26893 -13976 26917
rect -14045 26793 -14039 26841
rect -14029 26793 -14026 26841
rect -14008 26833 -14002 26841
rect -14028 26658 -14026 26793
rect -13996 26793 -13990 26833
rect -13996 26667 -13992 26793
rect -14418 26650 -14412 26658
rect -14390 26650 -14384 26658
rect -14358 26650 -14350 26658
rect -14330 26650 -14314 26658
rect -14298 26650 -14286 26658
rect -14270 26650 -14258 26658
rect -14238 26650 -14230 26658
rect -14210 26650 -14194 26658
rect -14178 26650 -14166 26658
rect -14150 26650 -14138 26658
rect -14118 26650 -14110 26658
rect -14090 26650 -14074 26658
rect -14060 26650 -14048 26658
rect -14032 26650 -14020 26658
rect -14428 26642 -14418 26650
rect -14400 26642 -14390 26650
rect -14388 26639 -14386 26650
rect -14350 26642 -14342 26650
rect -14302 26642 -14298 26650
rect -14274 26642 -14270 26650
rect -14268 26639 -14266 26650
rect -14230 26642 -14222 26650
rect -14182 26642 -14178 26650
rect -14172 26639 -14170 26650
rect -14154 26642 -14150 26650
rect -14110 26642 -14102 26650
rect -14076 26639 -14074 26650
rect -14062 26642 -14060 26650
rect -14048 26642 -14046 26650
rect -14034 26642 -14032 26650
rect -14028 26639 -14026 26650
rect -14020 26642 -14018 26650
rect -13980 26639 -13978 26893
rect -13976 26667 -13970 26841
rect -13956 26833 -13954 26953
rect -13943 26841 -13940 26851
rect -13932 26841 -13930 26979
rect -13860 26969 -13855 26979
rect -13860 26953 -13857 26969
rect -13856 26967 -13855 26969
rect -13764 26969 -13760 26979
rect -13856 26953 -13848 26967
rect -13951 26833 -13943 26841
rect -13933 26833 -13930 26841
rect -13969 26793 -13960 26833
rect -13958 26793 -13953 26833
rect -13949 26793 -13943 26833
rect -13942 26793 -13926 26833
rect -13958 26785 -13951 26793
rect -13932 26785 -13926 26793
rect -13956 26658 -13954 26785
rect -13932 26658 -13930 26785
rect -13922 26667 -13916 26841
rect -13912 26833 -13906 26841
rect -13900 26793 -13894 26833
rect -13900 26667 -13896 26793
rect -13860 26658 -13858 26953
rect -13855 26919 -13848 26953
rect -13764 26959 -13754 26969
rect -13764 26913 -13762 26959
rect -13777 26911 -13762 26913
rect -13777 26903 -13772 26911
rect -13764 26903 -13762 26911
rect -13753 26911 -13738 26959
rect -13727 26953 -13724 26963
rect -13716 26953 -13714 26979
rect -13656 26956 -13652 26966
rect -13644 26956 -13642 26979
rect -13717 26937 -13714 26953
rect -13646 26942 -13642 26956
rect -13640 26945 -13632 26956
rect -13641 26942 -13632 26945
rect -13753 26903 -13744 26911
rect -13767 26889 -13762 26903
rect -13829 26667 -13820 26843
rect -13964 26650 -13954 26658
rect -13936 26650 -13928 26658
rect -13866 26650 -13858 26658
rect -13838 26650 -13832 26658
rect -13806 26650 -13798 26658
rect -13778 26650 -13766 26658
rect -13764 26650 -13762 26889
rect -13746 26839 -13737 26849
rect -13736 26667 -13727 26839
rect -13716 26658 -13714 26937
rect -13701 26895 -13699 26899
rect -13691 26881 -13689 26895
rect -13687 26791 -13683 26849
rect -13670 26831 -13666 26839
rect -13644 26837 -13642 26942
rect -13634 26932 -13625 26942
rect -13615 26932 -13608 26979
rect -13606 26977 -13604 26979
rect -13607 26955 -13604 26965
rect -13596 26955 -13594 26979
rect -13597 26939 -13594 26955
rect -13556 26948 -13547 26979
rect -13500 26971 -13498 26979
rect -13480 26977 -13476 26979
rect -13500 26957 -13496 26971
rect -13480 26967 -13470 26977
rect -13495 26957 -13488 26967
rect -13500 26947 -13488 26957
rect -13624 26929 -13615 26932
rect -13633 26847 -13624 26881
rect -13633 26837 -13623 26847
rect -13615 26837 -13608 26916
rect -13654 26831 -13635 26837
rect -13682 26791 -13671 26831
rect -13669 26791 -13666 26831
rect -13644 26827 -13635 26831
rect -13687 26783 -13684 26791
rect -13660 26667 -13656 26791
rect -13644 26789 -13634 26827
rect -13633 26789 -13627 26831
rect -13750 26650 -13738 26658
rect -13722 26650 -13710 26658
rect -13690 26650 -13682 26658
rect -13972 26642 -13964 26650
rect -13956 26639 -13954 26650
rect -13944 26642 -13936 26650
rect -13932 26639 -13930 26650
rect -13876 26642 -13866 26650
rect -13860 26639 -13858 26650
rect -13848 26642 -13838 26650
rect -13798 26642 -13790 26650
rect -13766 26642 -13762 26650
rect -13738 26642 -13734 26650
rect -13764 26639 -13762 26642
rect -13716 26639 -13714 26650
rect -13710 26642 -13706 26650
rect -13682 26642 -13674 26650
rect -13644 26639 -13642 26789
rect -13625 26783 -13618 26831
rect -13616 26783 -13607 26837
rect -13596 26831 -13594 26939
rect -13570 26934 -13568 26939
rect -13558 26934 -13556 26939
rect -13556 26929 -13548 26934
rect -13546 26924 -13538 26929
rect -13549 26883 -13543 26909
rect -13606 26789 -13600 26831
rect -13598 26783 -13591 26831
rect -13589 26789 -13580 26841
rect -13568 26819 -13563 26847
rect -13550 26829 -13546 26837
rect -13567 26789 -13563 26819
rect -13562 26789 -13551 26829
rect -13549 26789 -13546 26829
rect -13615 26781 -13608 26783
rect -13596 26658 -13594 26783
rect -13567 26781 -13564 26789
rect -13540 26667 -13536 26789
rect -13500 26658 -13498 26947
rect -13496 26931 -13488 26947
rect -13495 26919 -13488 26931
rect -13469 26911 -13460 26967
rect -13404 26921 -13402 26979
rect -13401 26969 -13400 26979
rect -13401 26921 -13394 26969
rect -13381 26961 -13367 26969
rect -13404 26915 -13394 26921
rect -13469 26861 -13467 26901
rect -13469 26667 -13460 26839
rect -13404 26658 -13402 26915
rect -13393 26911 -13390 26915
rect -13382 26911 -13377 26959
rect -13383 26841 -13377 26851
rect -13367 26841 -13364 26851
rect -13356 26841 -13354 26979
rect -13284 26969 -13279 26979
rect -13284 26953 -13281 26969
rect -13280 26967 -13279 26969
rect -13160 26967 -13151 26969
rect -13040 26967 -13031 26969
rect -12920 26967 -12911 26969
rect -13280 26953 -13272 26967
rect -13373 26793 -13367 26841
rect -13357 26793 -13354 26841
rect -13336 26833 -13330 26841
rect -13356 26658 -13354 26793
rect -13324 26793 -13318 26833
rect -13324 26667 -13320 26793
rect -13284 26658 -13282 26953
rect -13279 26919 -13272 26953
rect -13160 26919 -13149 26967
rect -13040 26919 -13029 26967
rect -12920 26919 -12909 26967
rect -13253 26667 -13244 26843
rect -13626 26650 -13618 26658
rect -13598 26650 -13590 26658
rect -13566 26650 -13558 26658
rect -13538 26650 -13522 26658
rect -13506 26650 -13494 26658
rect -13478 26650 -13466 26658
rect -13446 26650 -13438 26658
rect -13418 26650 -13402 26658
rect -13388 26650 -13376 26658
rect -13360 26650 -13348 26658
rect -13290 26650 -13282 26658
rect -13262 26650 -13256 26658
rect -13230 26650 -13222 26658
rect -13202 26650 -13186 26658
rect -13170 26650 -13158 26658
rect -13142 26650 -13130 26658
rect -13110 26650 -13102 26658
rect -13082 26650 -13066 26658
rect -13050 26650 -13038 26658
rect -13022 26650 -13010 26658
rect -12990 26650 -12982 26658
rect -12962 26650 -12946 26658
rect -12930 26650 -12918 26658
rect -12902 26650 -12890 26658
rect -12870 26650 -12862 26658
rect -12842 26650 -12830 26658
rect -12828 26650 -12826 26979
rect -12820 26964 -12818 26969
rect -12825 26916 -12818 26964
rect -12817 26916 -12801 26959
rect -12802 26911 -12801 26916
rect -12780 26658 -12778 26979
rect -12686 26977 -12679 26979
rect -12686 26966 -12677 26977
rect -12686 26961 -12669 26966
rect -12749 26916 -12737 26956
rect -12686 26900 -12679 26961
rect -12664 26908 -12661 26956
rect -12684 26851 -12682 26900
rect -12685 26667 -12678 26851
rect -12671 26841 -12668 26851
rect -12660 26841 -12658 26979
rect -12622 26915 -12619 26925
rect -12612 26917 -12610 26979
rect -12599 26977 -12594 26979
rect -12590 26953 -12583 26979
rect -12612 26893 -12608 26917
rect -12661 26793 -12658 26841
rect -12640 26833 -12634 26841
rect -12684 26658 -12682 26667
rect -12660 26658 -12658 26793
rect -12628 26793 -12622 26833
rect -12628 26667 -12624 26793
rect -12814 26650 -12802 26658
rect -12786 26650 -12774 26658
rect -12754 26650 -12746 26658
rect -12692 26650 -12682 26658
rect -12664 26650 -12654 26658
rect -13634 26642 -13626 26650
rect -13606 26642 -13598 26650
rect -13596 26639 -13594 26650
rect -13558 26642 -13550 26650
rect -13510 26642 -13506 26650
rect -13500 26639 -13498 26650
rect -13482 26642 -13478 26650
rect -13438 26642 -13430 26650
rect -13404 26639 -13402 26650
rect -13390 26642 -13388 26650
rect -13376 26642 -13374 26650
rect -13362 26642 -13360 26650
rect -13356 26639 -13354 26650
rect -13348 26642 -13346 26650
rect -13300 26642 -13290 26650
rect -13284 26639 -13282 26650
rect -13272 26642 -13262 26650
rect -13222 26642 -13214 26650
rect -13174 26642 -13170 26650
rect -13146 26642 -13142 26650
rect -13102 26642 -13094 26650
rect -13054 26642 -13050 26650
rect -13026 26642 -13022 26650
rect -12982 26642 -12974 26650
rect -12934 26642 -12930 26650
rect -12906 26642 -12902 26650
rect -12862 26642 -12854 26650
rect -12830 26642 -12826 26650
rect -12802 26642 -12798 26650
rect -12828 26639 -12826 26642
rect -12780 26639 -12778 26650
rect -12774 26642 -12770 26650
rect -12746 26642 -12738 26650
rect -12698 26642 -12692 26650
rect -12684 26639 -12682 26650
rect -12670 26642 -12664 26650
rect -12660 26639 -12658 26650
rect -12612 26639 -12610 26893
rect -12608 26667 -12602 26841
rect -12588 26833 -12586 26953
rect -12575 26841 -12572 26851
rect -12564 26841 -12562 26979
rect -12492 26969 -12487 26979
rect -12492 26953 -12489 26969
rect -12488 26967 -12487 26969
rect -12396 26969 -12392 26979
rect -12488 26953 -12480 26967
rect -12583 26833 -12575 26841
rect -12565 26833 -12562 26841
rect -12601 26793 -12592 26833
rect -12590 26793 -12585 26833
rect -12581 26793 -12575 26833
rect -12574 26793 -12558 26833
rect -12590 26785 -12583 26793
rect -12564 26785 -12558 26793
rect -12588 26658 -12586 26785
rect -12564 26658 -12562 26785
rect -12554 26667 -12548 26841
rect -12544 26833 -12538 26841
rect -12532 26793 -12526 26833
rect -12532 26667 -12528 26793
rect -12492 26658 -12490 26953
rect -12487 26919 -12480 26953
rect -12396 26959 -12386 26969
rect -12396 26913 -12394 26959
rect -12409 26911 -12394 26913
rect -12409 26903 -12404 26911
rect -12396 26903 -12394 26911
rect -12385 26911 -12370 26959
rect -12359 26953 -12356 26963
rect -12348 26953 -12346 26979
rect -12349 26937 -12346 26953
rect -12385 26903 -12376 26911
rect -12399 26889 -12394 26903
rect -12461 26667 -12452 26843
rect -12596 26650 -12586 26658
rect -12568 26650 -12560 26658
rect -12498 26650 -12490 26658
rect -12470 26650 -12464 26658
rect -12438 26650 -12430 26658
rect -12410 26650 -12398 26658
rect -12396 26650 -12394 26889
rect -12378 26839 -12369 26849
rect -12368 26667 -12359 26839
rect -12348 26658 -12346 26937
rect -12333 26895 -12331 26899
rect -12323 26881 -12321 26895
rect -12319 26791 -12315 26849
rect -12302 26831 -12298 26839
rect -12314 26791 -12303 26831
rect -12301 26791 -12298 26831
rect -12319 26783 -12316 26791
rect -12292 26667 -12288 26791
rect -12382 26650 -12370 26658
rect -12354 26650 -12342 26658
rect -12322 26650 -12314 26658
rect -12604 26642 -12596 26650
rect -12588 26639 -12586 26650
rect -12576 26642 -12568 26650
rect -12564 26639 -12562 26650
rect -12508 26642 -12498 26650
rect -12492 26639 -12490 26650
rect -12480 26642 -12470 26650
rect -12430 26642 -12422 26650
rect -12398 26642 -12394 26650
rect -12370 26642 -12366 26650
rect -12396 26639 -12394 26642
rect -12348 26639 -12346 26650
rect -12342 26642 -12338 26650
rect -12314 26642 -12306 26650
rect -12276 26639 -12274 26979
rect -12252 26977 -12238 26979
rect -12252 26969 -12250 26977
rect -12253 26961 -12248 26969
rect -12252 26955 -12248 26961
rect -12254 26929 -12247 26955
rect -12272 26667 -12266 26841
rect -12252 26831 -12250 26929
rect -12239 26841 -12236 26851
rect -12228 26841 -12226 26979
rect -12156 26969 -12151 26979
rect -12156 26953 -12153 26969
rect -12152 26967 -12151 26969
rect -12152 26953 -12144 26967
rect -12247 26831 -12239 26841
rect -12229 26831 -12226 26841
rect -12265 26793 -12256 26831
rect -12254 26793 -12249 26831
rect -12245 26793 -12239 26831
rect -12238 26793 -12222 26831
rect -12254 26785 -12247 26793
rect -12228 26785 -12222 26793
rect -12252 26658 -12250 26785
rect -12228 26658 -12226 26785
rect -12218 26667 -12212 26841
rect -12208 26833 -12202 26841
rect -12196 26793 -12190 26833
rect -12196 26667 -12192 26793
rect -12156 26658 -12154 26953
rect -12151 26919 -12144 26953
rect -12125 26667 -12116 26843
rect -12260 26650 -12250 26658
rect -12232 26650 -12222 26658
rect -12162 26650 -12154 26658
rect -12134 26650 -12128 26658
rect -12102 26650 -12094 26658
rect -12074 26650 -12062 26658
rect -12060 26650 -12058 26979
rect -12052 26964 -12050 26969
rect -12057 26916 -12050 26964
rect -12049 26916 -12033 26959
rect -12034 26911 -12033 26916
rect -12012 26658 -12010 26979
rect -11918 26977 -11911 26979
rect -11918 26966 -11909 26977
rect -11918 26961 -11901 26966
rect -11981 26916 -11969 26956
rect -11918 26900 -11911 26961
rect -11896 26908 -11893 26956
rect -11916 26851 -11914 26900
rect -11917 26667 -11910 26851
rect -11903 26841 -11900 26851
rect -11892 26841 -11890 26979
rect -11844 26917 -11842 26979
rect -11841 26953 -11825 26964
rect -11841 26917 -11835 26953
rect -11844 26916 -11835 26917
rect -11815 26916 -11813 26964
rect -11844 26893 -11840 26916
rect -11893 26793 -11890 26841
rect -11872 26833 -11866 26841
rect -11916 26658 -11914 26667
rect -11892 26658 -11890 26793
rect -11860 26793 -11854 26833
rect -11860 26667 -11856 26793
rect -12046 26650 -12034 26658
rect -12018 26650 -12006 26658
rect -11986 26650 -11978 26658
rect -11924 26650 -11914 26658
rect -11896 26650 -11886 26658
rect -12266 26642 -12260 26650
rect -12252 26639 -12250 26650
rect -12238 26642 -12232 26650
rect -12228 26639 -12226 26650
rect -12172 26642 -12162 26650
rect -12156 26639 -12154 26650
rect -12144 26642 -12134 26650
rect -12094 26642 -12086 26650
rect -12062 26642 -12058 26650
rect -12034 26642 -12030 26650
rect -12060 26639 -12058 26642
rect -12012 26639 -12010 26650
rect -12006 26642 -12002 26650
rect -11978 26642 -11970 26650
rect -11930 26642 -11924 26650
rect -11916 26639 -11914 26650
rect -11902 26642 -11896 26650
rect -11892 26639 -11890 26650
rect -11844 26639 -11842 26893
rect -11796 26658 -11794 26979
rect -11765 26916 -11753 26956
rect -11710 26916 -11703 26964
rect -11701 26916 -11695 26956
rect -11693 26908 -11686 26956
rect -11676 26658 -11674 26979
rect -11581 26972 -11578 26979
rect -11580 26956 -11578 26972
rect -11556 26966 -11554 26979
rect -11645 26916 -11633 26956
rect -11583 26908 -11578 26956
rect -11567 26953 -11564 26963
rect -11558 26953 -11557 26956
rect -11556 26953 -11547 26966
rect -11558 26937 -11554 26953
rect -11558 26908 -11557 26937
rect -11580 26849 -11578 26908
rect -11581 26791 -11577 26849
rect -11580 26658 -11578 26791
rect -11556 26658 -11554 26937
rect -11541 26895 -11539 26899
rect -11549 26791 -11547 26889
rect -11531 26881 -11529 26895
rect -11527 26791 -11523 26849
rect -11510 26831 -11506 26839
rect -11522 26791 -11511 26831
rect -11509 26791 -11506 26831
rect -11527 26783 -11524 26791
rect -11500 26667 -11496 26791
rect -11830 26650 -11820 26658
rect -11802 26650 -11792 26658
rect -11770 26650 -11762 26658
rect -11742 26650 -11726 26658
rect -11710 26650 -11698 26658
rect -11682 26650 -11670 26658
rect -11650 26650 -11642 26658
rect -11622 26650 -11606 26658
rect -11590 26650 -11578 26658
rect -11562 26650 -11550 26658
rect -11530 26650 -11522 26658
rect -11836 26642 -11830 26650
rect -11808 26642 -11802 26650
rect -11796 26639 -11794 26650
rect -11762 26642 -11754 26650
rect -11714 26642 -11710 26650
rect -11686 26642 -11682 26650
rect -11676 26639 -11674 26650
rect -11642 26642 -11634 26650
rect -11594 26642 -11590 26650
rect -11580 26639 -11578 26650
rect -11566 26642 -11562 26650
rect -11556 26639 -11554 26650
rect -11522 26642 -11514 26650
rect -11484 26639 -11482 26979
rect -11460 26977 -11446 26979
rect -11460 26969 -11458 26977
rect -11461 26961 -11456 26969
rect -11460 26955 -11456 26961
rect -11462 26929 -11455 26955
rect -11480 26667 -11474 26841
rect -11460 26831 -11458 26929
rect -11447 26841 -11444 26851
rect -11436 26841 -11434 26979
rect -11398 26915 -11395 26925
rect -11388 26917 -11386 26979
rect -11375 26977 -11370 26979
rect -11366 26953 -11359 26979
rect -11388 26893 -11384 26917
rect -11455 26831 -11447 26841
rect -11437 26831 -11434 26841
rect -11473 26793 -11464 26831
rect -11462 26793 -11457 26831
rect -11453 26793 -11447 26831
rect -11446 26793 -11430 26831
rect -11462 26785 -11455 26793
rect -11436 26785 -11430 26793
rect -11460 26658 -11458 26785
rect -11436 26658 -11434 26785
rect -11426 26667 -11420 26841
rect -11416 26833 -11410 26841
rect -11404 26793 -11398 26833
rect -11404 26667 -11400 26793
rect -11468 26650 -11458 26658
rect -11440 26650 -11430 26658
rect -11474 26642 -11468 26650
rect -11460 26639 -11458 26650
rect -11446 26642 -11440 26650
rect -11436 26639 -11434 26650
rect -11388 26639 -11386 26893
rect -11384 26667 -11378 26841
rect -11364 26833 -11362 26953
rect -11351 26841 -11348 26851
rect -11340 26841 -11338 26979
rect -11268 26969 -11263 26979
rect -11268 26953 -11265 26969
rect -11264 26967 -11263 26969
rect -11264 26953 -11256 26967
rect -11359 26833 -11351 26841
rect -11341 26833 -11338 26841
rect -11377 26793 -11368 26833
rect -11366 26793 -11361 26833
rect -11357 26793 -11351 26833
rect -11350 26793 -11334 26833
rect -11366 26785 -11359 26793
rect -11340 26785 -11334 26793
rect -11364 26658 -11362 26785
rect -11340 26658 -11338 26785
rect -11330 26667 -11324 26841
rect -11320 26833 -11314 26841
rect -11308 26793 -11302 26833
rect -11308 26667 -11304 26793
rect -11268 26658 -11266 26953
rect -11263 26919 -11256 26953
rect -11172 26921 -11170 26979
rect -11169 26969 -11168 26979
rect -11169 26921 -11162 26969
rect -11149 26961 -11135 26969
rect -11172 26915 -11162 26921
rect -11237 26667 -11228 26843
rect -11172 26658 -11170 26915
rect -11161 26911 -11158 26915
rect -11150 26911 -11145 26959
rect -11151 26841 -11145 26851
rect -11135 26841 -11132 26851
rect -11124 26841 -11122 26979
rect -11088 26956 -11083 26966
rect -11076 26956 -11073 26979
rect -11078 26953 -11064 26956
rect -11078 26942 -11073 26953
rect -11076 26917 -11073 26942
rect -11047 26932 -11040 26979
rect -11039 26955 -11036 26965
rect -11028 26955 -11026 26979
rect -11029 26939 -11026 26955
rect -10988 26948 -10979 26979
rect -10932 26971 -10930 26979
rect -10912 26977 -10908 26979
rect -10932 26957 -10928 26971
rect -10912 26967 -10902 26977
rect -10927 26957 -10920 26967
rect -10932 26947 -10920 26957
rect -11076 26893 -11072 26917
rect -11141 26793 -11135 26841
rect -11125 26793 -11122 26841
rect -11104 26833 -11098 26841
rect -11076 26837 -11074 26893
rect -11059 26847 -11056 26893
rect -11059 26837 -11049 26847
rect -11047 26837 -11040 26916
rect -11086 26833 -11067 26837
rect -11124 26658 -11122 26793
rect -11092 26793 -11086 26833
rect -11076 26827 -11067 26833
rect -11092 26667 -11088 26793
rect -11076 26789 -11066 26827
rect -11065 26789 -11059 26833
rect -11372 26650 -11362 26658
rect -11344 26650 -11336 26658
rect -11274 26650 -11266 26658
rect -11246 26650 -11240 26658
rect -11214 26650 -11206 26658
rect -11186 26650 -11170 26658
rect -11156 26650 -11144 26658
rect -11128 26650 -11116 26658
rect -11380 26642 -11372 26650
rect -11364 26639 -11362 26650
rect -11352 26642 -11344 26650
rect -11340 26639 -11338 26650
rect -11284 26642 -11274 26650
rect -11268 26639 -11266 26650
rect -11256 26642 -11246 26650
rect -11206 26642 -11198 26650
rect -11172 26639 -11170 26650
rect -11158 26642 -11156 26650
rect -11144 26642 -11142 26650
rect -11130 26642 -11128 26650
rect -11124 26639 -11122 26650
rect -11116 26642 -11114 26650
rect -11076 26639 -11074 26789
rect -11057 26785 -11050 26833
rect -11048 26785 -11039 26837
rect -11028 26833 -11026 26939
rect -11002 26934 -11000 26939
rect -10990 26934 -10988 26939
rect -10988 26929 -10980 26934
rect -10978 26924 -10970 26929
rect -10981 26883 -10975 26909
rect -11038 26789 -11032 26833
rect -11030 26785 -11023 26833
rect -11021 26789 -11012 26843
rect -11000 26819 -10995 26847
rect -10982 26829 -10978 26837
rect -10999 26789 -10995 26819
rect -10994 26789 -10983 26829
rect -10981 26789 -10978 26829
rect -11047 26781 -11040 26785
rect -11028 26658 -11026 26785
rect -10999 26781 -10996 26789
rect -10972 26667 -10968 26789
rect -10932 26658 -10930 26947
rect -10928 26931 -10920 26947
rect -10927 26919 -10920 26931
rect -10901 26911 -10892 26967
rect -10901 26861 -10899 26901
rect -10901 26667 -10892 26839
rect -11058 26650 -11052 26658
rect -11030 26650 -11024 26658
rect -10998 26650 -10990 26658
rect -10970 26650 -10954 26658
rect -10938 26650 -10926 26658
rect -10910 26650 -10898 26658
rect -10878 26650 -10870 26658
rect -10850 26650 -10838 26658
rect -10836 26650 -10834 26979
rect -10828 26964 -10826 26969
rect -10833 26916 -10826 26964
rect -10825 26916 -10809 26959
rect -10810 26911 -10809 26916
rect -10788 26658 -10786 26979
rect -10757 26916 -10745 26956
rect -10702 26916 -10695 26964
rect -10693 26916 -10687 26956
rect -10685 26908 -10678 26956
rect -10668 26658 -10666 26979
rect -10637 26916 -10625 26956
rect -10562 26908 -10555 26956
rect -10486 26882 -10479 26979
rect -10436 26976 -10433 26979
rect -10360 26968 -10357 26979
rect -10319 26970 -10316 26979
rect -10301 26978 -10215 26979
rect -10266 26960 -10263 26961
rect -10456 26952 -10450 26960
rect -10443 26952 -10429 26960
rect -10369 26952 -10360 26953
rect -10300 26952 -10298 26960
rect -10291 26952 -10257 26960
rect -10436 26950 -10433 26952
rect -10360 26950 -10357 26952
rect -10450 26902 -10443 26950
rect -10440 26902 -10439 26942
rect -10455 26894 -10446 26902
rect -10436 26894 -10429 26942
rect -10418 26902 -10411 26950
rect -10367 26947 -10353 26950
rect -10360 26942 -10353 26947
rect -10379 26902 -10376 26942
rect -10424 26894 -10379 26902
rect -10374 26894 -10367 26942
rect -10359 26894 -10353 26942
rect -10302 26902 -10300 26942
rect -10298 26902 -10291 26950
rect -10271 26947 -10250 26950
rect -10257 26942 -10250 26947
rect -10204 26942 -10200 26978
rect -10283 26902 -10282 26942
rect -10333 26894 -10326 26902
rect -10280 26894 -10273 26942
rect -10269 26902 -10265 26942
rect -10257 26902 -10253 26942
rect -10226 26902 -10225 26942
rect -10250 26894 -10243 26902
rect -10217 26894 -10210 26942
rect -10436 26882 -10433 26894
rect -10360 26892 -10353 26894
rect -10360 26882 -10357 26892
rect -10496 26874 -10424 26882
rect -10379 26874 -10302 26882
rect -10486 26872 -10479 26874
rect -10476 26856 -10472 26862
rect -10486 26816 -10479 26856
rect -10436 26841 -10433 26874
rect -10432 26864 -10429 26874
rect -10422 26854 -10419 26864
rect -10422 26848 -10406 26854
rect -10378 26848 -10366 26854
rect -10464 26824 -10460 26834
rect -10450 26826 -10428 26834
rect -10450 26825 -10434 26826
rect -10360 26824 -10357 26874
rect -10334 26854 -10212 26859
rect -10308 26839 -10290 26846
rect -10353 26826 -10333 26834
rect -10204 26826 -10200 26894
rect -10454 26820 -10436 26824
rect -10494 26768 -10487 26816
rect -10454 26776 -10448 26820
rect -10418 26776 -10411 26824
rect -10360 26816 -10352 26824
rect -10298 26816 -10291 26824
rect -10378 26776 -10376 26816
rect -10476 26768 -10460 26775
rect -10454 26768 -10450 26776
rect -10374 26768 -10367 26816
rect -10359 26768 -10352 26816
rect -10316 26777 -10308 26816
rect -10316 26776 -10300 26777
rect -10486 26705 -10479 26768
rect -10360 26765 -10352 26768
rect -10333 26765 -10326 26776
rect -10308 26768 -10300 26776
rect -10280 26768 -10273 26816
rect -10271 26776 -10267 26816
rect -10257 26776 -10255 26824
rect -10250 26768 -10243 26816
rect -10238 26778 -10232 26816
rect -10204 26778 -10197 26826
rect -10195 26778 -10191 26816
rect -10217 26768 -10210 26778
rect -10134 26771 -10130 26818
rect -10061 26815 -10058 26841
rect -10050 26815 -10044 26979
rect -10020 26824 -10013 26979
rect -9876 26917 -9874 26979
rect -9873 26953 -9857 26964
rect -9873 26917 -9867 26953
rect -9876 26916 -9867 26917
rect -9847 26916 -9845 26964
rect -9876 26893 -9872 26916
rect -10116 26783 -10115 26813
rect -10069 26805 -10067 26815
rect -10050 26805 -10043 26815
rect -10030 26805 -10023 26824
rect -10007 26823 -9995 26824
rect -10008 26807 -9995 26823
rect -10059 26789 -10057 26805
rect -10040 26789 -10023 26805
rect -10134 26770 -10117 26771
rect -10248 26767 -10245 26768
rect -10204 26767 -10200 26768
rect -10472 26747 -10436 26755
rect -10360 26753 -10357 26765
rect -10050 26763 -10044 26789
rect -10038 26776 -10023 26789
rect -10003 26776 -9996 26807
rect -9968 26793 -9967 26841
rect -9943 26826 -9937 26841
rect -9904 26833 -9898 26841
rect -9943 26816 -9936 26826
rect -9962 26793 -9952 26816
rect -9950 26793 -9946 26816
rect -9944 26793 -9943 26816
rect -9941 26793 -9936 26816
rect -9935 26793 -9925 26816
rect -9950 26785 -9944 26793
rect -9923 26785 -9919 26816
rect -10384 26747 -10336 26753
rect -10278 26747 -10267 26755
rect -10437 26737 -10436 26747
rect -10412 26745 -10411 26747
rect -10418 26737 -10411 26745
rect -10360 26743 -10357 26747
rect -10486 26697 -10470 26705
rect -10496 26685 -10488 26695
rect -10486 26689 -10477 26697
rect -10462 26687 -10460 26715
rect -10437 26689 -10429 26737
rect -10412 26697 -10411 26737
rect -10391 26689 -10384 26737
rect -10374 26727 -10358 26737
rect -10298 26735 -10291 26745
rect -10248 26735 -10242 26755
rect -10234 26737 -10225 26745
rect -10222 26737 -10215 26755
rect -10170 26747 -10153 26755
rect -10143 26747 -10130 26755
rect -10132 26746 -10130 26747
rect -10298 26719 -10282 26735
rect -10320 26693 -10314 26699
rect -10222 26697 -10213 26737
rect -10160 26697 -10149 26737
rect -10131 26697 -10130 26746
rect -10077 26737 -10071 26755
rect -10065 26747 -10057 26759
rect -10020 26755 -10013 26776
rect -10054 26751 -10030 26755
rect -10023 26751 -10012 26755
rect -10054 26747 -10041 26751
rect -10065 26745 -10055 26747
rect -10050 26745 -10044 26747
rect -10020 26745 -10013 26751
rect -10002 26745 -9995 26747
rect -10061 26742 -10050 26745
rect -10043 26742 -10036 26745
rect -10061 26737 -10052 26742
rect -10031 26737 -10022 26745
rect -10003 26737 -9995 26745
rect -9989 26737 -9985 26751
rect -10084 26697 -10081 26737
rect -10079 26697 -10072 26737
rect -10068 26697 -10064 26737
rect -10061 26697 -10054 26737
rect -10049 26697 -10042 26737
rect -10038 26697 -10033 26737
rect -10030 26697 -10023 26737
rect -10021 26697 -10012 26737
rect -10011 26697 -10005 26737
rect -10003 26697 -9996 26737
rect -10324 26689 -10320 26693
rect -10258 26685 -10252 26695
rect -10222 26689 -10215 26697
rect -10084 26689 -10064 26697
rect -10050 26689 -10043 26697
rect -10021 26689 -10013 26697
rect -9992 26689 -9985 26737
rect -9968 26689 -9966 26747
rect -10486 26677 -10478 26685
rect -10248 26677 -10242 26685
rect -10018 26677 -10015 26689
rect -10486 26669 -10370 26677
rect -10248 26669 -10241 26677
rect -10225 26669 -10207 26677
rect -10191 26669 -10176 26677
rect -10018 26669 -10011 26677
rect -9995 26669 -9968 26677
rect -9952 26669 -9949 26677
rect -9914 26667 -9909 26826
rect -9892 26793 -9886 26833
rect -9892 26667 -9888 26793
rect -10822 26650 -10810 26658
rect -10794 26650 -10782 26658
rect -10762 26650 -10754 26658
rect -10734 26650 -10718 26658
rect -10702 26650 -10690 26658
rect -10674 26650 -10662 26658
rect -10642 26650 -10634 26658
rect -10578 26650 -10570 26658
rect -10550 26650 -10542 26658
rect -10518 26650 -10510 26658
rect -10490 26650 -10482 26658
rect -10462 26650 -10454 26658
rect -10434 26650 -10426 26658
rect -10423 26656 -10410 26658
rect -10406 26650 -10398 26658
rect -10378 26650 -10370 26658
rect -10365 26656 -10354 26658
rect -10350 26650 -10342 26658
rect -10322 26650 -10314 26658
rect -10294 26650 -10286 26658
rect -10266 26650 -10258 26658
rect -10238 26650 -10230 26658
rect -10210 26656 -10192 26658
rect -10210 26650 -10202 26656
rect -10154 26650 -10148 26661
rect -10126 26650 -10120 26661
rect -10084 26653 -10076 26661
rect -10072 26653 -10064 26661
rect -10056 26653 -10048 26661
rect -10044 26653 -10036 26661
rect -10028 26653 -10020 26661
rect -10016 26653 -10008 26661
rect -10000 26653 -9992 26661
rect -9988 26653 -9972 26658
rect -9956 26653 -9944 26658
rect -9928 26653 -9916 26658
rect -10072 26652 -10056 26653
rect -10044 26652 -10028 26653
rect -10016 26652 -10000 26653
rect -9988 26652 -9980 26653
rect -11068 26642 -11058 26650
rect -11040 26642 -11030 26650
rect -11028 26639 -11026 26650
rect -10990 26642 -10982 26650
rect -10942 26642 -10938 26650
rect -10932 26639 -10930 26650
rect -10914 26642 -10910 26650
rect -10870 26642 -10862 26650
rect -10838 26642 -10834 26650
rect -10810 26642 -10806 26650
rect -10836 26639 -10834 26642
rect -10788 26639 -10786 26650
rect -10782 26642 -10778 26650
rect -10754 26642 -10746 26650
rect -10706 26642 -10702 26650
rect -10678 26642 -10674 26650
rect -10668 26639 -10666 26650
rect -10634 26642 -10626 26650
rect -10586 26642 -10578 26650
rect -10558 26642 -10550 26650
rect -10510 26642 -10502 26650
rect -10482 26642 -10474 26650
rect -10454 26642 -10446 26650
rect -10426 26642 -10418 26650
rect -10398 26642 -10390 26650
rect -10370 26642 -10362 26650
rect -10342 26642 -10334 26650
rect -10314 26642 -10306 26650
rect -10286 26642 -10278 26650
rect -10258 26642 -10250 26650
rect -10230 26642 -10222 26650
rect -10202 26642 -10194 26650
rect -10148 26645 -10138 26650
rect -10120 26645 -10110 26650
rect -10064 26645 -10056 26652
rect -10036 26645 -10028 26652
rect -10008 26645 -10000 26652
rect -9960 26642 -9956 26653
rect -9932 26642 -9928 26653
rect -10512 26639 -10476 26642
rect -10126 26639 -10092 26641
rect -9876 26639 -9874 26893
rect -9828 26658 -9826 26979
rect -9733 26972 -9730 26979
rect -9732 26956 -9730 26972
rect -9708 26966 -9706 26979
rect -9612 26969 -9610 26979
rect -9797 26916 -9785 26956
rect -9735 26908 -9730 26956
rect -9719 26953 -9716 26963
rect -9710 26953 -9709 26956
rect -9708 26953 -9699 26966
rect -9612 26955 -9608 26969
rect -9607 26955 -9600 26967
rect -9710 26937 -9706 26953
rect -9710 26908 -9709 26937
rect -9732 26849 -9730 26908
rect -9733 26791 -9729 26849
rect -9732 26658 -9730 26791
rect -9708 26658 -9706 26937
rect -9612 26945 -9600 26955
rect -9693 26895 -9691 26899
rect -9701 26791 -9699 26889
rect -9683 26881 -9681 26895
rect -9679 26791 -9675 26849
rect -9662 26831 -9658 26839
rect -9674 26791 -9663 26831
rect -9661 26791 -9658 26831
rect -9679 26783 -9676 26791
rect -9652 26667 -9648 26791
rect -9612 26658 -9610 26945
rect -9608 26929 -9600 26945
rect -9607 26919 -9600 26929
rect -9516 26921 -9514 26979
rect -9513 26969 -9512 26979
rect -9513 26921 -9506 26969
rect -9493 26961 -9479 26969
rect -9516 26915 -9506 26921
rect -9581 26667 -9572 26841
rect -9516 26658 -9514 26915
rect -9505 26911 -9502 26915
rect -9494 26911 -9489 26959
rect -9495 26841 -9489 26851
rect -9479 26841 -9476 26851
rect -9468 26841 -9466 26979
rect -9420 26917 -9417 26979
rect -9400 26972 -9391 26979
rect -9396 26969 -9392 26972
rect -9396 26953 -9393 26969
rect -9433 26907 -9428 26913
rect -9433 26903 -9426 26907
rect -9420 26903 -9416 26917
rect -9423 26893 -9416 26903
rect -9423 26889 -9418 26893
rect -9420 26843 -9418 26889
rect -9403 26849 -9399 26889
rect -9396 26849 -9394 26953
rect -9485 26793 -9479 26841
rect -9469 26793 -9466 26841
rect -9448 26833 -9442 26841
rect -9468 26658 -9466 26793
rect -9436 26793 -9430 26833
rect -9436 26667 -9432 26793
rect -9420 26791 -9410 26843
rect -9403 26839 -9393 26849
rect -9391 26839 -9384 26972
rect -9383 26953 -9380 26963
rect -9372 26953 -9370 26979
rect -9373 26937 -9370 26953
rect -9396 26833 -9394 26839
rect -9409 26791 -9403 26833
rect -9862 26650 -9852 26658
rect -9834 26650 -9824 26658
rect -9802 26650 -9794 26658
rect -9774 26650 -9758 26658
rect -9742 26650 -9730 26658
rect -9714 26650 -9702 26658
rect -9682 26650 -9674 26658
rect -9618 26650 -9610 26658
rect -9590 26650 -9582 26658
rect -9558 26650 -9550 26658
rect -9530 26650 -9514 26658
rect -9500 26650 -9488 26658
rect -9472 26650 -9460 26658
rect -9868 26642 -9862 26650
rect -9840 26642 -9834 26650
rect -9828 26639 -9826 26650
rect -9794 26642 -9786 26650
rect -9746 26642 -9742 26650
rect -9732 26639 -9730 26650
rect -9718 26642 -9714 26650
rect -9708 26639 -9706 26650
rect -9674 26642 -9666 26650
rect -9626 26642 -9618 26650
rect -9612 26639 -9610 26650
rect -9598 26642 -9590 26650
rect -9550 26642 -9542 26650
rect -9516 26639 -9514 26650
rect -9502 26642 -9500 26650
rect -9488 26642 -9486 26650
rect -9474 26642 -9472 26650
rect -9468 26639 -9466 26650
rect -9460 26642 -9458 26650
rect -9420 26639 -9418 26791
rect -9401 26785 -9394 26833
rect -9392 26785 -9383 26839
rect -9372 26833 -9370 26937
rect -9357 26895 -9355 26899
rect -9347 26881 -9345 26895
rect -9382 26791 -9376 26833
rect -9374 26785 -9367 26833
rect -9365 26791 -9356 26843
rect -9343 26791 -9339 26849
rect -9326 26831 -9322 26839
rect -9338 26791 -9327 26831
rect -9325 26791 -9322 26831
rect -9396 26658 -9394 26785
rect -9391 26783 -9384 26785
rect -9372 26658 -9370 26785
rect -9343 26783 -9340 26791
rect -9316 26667 -9312 26791
rect -9406 26650 -9394 26658
rect -9378 26650 -9368 26658
rect -9346 26650 -9338 26658
rect -9318 26650 -9302 26658
rect -9412 26642 -9406 26650
rect -9396 26639 -9394 26650
rect -9384 26642 -9378 26650
rect -9372 26639 -9370 26650
rect -9338 26642 -9330 26650
rect -9300 26639 -9298 26979
rect -9274 26977 -9272 26979
rect -9297 26959 -9291 26964
rect -9297 26945 -9282 26959
rect -9297 26929 -9281 26945
rect -9297 26916 -9291 26929
rect -9271 26916 -9269 26964
rect -9252 26658 -9250 26979
rect -9158 26977 -9151 26979
rect -9158 26966 -9149 26977
rect -9158 26961 -9141 26966
rect -9221 26916 -9209 26956
rect -9158 26900 -9151 26961
rect -9136 26908 -9133 26956
rect -9156 26851 -9154 26900
rect -9157 26667 -9150 26851
rect -9143 26841 -9140 26851
rect -9132 26841 -9130 26979
rect -9094 26915 -9091 26925
rect -9084 26917 -9082 26979
rect -9071 26977 -9066 26979
rect -9062 26953 -9055 26979
rect -9084 26893 -9080 26917
rect -9133 26793 -9130 26841
rect -9112 26833 -9106 26841
rect -9156 26658 -9154 26667
rect -9132 26658 -9130 26793
rect -9100 26793 -9094 26833
rect -9100 26667 -9096 26793
rect -9286 26650 -9274 26658
rect -9258 26650 -9246 26658
rect -9226 26650 -9218 26658
rect -9164 26650 -9154 26658
rect -9136 26650 -9126 26658
rect -9290 26642 -9286 26650
rect -9262 26642 -9258 26650
rect -9252 26639 -9250 26650
rect -9218 26642 -9210 26650
rect -9170 26642 -9164 26650
rect -9156 26639 -9154 26650
rect -9142 26642 -9136 26650
rect -9132 26639 -9130 26650
rect -9084 26639 -9082 26893
rect -9080 26667 -9074 26841
rect -9060 26833 -9058 26953
rect -9047 26841 -9044 26851
rect -9036 26841 -9034 26979
rect -8991 26917 -8985 26979
rect -8972 26969 -8969 26979
rect -8964 26969 -8960 26979
rect -8964 26953 -8961 26969
rect -9001 26907 -8996 26913
rect -9001 26903 -8994 26907
rect -8991 26893 -8984 26917
rect -8991 26889 -8986 26893
rect -8988 26841 -8986 26889
rect -8972 26891 -8969 26953
rect -8972 26889 -8967 26891
rect -8972 26851 -8969 26889
rect -8964 26851 -8962 26953
rect -8975 26841 -8962 26851
rect -9055 26833 -9047 26841
rect -9037 26833 -9034 26841
rect -9073 26793 -9064 26833
rect -9062 26793 -9057 26833
rect -9053 26793 -9047 26833
rect -9046 26793 -9030 26833
rect -9062 26785 -9055 26793
rect -9036 26785 -9030 26793
rect -9060 26658 -9058 26785
rect -9036 26658 -9034 26785
rect -9026 26667 -9020 26841
rect -9016 26833 -9010 26841
rect -8988 26833 -8979 26841
rect -8971 26833 -8962 26841
rect -8959 26841 -8955 26979
rect -8945 26841 -8942 26979
rect -9004 26793 -8998 26833
rect -8990 26793 -8979 26833
rect -8977 26793 -8974 26833
rect -8972 26793 -8961 26833
rect -8959 26793 -8952 26841
rect -8940 26833 -8938 26979
rect -8896 26978 -8890 26979
rect -8903 26841 -8900 26851
rect -8892 26841 -8890 26978
rect -8856 26956 -8852 26966
rect -8844 26956 -8842 26979
rect -8846 26942 -8842 26956
rect -8924 26833 -8920 26841
rect -8896 26833 -8890 26841
rect -8870 26833 -8866 26841
rect -8844 26837 -8842 26942
rect -8815 26932 -8808 26979
rect -8807 26955 -8804 26965
rect -8796 26955 -8794 26979
rect -8797 26939 -8794 26955
rect -8756 26948 -8747 26979
rect -8700 26971 -8698 26979
rect -8680 26977 -8676 26979
rect -8700 26957 -8696 26971
rect -8680 26967 -8670 26977
rect -8695 26957 -8688 26967
rect -8700 26947 -8688 26957
rect -8833 26847 -8824 26883
rect -8833 26837 -8823 26847
rect -8815 26837 -8808 26916
rect -8854 26833 -8835 26837
rect -8950 26793 -8947 26833
rect -9004 26667 -9000 26793
rect -9068 26650 -9058 26658
rect -9040 26650 -9032 26658
rect -9008 26650 -8992 26658
rect -9076 26642 -9068 26650
rect -9060 26639 -9058 26650
rect -9048 26642 -9040 26650
rect -9036 26639 -9034 26650
rect -8988 26639 -8986 26793
rect -8972 26785 -8965 26793
rect -8964 26658 -8962 26793
rect -8945 26785 -8938 26833
rect -8936 26793 -8934 26833
rect -8940 26658 -8938 26785
rect -8914 26667 -8910 26833
rect -8909 26793 -8898 26833
rect -8896 26793 -8889 26833
rect -8887 26793 -8884 26833
rect -8882 26793 -8871 26833
rect -8869 26793 -8866 26833
rect -8844 26827 -8835 26833
rect -8976 26650 -8962 26658
rect -8948 26650 -8936 26658
rect -8916 26650 -8908 26658
rect -8980 26642 -8976 26650
rect -8964 26639 -8962 26650
rect -8952 26642 -8948 26650
rect -8940 26639 -8938 26650
rect -8908 26642 -8900 26650
rect -8892 26639 -8890 26793
rect -8889 26785 -8884 26793
rect -8860 26667 -8856 26793
rect -8844 26789 -8834 26827
rect -8833 26789 -8827 26833
rect -8888 26650 -8880 26658
rect -8880 26642 -8872 26650
rect -8844 26639 -8842 26789
rect -8825 26785 -8818 26833
rect -8816 26785 -8807 26837
rect -8796 26833 -8794 26939
rect -8770 26934 -8768 26939
rect -8758 26934 -8756 26939
rect -8756 26929 -8748 26934
rect -8746 26924 -8738 26929
rect -8749 26883 -8743 26909
rect -8806 26789 -8800 26833
rect -8798 26785 -8791 26833
rect -8789 26789 -8780 26843
rect -8768 26819 -8763 26847
rect -8750 26829 -8746 26837
rect -8767 26789 -8763 26819
rect -8762 26789 -8751 26829
rect -8749 26789 -8746 26829
rect -8815 26781 -8808 26785
rect -8796 26658 -8794 26785
rect -8767 26781 -8764 26789
rect -8740 26667 -8736 26789
rect -8700 26658 -8698 26947
rect -8696 26931 -8688 26947
rect -8695 26919 -8688 26931
rect -8669 26911 -8660 26967
rect -8604 26921 -8602 26979
rect -8601 26969 -8600 26979
rect -8601 26921 -8594 26969
rect -8581 26961 -8567 26969
rect -8604 26915 -8594 26921
rect -8669 26861 -8667 26901
rect -8669 26667 -8660 26839
rect -8604 26658 -8602 26915
rect -8593 26911 -8590 26915
rect -8582 26911 -8577 26959
rect -8583 26841 -8577 26851
rect -8567 26841 -8564 26851
rect -8556 26841 -8554 26979
rect -8518 26915 -8515 26925
rect -8508 26917 -8506 26979
rect -8495 26977 -8490 26979
rect -8486 26953 -8479 26979
rect -8508 26893 -8504 26917
rect -8573 26793 -8567 26841
rect -8557 26793 -8554 26841
rect -8536 26833 -8530 26841
rect -8556 26658 -8554 26793
rect -8524 26793 -8518 26833
rect -8524 26667 -8520 26793
rect -8826 26650 -8816 26658
rect -8798 26650 -8788 26658
rect -8766 26650 -8758 26658
rect -8738 26650 -8722 26658
rect -8706 26650 -8694 26658
rect -8678 26650 -8666 26658
rect -8646 26650 -8638 26658
rect -8618 26650 -8602 26658
rect -8588 26650 -8576 26658
rect -8560 26650 -8548 26658
rect -8832 26642 -8826 26650
rect -8804 26642 -8798 26650
rect -8796 26639 -8794 26650
rect -8758 26642 -8750 26650
rect -8710 26642 -8706 26650
rect -8700 26639 -8698 26650
rect -8682 26642 -8678 26650
rect -8638 26642 -8630 26650
rect -8604 26639 -8602 26650
rect -8590 26642 -8588 26650
rect -8576 26642 -8574 26650
rect -8562 26642 -8560 26650
rect -8556 26639 -8554 26650
rect -8548 26642 -8546 26650
rect -8508 26639 -8506 26893
rect -8504 26667 -8498 26841
rect -8484 26833 -8482 26953
rect -8471 26841 -8468 26851
rect -8460 26841 -8458 26979
rect -8422 26915 -8419 26925
rect -8412 26917 -8410 26979
rect -8399 26977 -8394 26979
rect -8390 26953 -8383 26979
rect -8412 26893 -8408 26917
rect -8479 26833 -8471 26841
rect -8461 26833 -8458 26841
rect -8497 26793 -8488 26833
rect -8486 26793 -8481 26833
rect -8477 26793 -8471 26833
rect -8470 26793 -8454 26833
rect -8486 26785 -8479 26793
rect -8460 26785 -8454 26793
rect -8484 26658 -8482 26785
rect -8460 26658 -8458 26785
rect -8450 26667 -8444 26841
rect -8440 26833 -8434 26841
rect -8428 26793 -8422 26833
rect -8428 26667 -8424 26793
rect -8492 26650 -8482 26658
rect -8464 26650 -8456 26658
rect -8500 26642 -8492 26650
rect -8484 26639 -8482 26650
rect -8472 26642 -8464 26650
rect -8460 26639 -8458 26650
rect -8412 26639 -8410 26893
rect -8408 26667 -8402 26841
rect -8388 26833 -8386 26953
rect -8375 26841 -8372 26851
rect -8364 26841 -8362 26979
rect -8326 26915 -8323 26925
rect -8316 26917 -8314 26979
rect -8303 26977 -8298 26979
rect -8294 26953 -8287 26979
rect -8316 26893 -8312 26917
rect -8383 26833 -8375 26841
rect -8365 26833 -8362 26841
rect -8401 26793 -8392 26833
rect -8390 26793 -8385 26833
rect -8381 26793 -8375 26833
rect -8374 26793 -8358 26833
rect -8390 26785 -8383 26793
rect -8364 26785 -8358 26793
rect -8388 26658 -8386 26785
rect -8364 26658 -8362 26785
rect -8354 26667 -8348 26841
rect -8344 26833 -8338 26841
rect -8332 26793 -8326 26833
rect -8332 26667 -8328 26793
rect -8396 26650 -8386 26658
rect -8368 26650 -8360 26658
rect -8404 26642 -8396 26650
rect -8388 26639 -8386 26650
rect -8376 26642 -8368 26650
rect -8364 26639 -8362 26650
rect -8316 26639 -8314 26893
rect -8312 26667 -8306 26841
rect -8292 26833 -8290 26953
rect -8279 26841 -8276 26851
rect -8268 26841 -8266 26979
rect -8196 26969 -8191 26979
rect -8196 26953 -8193 26969
rect -8192 26967 -8191 26969
rect -8192 26953 -8184 26967
rect -8287 26833 -8279 26841
rect -8269 26833 -8266 26841
rect -8305 26793 -8296 26833
rect -8294 26793 -8289 26833
rect -8285 26793 -8279 26833
rect -8278 26793 -8262 26833
rect -8294 26785 -8287 26793
rect -8268 26785 -8262 26793
rect -8292 26658 -8290 26785
rect -8268 26658 -8266 26785
rect -8258 26667 -8252 26841
rect -8248 26833 -8242 26841
rect -8236 26793 -8230 26833
rect -8236 26667 -8232 26793
rect -8196 26658 -8194 26953
rect -8191 26919 -8184 26953
rect -8165 26667 -8156 26843
rect -8300 26650 -8290 26658
rect -8272 26650 -8264 26658
rect -8202 26650 -8194 26658
rect -8174 26650 -8168 26658
rect -8142 26650 -8134 26658
rect -8114 26650 -8102 26658
rect -8100 26650 -8098 26979
rect -8092 26964 -8090 26969
rect -8097 26916 -8090 26964
rect -8089 26916 -8073 26959
rect -8074 26911 -8073 26916
rect -8052 26658 -8050 26979
rect -7932 26966 -7930 26979
rect -8021 26916 -8009 26956
rect -7959 26932 -7954 26956
rect -7943 26955 -7940 26965
rect -7934 26955 -7933 26956
rect -7932 26955 -7923 26966
rect -7934 26939 -7930 26955
rect -7892 26948 -7883 26979
rect -7836 26971 -7834 26979
rect -7816 26977 -7812 26979
rect -7836 26957 -7832 26971
rect -7816 26967 -7806 26977
rect -7831 26957 -7824 26967
rect -7836 26947 -7824 26957
rect -7960 26916 -7944 26932
rect -7959 26908 -7954 26916
rect -7934 26908 -7933 26939
rect -7957 26789 -7953 26847
rect -7932 26658 -7930 26939
rect -7906 26934 -7904 26939
rect -7894 26934 -7892 26939
rect -7892 26929 -7884 26934
rect -7882 26924 -7874 26929
rect -7925 26789 -7923 26919
rect -7885 26883 -7879 26909
rect -7904 26819 -7899 26847
rect -7886 26829 -7882 26837
rect -7903 26789 -7899 26819
rect -7898 26789 -7887 26829
rect -7885 26789 -7882 26829
rect -7903 26781 -7900 26789
rect -7876 26667 -7872 26789
rect -7836 26658 -7834 26947
rect -7832 26931 -7824 26947
rect -7831 26919 -7824 26931
rect -7805 26911 -7796 26967
rect -7740 26921 -7738 26979
rect -7737 26969 -7736 26979
rect -7737 26921 -7730 26969
rect -7717 26961 -7703 26969
rect -7740 26915 -7730 26921
rect -7805 26861 -7803 26901
rect -7805 26667 -7796 26839
rect -7740 26658 -7738 26915
rect -7729 26911 -7726 26915
rect -7718 26911 -7713 26959
rect -7719 26841 -7713 26851
rect -7703 26841 -7700 26851
rect -7692 26841 -7690 26979
rect -7620 26969 -7615 26979
rect -7620 26953 -7617 26969
rect -7616 26967 -7615 26969
rect -7496 26967 -7487 26969
rect -7616 26953 -7608 26967
rect -7709 26793 -7703 26841
rect -7693 26793 -7690 26841
rect -7672 26833 -7666 26841
rect -7692 26658 -7690 26793
rect -7660 26793 -7654 26833
rect -7660 26667 -7656 26793
rect -7620 26658 -7618 26953
rect -7615 26919 -7608 26953
rect -7496 26919 -7485 26967
rect -7396 26911 -7394 26969
rect -7380 26933 -7377 26959
rect -7389 26919 -7377 26933
rect -7380 26911 -7377 26919
rect -7367 26900 -7364 26910
rect -7356 26900 -7354 26979
rect -7310 26911 -7298 26914
rect -7357 26886 -7354 26900
rect -7304 26888 -7298 26911
rect -7589 26667 -7580 26843
rect -7386 26771 -7377 26781
rect -7376 26755 -7367 26771
rect -7378 26745 -7377 26755
rect -7368 26667 -7367 26745
rect -8086 26650 -8074 26658
rect -8058 26650 -8046 26658
rect -8026 26650 -8018 26658
rect -7962 26650 -7954 26658
rect -7934 26650 -7926 26658
rect -7902 26650 -7894 26658
rect -7874 26650 -7858 26658
rect -7842 26650 -7830 26658
rect -7814 26650 -7802 26658
rect -7782 26650 -7774 26658
rect -7754 26650 -7738 26658
rect -7724 26650 -7712 26658
rect -7696 26650 -7684 26658
rect -7626 26650 -7618 26658
rect -7598 26650 -7592 26658
rect -7566 26650 -7558 26658
rect -7538 26650 -7522 26658
rect -7506 26650 -7494 26658
rect -7478 26650 -7466 26658
rect -7446 26650 -7438 26658
rect -7390 26650 -7389 26661
rect -7362 26650 -7361 26661
rect -7356 26650 -7354 26886
rect -7314 26805 -7310 26815
rect -7295 26805 -7288 26979
rect -7284 26919 -7282 26979
rect -7265 26919 -7258 26979
rect -7284 26908 -7270 26919
rect -7284 26904 -7266 26908
rect -7284 26892 -7278 26904
rect -7270 26903 -7266 26904
rect -7258 26903 -7254 26906
rect -7246 26903 -7244 26929
rect -7212 26905 -7210 26979
rect -7188 26920 -7186 26979
rect -7198 26910 -7194 26915
rect -7208 26905 -7198 26910
rect -7304 26789 -7300 26805
rect -7295 26763 -7288 26789
rect -7284 26755 -7282 26892
rect -7265 26824 -7258 26903
rect -7212 26901 -7198 26905
rect -7212 26881 -7208 26901
rect -7188 26896 -7184 26920
rect -7116 26917 -7113 26979
rect -7096 26972 -7087 26979
rect -7092 26969 -7088 26972
rect -7092 26953 -7089 26969
rect -7129 26907 -7124 26913
rect -7129 26903 -7122 26907
rect -7116 26903 -7112 26917
rect -7273 26776 -7266 26824
rect -7246 26776 -7240 26824
rect -7333 26737 -7324 26745
rect -7320 26737 -7314 26755
rect -7293 26751 -7273 26755
rect -7293 26748 -7282 26751
rect -7297 26747 -7282 26748
rect -7302 26745 -7300 26747
rect -7295 26745 -7288 26747
rect -7284 26745 -7282 26747
rect -7265 26745 -7258 26776
rect -7304 26742 -7295 26745
rect -7288 26742 -7279 26745
rect -7323 26697 -7314 26737
rect -7313 26697 -7307 26737
rect -7304 26697 -7297 26742
rect -7284 26737 -7282 26742
rect -7274 26737 -7266 26745
rect -7247 26737 -7240 26747
rect -7234 26745 -7230 26751
rect -7292 26697 -7288 26737
rect -7323 26689 -7307 26697
rect -7295 26689 -7288 26697
rect -7284 26697 -7276 26737
rect -7273 26697 -7267 26737
rect -7284 26661 -7282 26697
rect -7265 26689 -7258 26737
rect -7256 26697 -7248 26737
rect -7246 26697 -7240 26737
rect -7237 26689 -7230 26697
rect -7261 26677 -7260 26689
rect -7212 26677 -7210 26881
rect -7208 26816 -7207 26841
rect -7190 26816 -7189 26818
rect -7188 26816 -7186 26896
rect -7175 26895 -7168 26901
rect -7119 26893 -7112 26903
rect -7119 26889 -7114 26893
rect -7116 26843 -7114 26889
rect -7099 26849 -7095 26889
rect -7092 26849 -7090 26953
rect -7183 26816 -7182 26841
rect -7144 26833 -7138 26841
rect -7208 26793 -7192 26816
rect -7190 26793 -7183 26816
rect -7181 26793 -7165 26816
rect -7163 26793 -7162 26818
rect -7132 26793 -7126 26833
rect -7190 26785 -7189 26793
rect -7261 26669 -7256 26677
rect -7240 26669 -7208 26677
rect -7325 26653 -7316 26661
rect -7313 26653 -7304 26661
rect -7297 26653 -7288 26661
rect -7285 26653 -7276 26661
rect -7268 26653 -7260 26661
rect -7256 26653 -7248 26661
rect -7240 26653 -7232 26661
rect -7212 26658 -7210 26669
rect -7188 26658 -7186 26793
rect -7168 26780 -7164 26793
rect -7132 26667 -7128 26793
rect -7116 26791 -7106 26843
rect -7099 26839 -7089 26849
rect -7087 26839 -7080 26972
rect -7079 26953 -7076 26963
rect -7068 26953 -7066 26979
rect -7069 26937 -7066 26953
rect -7092 26833 -7090 26839
rect -7105 26791 -7099 26833
rect -7228 26653 -7210 26658
rect -7196 26653 -7184 26658
rect -7168 26653 -7156 26658
rect -7313 26652 -7297 26653
rect -7285 26652 -7269 26653
rect -7256 26652 -7240 26653
rect -7228 26652 -7220 26653
rect -8308 26642 -8300 26650
rect -8292 26639 -8290 26650
rect -8280 26642 -8272 26650
rect -8268 26639 -8266 26650
rect -8212 26642 -8202 26650
rect -8196 26639 -8194 26650
rect -8184 26642 -8174 26650
rect -8134 26642 -8126 26650
rect -8102 26642 -8098 26650
rect -8074 26642 -8070 26650
rect -8100 26639 -8098 26642
rect -8052 26639 -8050 26650
rect -8046 26642 -8042 26650
rect -8018 26642 -8010 26650
rect -7970 26642 -7962 26650
rect -7942 26642 -7934 26650
rect -7932 26639 -7930 26650
rect -7894 26642 -7886 26650
rect -7846 26642 -7842 26650
rect -7836 26639 -7834 26650
rect -7818 26642 -7814 26650
rect -7774 26642 -7766 26650
rect -7740 26639 -7738 26650
rect -7726 26642 -7724 26650
rect -7712 26642 -7710 26650
rect -7698 26642 -7696 26650
rect -7692 26639 -7690 26650
rect -7684 26642 -7682 26650
rect -7636 26642 -7626 26650
rect -7620 26639 -7618 26650
rect -7608 26642 -7598 26650
rect -7558 26642 -7550 26650
rect -7510 26642 -7506 26650
rect -7482 26642 -7478 26650
rect -7438 26642 -7430 26650
rect -7389 26645 -7374 26650
rect -7361 26645 -7346 26650
rect -7304 26645 -7297 26652
rect -7356 26639 -7354 26645
rect -7284 26639 -7282 26652
rect -7276 26645 -7269 26652
rect -7248 26645 -7240 26652
rect -7212 26639 -7210 26653
rect -7200 26642 -7196 26653
rect -7188 26639 -7186 26653
rect -7172 26642 -7168 26653
rect -7116 26639 -7114 26791
rect -7097 26785 -7090 26833
rect -7088 26785 -7079 26839
rect -7068 26833 -7066 26937
rect -7053 26895 -7051 26899
rect -7043 26881 -7041 26895
rect -7078 26791 -7072 26833
rect -7070 26785 -7063 26833
rect -7061 26791 -7052 26843
rect -7039 26791 -7035 26849
rect -7022 26831 -7018 26839
rect -7034 26791 -7023 26831
rect -7021 26791 -7018 26831
rect -7092 26658 -7090 26785
rect -7087 26783 -7080 26785
rect -7068 26658 -7066 26785
rect -7039 26783 -7036 26791
rect -7012 26667 -7008 26791
rect -7102 26650 -7090 26658
rect -7074 26650 -7064 26658
rect -7042 26650 -7034 26658
rect -7108 26642 -7102 26650
rect -7092 26639 -7090 26650
rect -7080 26642 -7074 26650
rect -7068 26639 -7066 26650
rect -7034 26642 -7026 26650
rect -6996 26639 -6994 26979
rect -6972 26977 -6958 26979
rect -6972 26969 -6970 26977
rect -6973 26961 -6968 26969
rect -6972 26955 -6968 26961
rect -6974 26929 -6967 26955
rect -6992 26667 -6986 26841
rect -6972 26831 -6970 26929
rect -6959 26841 -6956 26851
rect -6948 26841 -6946 26979
rect -6910 26915 -6907 26925
rect -6900 26917 -6898 26979
rect -6887 26977 -6882 26979
rect -6878 26953 -6871 26979
rect -6900 26893 -6896 26917
rect -6967 26831 -6959 26841
rect -6949 26831 -6946 26841
rect -6985 26793 -6976 26831
rect -6974 26793 -6969 26831
rect -6965 26793 -6959 26831
rect -6958 26793 -6942 26831
rect -6974 26785 -6967 26793
rect -6948 26785 -6942 26793
rect -6972 26658 -6970 26785
rect -6948 26658 -6946 26785
rect -6938 26667 -6932 26841
rect -6928 26833 -6922 26841
rect -6916 26793 -6910 26833
rect -6916 26667 -6912 26793
rect -6980 26650 -6970 26658
rect -6952 26650 -6942 26658
rect -6986 26642 -6980 26650
rect -6972 26639 -6970 26650
rect -6958 26642 -6952 26650
rect -6948 26639 -6946 26650
rect -6900 26639 -6898 26893
rect -6896 26667 -6890 26841
rect -6876 26833 -6874 26953
rect -6863 26841 -6860 26851
rect -6852 26841 -6850 26979
rect -6814 26915 -6811 26925
rect -6804 26917 -6802 26979
rect -6791 26977 -6786 26979
rect -6782 26953 -6775 26979
rect -6804 26893 -6800 26917
rect -6871 26833 -6863 26841
rect -6853 26833 -6850 26841
rect -6889 26793 -6880 26833
rect -6878 26793 -6873 26833
rect -6869 26793 -6863 26833
rect -6862 26793 -6846 26833
rect -6878 26785 -6871 26793
rect -6852 26785 -6846 26793
rect -6876 26658 -6874 26785
rect -6852 26658 -6850 26785
rect -6842 26667 -6836 26841
rect -6832 26833 -6826 26841
rect -6820 26793 -6814 26833
rect -6820 26667 -6816 26793
rect -6884 26650 -6874 26658
rect -6856 26650 -6848 26658
rect -6892 26642 -6884 26650
rect -6876 26639 -6874 26650
rect -6864 26642 -6856 26650
rect -6852 26639 -6850 26650
rect -6804 26639 -6802 26893
rect -6800 26667 -6794 26841
rect -6780 26833 -6778 26953
rect -6767 26841 -6764 26851
rect -6756 26841 -6754 26979
rect -6718 26915 -6715 26925
rect -6708 26917 -6706 26979
rect -6695 26977 -6690 26979
rect -6686 26953 -6679 26979
rect -6708 26893 -6704 26917
rect -6775 26833 -6767 26841
rect -6757 26833 -6754 26841
rect -6793 26793 -6784 26833
rect -6782 26793 -6777 26833
rect -6773 26793 -6767 26833
rect -6766 26793 -6750 26833
rect -6782 26785 -6775 26793
rect -6756 26785 -6750 26793
rect -6780 26658 -6778 26785
rect -6756 26658 -6754 26785
rect -6746 26667 -6740 26841
rect -6736 26833 -6730 26841
rect -6724 26793 -6718 26833
rect -6724 26667 -6720 26793
rect -6788 26650 -6778 26658
rect -6760 26650 -6752 26658
rect -6796 26642 -6788 26650
rect -6780 26639 -6778 26650
rect -6768 26642 -6760 26650
rect -6756 26639 -6754 26650
rect -6708 26639 -6706 26893
rect -6704 26667 -6698 26841
rect -6684 26833 -6682 26953
rect -6671 26841 -6668 26851
rect -6660 26841 -6658 26979
rect -6622 26915 -6619 26925
rect -6612 26917 -6610 26979
rect -6599 26977 -6594 26979
rect -6590 26953 -6583 26979
rect -6612 26893 -6608 26917
rect -6679 26833 -6671 26841
rect -6661 26833 -6658 26841
rect -6697 26793 -6688 26833
rect -6686 26793 -6681 26833
rect -6677 26793 -6671 26833
rect -6670 26793 -6654 26833
rect -6686 26785 -6679 26793
rect -6660 26785 -6654 26793
rect -6684 26658 -6682 26785
rect -6660 26658 -6658 26785
rect -6650 26667 -6644 26841
rect -6640 26833 -6634 26841
rect -6628 26793 -6622 26833
rect -6628 26667 -6624 26793
rect -6692 26650 -6682 26658
rect -6664 26650 -6656 26658
rect -6700 26642 -6692 26650
rect -6684 26639 -6682 26650
rect -6672 26642 -6664 26650
rect -6660 26639 -6658 26650
rect -6612 26639 -6610 26893
rect -6608 26667 -6602 26841
rect -6588 26833 -6586 26953
rect -6575 26841 -6572 26851
rect -6564 26841 -6562 26979
rect -6526 26915 -6523 26925
rect -6516 26917 -6514 26979
rect -6503 26977 -6498 26979
rect -6494 26953 -6487 26979
rect -6516 26893 -6512 26917
rect -6583 26833 -6575 26841
rect -6565 26833 -6562 26841
rect -6601 26793 -6592 26833
rect -6590 26793 -6585 26833
rect -6581 26793 -6575 26833
rect -6574 26793 -6558 26833
rect -6590 26785 -6583 26793
rect -6564 26785 -6558 26793
rect -6588 26658 -6586 26785
rect -6564 26658 -6562 26785
rect -6554 26667 -6548 26841
rect -6544 26833 -6538 26841
rect -6532 26793 -6526 26833
rect -6532 26667 -6528 26793
rect -6596 26650 -6586 26658
rect -6568 26650 -6560 26658
rect -6604 26642 -6596 26650
rect -6588 26639 -6586 26650
rect -6576 26642 -6568 26650
rect -6564 26639 -6562 26650
rect -6516 26639 -6514 26893
rect -6512 26667 -6506 26841
rect -6492 26833 -6490 26953
rect -6479 26841 -6476 26851
rect -6468 26841 -6466 26979
rect -6430 26915 -6427 26925
rect -6420 26917 -6418 26979
rect -6407 26977 -6402 26979
rect -6398 26953 -6391 26979
rect -6420 26893 -6416 26917
rect -6487 26833 -6479 26841
rect -6469 26833 -6466 26841
rect -6505 26793 -6496 26833
rect -6494 26793 -6489 26833
rect -6485 26793 -6479 26833
rect -6478 26793 -6462 26833
rect -6494 26785 -6487 26793
rect -6468 26785 -6462 26793
rect -6492 26658 -6490 26785
rect -6468 26658 -6466 26785
rect -6458 26667 -6452 26841
rect -6448 26833 -6442 26841
rect -6436 26793 -6430 26833
rect -6436 26667 -6432 26793
rect -6500 26650 -6490 26658
rect -6472 26650 -6464 26658
rect -6508 26642 -6500 26650
rect -6492 26639 -6490 26650
rect -6480 26642 -6472 26650
rect -6468 26639 -6466 26650
rect -6420 26639 -6418 26893
rect -6416 26667 -6410 26841
rect -6396 26833 -6394 26953
rect -6383 26841 -6380 26851
rect -6372 26841 -6370 26979
rect -6334 26915 -6331 26925
rect -6324 26917 -6322 26979
rect -6311 26977 -6306 26979
rect -6302 26953 -6295 26979
rect -6324 26893 -6320 26917
rect -6391 26833 -6383 26841
rect -6373 26833 -6370 26841
rect -6409 26793 -6400 26833
rect -6398 26793 -6393 26833
rect -6389 26793 -6383 26833
rect -6382 26793 -6366 26833
rect -6398 26785 -6391 26793
rect -6372 26785 -6366 26793
rect -6396 26658 -6394 26785
rect -6372 26658 -6370 26785
rect -6362 26667 -6356 26841
rect -6352 26833 -6346 26841
rect -6340 26793 -6334 26833
rect -6340 26667 -6336 26793
rect -6404 26650 -6394 26658
rect -6376 26650 -6368 26658
rect -6412 26642 -6404 26650
rect -6396 26639 -6394 26650
rect -6384 26642 -6376 26650
rect -6372 26639 -6370 26650
rect -6324 26639 -6322 26893
rect -6320 26667 -6314 26841
rect -6300 26833 -6298 26953
rect -6287 26841 -6284 26851
rect -6276 26841 -6274 26979
rect -6228 26917 -6226 26979
rect -6225 26953 -6209 26964
rect -6225 26917 -6219 26953
rect -6228 26916 -6219 26917
rect -6199 26916 -6197 26964
rect -6228 26893 -6224 26916
rect -6295 26833 -6287 26841
rect -6277 26833 -6274 26841
rect -6313 26793 -6304 26833
rect -6302 26793 -6297 26833
rect -6293 26793 -6287 26833
rect -6286 26793 -6270 26833
rect -6302 26785 -6295 26793
rect -6276 26785 -6270 26793
rect -6300 26658 -6298 26785
rect -6276 26658 -6274 26785
rect -6266 26667 -6260 26841
rect -6256 26833 -6250 26841
rect -6244 26793 -6238 26833
rect -6244 26667 -6240 26793
rect -6308 26650 -6298 26658
rect -6280 26650 -6272 26658
rect -6316 26642 -6308 26650
rect -6300 26639 -6298 26650
rect -6288 26642 -6280 26650
rect -6276 26639 -6274 26650
rect -6228 26639 -6226 26893
rect -6180 26658 -6178 26979
rect -6149 26916 -6137 26956
rect -6094 26916 -6087 26964
rect -6085 26916 -6079 26956
rect -6077 26908 -6070 26956
rect -6060 26658 -6058 26979
rect -5975 26956 -5970 26966
rect -5964 26956 -5957 26979
rect -6029 26916 -6017 26956
rect -5965 26900 -5957 26956
rect -5951 26900 -5948 26910
rect -5942 26908 -5941 26916
rect -5940 26900 -5938 26979
rect -5894 26911 -5882 26914
rect -5965 26755 -5960 26900
rect -5941 26886 -5938 26900
rect -5888 26888 -5882 26911
rect -5965 26697 -5957 26755
rect -6214 26650 -6204 26658
rect -6186 26650 -6176 26658
rect -6154 26650 -6146 26658
rect -6126 26650 -6110 26658
rect -6094 26650 -6082 26658
rect -6066 26650 -6054 26658
rect -6034 26650 -6026 26658
rect -5978 26650 -5973 26661
rect -5964 26650 -5962 26697
rect -5950 26650 -5945 26661
rect -5940 26650 -5938 26886
rect -5898 26805 -5894 26815
rect -5879 26805 -5872 26979
rect -5868 26919 -5866 26979
rect -5849 26919 -5842 26979
rect -5808 26956 -5804 26966
rect -5796 26956 -5794 26979
rect -5798 26942 -5794 26956
rect -5708 26948 -5699 26979
rect -5652 26971 -5650 26979
rect -5632 26977 -5628 26979
rect -5652 26957 -5648 26971
rect -5632 26967 -5622 26977
rect -5528 26967 -5519 26969
rect -5408 26967 -5399 26969
rect -5647 26957 -5640 26967
rect -5868 26908 -5854 26919
rect -5868 26904 -5850 26908
rect -5868 26892 -5862 26904
rect -5854 26903 -5850 26904
rect -5842 26903 -5838 26906
rect -5830 26903 -5828 26929
rect -5796 26905 -5794 26942
rect -5652 26947 -5640 26957
rect -5722 26934 -5720 26939
rect -5710 26934 -5708 26939
rect -5708 26929 -5700 26934
rect -5698 26924 -5690 26929
rect -5788 26911 -5786 26921
rect -5776 26919 -5752 26921
rect -5776 26916 -5760 26919
rect -5778 26910 -5776 26911
rect -5888 26789 -5884 26805
rect -5879 26763 -5872 26789
rect -5868 26755 -5866 26892
rect -5849 26824 -5842 26903
rect -5796 26881 -5792 26905
rect -5778 26895 -5776 26896
rect -5701 26883 -5695 26909
rect -5796 26837 -5794 26881
rect -5857 26776 -5850 26824
rect -5830 26776 -5824 26824
rect -5796 26816 -5791 26837
rect -5770 26826 -5766 26837
rect -5770 26816 -5765 26826
rect -5796 26789 -5779 26816
rect -5777 26789 -5775 26816
rect -5773 26789 -5770 26816
rect -5917 26737 -5908 26745
rect -5904 26737 -5898 26755
rect -5877 26751 -5857 26755
rect -5877 26748 -5866 26751
rect -5881 26747 -5866 26748
rect -5886 26745 -5884 26747
rect -5879 26745 -5872 26747
rect -5868 26745 -5866 26747
rect -5849 26745 -5842 26776
rect -5888 26742 -5879 26745
rect -5872 26742 -5863 26745
rect -5907 26697 -5898 26737
rect -5897 26697 -5891 26737
rect -5888 26697 -5881 26742
rect -5868 26737 -5866 26742
rect -5858 26737 -5850 26745
rect -5831 26737 -5824 26747
rect -5818 26745 -5814 26751
rect -5876 26697 -5872 26737
rect -5907 26689 -5891 26697
rect -5879 26689 -5872 26697
rect -5868 26697 -5860 26737
rect -5857 26697 -5851 26737
rect -5868 26661 -5866 26697
rect -5849 26689 -5842 26737
rect -5840 26697 -5832 26737
rect -5830 26697 -5824 26737
rect -5821 26689 -5814 26697
rect -5845 26677 -5844 26689
rect -5796 26677 -5794 26789
rect -5777 26781 -5773 26789
rect -5768 26768 -5765 26816
rect -5764 26789 -5752 26816
rect -5750 26781 -5748 26816
rect -5741 26789 -5738 26826
rect -5720 26819 -5715 26847
rect -5702 26829 -5698 26837
rect -5719 26789 -5715 26819
rect -5714 26789 -5703 26829
rect -5701 26789 -5698 26829
rect -5719 26781 -5716 26789
rect -5768 26689 -5765 26747
rect -5845 26669 -5840 26677
rect -5824 26669 -5778 26677
rect -5909 26653 -5900 26661
rect -5897 26653 -5888 26661
rect -5881 26653 -5872 26661
rect -5869 26653 -5860 26661
rect -5852 26653 -5844 26661
rect -5840 26653 -5832 26661
rect -5824 26653 -5816 26661
rect -5796 26658 -5794 26669
rect -5692 26667 -5688 26789
rect -5652 26658 -5650 26947
rect -5648 26931 -5640 26947
rect -5647 26919 -5640 26931
rect -5621 26911 -5612 26967
rect -5528 26919 -5517 26967
rect -5408 26919 -5397 26967
rect -5316 26921 -5314 26979
rect -5313 26969 -5312 26979
rect -5313 26921 -5306 26969
rect -5293 26961 -5279 26969
rect -5316 26915 -5306 26921
rect -5621 26861 -5619 26901
rect -5621 26667 -5612 26839
rect -5316 26658 -5314 26915
rect -5305 26911 -5302 26915
rect -5294 26911 -5289 26959
rect -5295 26841 -5289 26851
rect -5279 26841 -5276 26851
rect -5268 26841 -5266 26979
rect -5230 26915 -5227 26925
rect -5220 26917 -5218 26979
rect -5207 26977 -5202 26979
rect -5198 26953 -5191 26979
rect -5220 26893 -5216 26917
rect -5285 26793 -5279 26841
rect -5269 26793 -5266 26841
rect -5248 26833 -5242 26841
rect -5268 26658 -5266 26793
rect -5236 26793 -5230 26833
rect -5236 26667 -5232 26793
rect -5796 26653 -5784 26658
rect -5778 26653 -5768 26658
rect -5766 26653 -5756 26658
rect -5750 26653 -5740 26658
rect -5897 26652 -5881 26653
rect -5869 26652 -5853 26653
rect -5840 26652 -5824 26653
rect -5812 26652 -5804 26653
rect -5796 26652 -5778 26653
rect -5766 26652 -5750 26653
rect -5738 26652 -5728 26658
rect -6220 26642 -6214 26650
rect -6192 26642 -6186 26650
rect -6180 26639 -6178 26650
rect -6146 26642 -6138 26650
rect -6098 26642 -6094 26650
rect -6070 26642 -6066 26650
rect -6060 26639 -6058 26650
rect -6026 26642 -6018 26650
rect -5973 26645 -5962 26650
rect -5945 26645 -5934 26650
rect -5888 26645 -5881 26652
rect -5964 26639 -5962 26645
rect -5940 26639 -5938 26645
rect -5868 26639 -5866 26652
rect -5860 26645 -5853 26652
rect -5832 26645 -5824 26652
rect -5796 26639 -5794 26652
rect -5784 26642 -5778 26652
rect -5756 26642 -5750 26652
rect -5718 26650 -5710 26658
rect -5690 26650 -5674 26658
rect -5658 26650 -5646 26658
rect -5630 26650 -5618 26658
rect -5598 26650 -5590 26658
rect -5570 26650 -5554 26658
rect -5538 26650 -5526 26658
rect -5510 26650 -5498 26658
rect -5478 26650 -5470 26658
rect -5450 26650 -5434 26658
rect -5418 26650 -5406 26658
rect -5390 26650 -5378 26658
rect -5358 26650 -5350 26658
rect -5330 26650 -5314 26658
rect -5300 26650 -5288 26658
rect -5272 26650 -5260 26658
rect -5710 26642 -5702 26650
rect -5662 26642 -5658 26650
rect -5652 26639 -5650 26650
rect -5634 26642 -5630 26650
rect -5590 26642 -5582 26650
rect -5542 26642 -5538 26650
rect -5514 26642 -5510 26650
rect -5470 26642 -5462 26650
rect -5422 26642 -5418 26650
rect -5394 26642 -5390 26650
rect -5350 26642 -5342 26650
rect -5316 26639 -5314 26650
rect -5302 26642 -5300 26650
rect -5288 26642 -5286 26650
rect -5274 26642 -5272 26650
rect -5268 26639 -5266 26650
rect -5260 26642 -5258 26650
rect -5220 26639 -5218 26893
rect -5216 26667 -5210 26841
rect -5196 26833 -5194 26953
rect -5183 26841 -5180 26851
rect -5172 26841 -5170 26979
rect -5134 26915 -5131 26925
rect -5124 26917 -5122 26979
rect -5111 26977 -5106 26979
rect -5102 26953 -5095 26979
rect -5124 26893 -5120 26917
rect -5191 26833 -5183 26841
rect -5173 26833 -5170 26841
rect -5209 26793 -5200 26833
rect -5198 26793 -5193 26833
rect -5189 26793 -5183 26833
rect -5182 26793 -5166 26833
rect -5198 26785 -5191 26793
rect -5172 26785 -5166 26793
rect -5196 26658 -5194 26785
rect -5172 26658 -5170 26785
rect -5162 26667 -5156 26841
rect -5152 26833 -5146 26841
rect -5140 26793 -5134 26833
rect -5140 26667 -5136 26793
rect -5204 26650 -5194 26658
rect -5176 26650 -5168 26658
rect -5212 26642 -5204 26650
rect -5196 26639 -5194 26650
rect -5184 26642 -5176 26650
rect -5172 26639 -5170 26650
rect -5124 26639 -5122 26893
rect -5120 26667 -5114 26841
rect -5100 26833 -5098 26953
rect -5087 26841 -5084 26851
rect -5076 26841 -5074 26979
rect -5040 26956 -5035 26966
rect -5028 26956 -5025 26979
rect -5030 26953 -5016 26956
rect -5030 26942 -5025 26953
rect -5028 26917 -5025 26942
rect -4999 26932 -4992 26979
rect -4991 26955 -4988 26965
rect -4980 26955 -4978 26979
rect -4981 26939 -4978 26955
rect -4940 26948 -4931 26979
rect -4884 26971 -4882 26979
rect -4885 26961 -4880 26971
rect -4864 26961 -4858 26979
rect -4884 26957 -4880 26961
rect -5028 26893 -5024 26917
rect -5095 26833 -5087 26841
rect -5077 26833 -5074 26841
rect -5113 26793 -5104 26833
rect -5102 26793 -5097 26833
rect -5093 26793 -5087 26833
rect -5086 26793 -5070 26833
rect -5102 26785 -5095 26793
rect -5076 26785 -5070 26793
rect -5100 26658 -5098 26785
rect -5076 26658 -5074 26785
rect -5066 26667 -5060 26841
rect -5056 26833 -5050 26841
rect -5028 26837 -5026 26893
rect -5011 26847 -5008 26893
rect -5011 26837 -5001 26847
rect -4999 26837 -4992 26916
rect -5038 26833 -5019 26837
rect -5044 26793 -5038 26833
rect -5028 26827 -5019 26833
rect -5044 26667 -5040 26793
rect -5028 26789 -5018 26827
rect -5017 26789 -5011 26833
rect -5108 26650 -5098 26658
rect -5080 26650 -5072 26658
rect -5116 26642 -5108 26650
rect -5100 26639 -5098 26650
rect -5088 26642 -5080 26650
rect -5076 26639 -5074 26650
rect -5028 26639 -5026 26789
rect -5009 26785 -5002 26833
rect -5000 26785 -4991 26837
rect -4980 26833 -4978 26939
rect -4954 26934 -4952 26939
rect -4942 26934 -4940 26939
rect -4940 26929 -4932 26934
rect -4886 26931 -4879 26957
rect -4930 26924 -4922 26929
rect -4933 26883 -4927 26909
rect -4908 26908 -4906 26911
rect -4990 26789 -4984 26833
rect -4982 26785 -4975 26833
rect -4973 26789 -4964 26843
rect -4952 26819 -4947 26847
rect -4904 26839 -4899 26841
rect -4934 26829 -4930 26837
rect -4951 26789 -4947 26819
rect -4946 26789 -4935 26829
rect -4933 26789 -4930 26829
rect -4999 26781 -4992 26785
rect -4980 26658 -4978 26785
rect -4951 26781 -4948 26789
rect -4924 26667 -4920 26789
rect -4904 26667 -4898 26839
rect -4884 26829 -4882 26931
rect -4860 26901 -4858 26961
rect -4788 26969 -4783 26979
rect -4788 26953 -4785 26969
rect -4784 26967 -4783 26969
rect -4784 26953 -4776 26967
rect -4860 26885 -4852 26901
rect -4860 26861 -4851 26885
rect -4871 26841 -4868 26851
rect -4860 26841 -4858 26861
rect -4879 26839 -4872 26841
rect -4879 26829 -4871 26839
rect -4861 26829 -4858 26841
rect -4897 26793 -4888 26829
rect -4886 26793 -4881 26829
rect -4877 26793 -4871 26829
rect -4870 26793 -4854 26829
rect -4886 26785 -4879 26793
rect -4860 26785 -4854 26793
rect -4884 26658 -4882 26785
rect -4860 26658 -4858 26785
rect -4850 26667 -4844 26839
rect -4840 26833 -4834 26841
rect -4828 26793 -4822 26833
rect -4828 26667 -4824 26793
rect -4788 26658 -4786 26953
rect -4783 26919 -4776 26953
rect -4692 26921 -4690 26979
rect -4689 26969 -4688 26979
rect -4689 26921 -4682 26969
rect -4669 26961 -4655 26969
rect -4692 26915 -4682 26921
rect -4757 26667 -4748 26843
rect -4692 26658 -4690 26915
rect -4681 26911 -4678 26915
rect -4670 26911 -4665 26959
rect -4671 26841 -4665 26851
rect -4655 26841 -4652 26851
rect -4644 26841 -4642 26979
rect -4608 26956 -4603 26966
rect -4596 26956 -4593 26979
rect -4598 26953 -4584 26956
rect -4598 26942 -4593 26953
rect -4596 26917 -4593 26942
rect -4567 26932 -4560 26979
rect -4559 26955 -4556 26965
rect -4548 26955 -4546 26979
rect -4549 26939 -4546 26955
rect -4508 26948 -4499 26979
rect -4473 26961 -4467 26964
rect -4473 26947 -4458 26961
rect -4596 26893 -4592 26917
rect -4661 26793 -4655 26841
rect -4645 26793 -4642 26841
rect -4624 26833 -4618 26841
rect -4596 26837 -4594 26893
rect -4579 26847 -4576 26893
rect -4579 26837 -4569 26847
rect -4567 26837 -4560 26916
rect -4606 26833 -4587 26837
rect -4644 26658 -4642 26793
rect -4612 26793 -4606 26833
rect -4596 26827 -4587 26833
rect -4612 26667 -4608 26793
rect -4596 26789 -4586 26827
rect -4585 26789 -4579 26833
rect -5010 26650 -5004 26658
rect -4982 26650 -4976 26658
rect -4950 26650 -4942 26658
rect -4922 26650 -4908 26658
rect -4892 26650 -4880 26658
rect -4864 26650 -4852 26658
rect -4794 26650 -4786 26658
rect -4766 26650 -4760 26658
rect -4734 26650 -4726 26658
rect -4706 26650 -4690 26658
rect -4676 26650 -4664 26658
rect -4648 26650 -4636 26658
rect -5020 26642 -5010 26650
rect -4992 26642 -4982 26650
rect -4980 26639 -4978 26650
rect -4942 26642 -4934 26650
rect -4908 26642 -4906 26650
rect -4894 26642 -4892 26650
rect -4884 26639 -4882 26650
rect -4880 26642 -4878 26650
rect -4866 26642 -4864 26650
rect -4860 26639 -4858 26650
rect -4852 26642 -4850 26650
rect -4804 26642 -4794 26650
rect -4788 26639 -4786 26650
rect -4776 26642 -4766 26650
rect -4726 26642 -4718 26650
rect -4692 26639 -4690 26650
rect -4678 26642 -4676 26650
rect -4664 26642 -4662 26650
rect -4650 26642 -4648 26650
rect -4644 26639 -4642 26650
rect -4636 26642 -4634 26650
rect -4596 26639 -4594 26789
rect -4577 26785 -4570 26833
rect -4568 26785 -4559 26837
rect -4548 26833 -4546 26939
rect -4522 26934 -4520 26939
rect -4510 26934 -4508 26939
rect -4508 26929 -4500 26934
rect -4473 26931 -4457 26947
rect -4498 26924 -4490 26929
rect -4473 26916 -4467 26931
rect -4447 26916 -4445 26964
rect -4501 26883 -4495 26909
rect -4428 26885 -4426 26979
rect -4334 26977 -4327 26979
rect -4334 26966 -4325 26977
rect -4334 26961 -4317 26966
rect -4397 26916 -4385 26956
rect -4334 26900 -4327 26961
rect -4312 26908 -4309 26956
rect -4428 26861 -4419 26885
rect -4558 26789 -4552 26833
rect -4550 26785 -4543 26833
rect -4541 26789 -4532 26843
rect -4520 26819 -4515 26847
rect -4502 26829 -4498 26837
rect -4519 26789 -4515 26819
rect -4514 26789 -4503 26829
rect -4501 26789 -4498 26829
rect -4567 26781 -4560 26785
rect -4548 26658 -4546 26785
rect -4519 26781 -4516 26789
rect -4492 26667 -4488 26789
rect -4428 26658 -4426 26861
rect -4332 26851 -4330 26900
rect -4333 26667 -4326 26851
rect -4319 26841 -4316 26851
rect -4308 26841 -4306 26979
rect -4272 26956 -4267 26966
rect -4260 26956 -4257 26979
rect -4262 26953 -4248 26956
rect -4262 26942 -4257 26953
rect -4260 26917 -4257 26942
rect -4231 26932 -4224 26979
rect -4223 26955 -4220 26965
rect -4212 26955 -4210 26979
rect -4213 26939 -4210 26955
rect -4172 26948 -4163 26979
rect -4116 26971 -4114 26979
rect -4117 26961 -4112 26971
rect -4096 26961 -4090 26979
rect -4116 26957 -4112 26961
rect -4260 26893 -4256 26917
rect -4309 26793 -4306 26841
rect -4288 26833 -4282 26841
rect -4260 26837 -4258 26893
rect -4243 26847 -4240 26893
rect -4243 26837 -4233 26847
rect -4231 26837 -4224 26916
rect -4270 26833 -4251 26837
rect -4332 26658 -4330 26667
rect -4308 26658 -4306 26793
rect -4276 26793 -4270 26833
rect -4260 26827 -4251 26833
rect -4276 26667 -4272 26793
rect -4260 26789 -4250 26827
rect -4249 26789 -4243 26833
rect -4578 26650 -4572 26658
rect -4550 26650 -4544 26658
rect -4518 26650 -4510 26658
rect -4490 26650 -4478 26658
rect -4462 26650 -4450 26658
rect -4434 26650 -4422 26658
rect -4402 26650 -4394 26658
rect -4340 26650 -4330 26658
rect -4312 26650 -4302 26658
rect -4588 26642 -4578 26650
rect -4560 26642 -4550 26650
rect -4548 26639 -4546 26650
rect -4510 26642 -4502 26650
rect -4478 26642 -4474 26650
rect -4450 26642 -4446 26650
rect -4428 26639 -4426 26650
rect -4422 26642 -4418 26650
rect -4394 26642 -4386 26650
rect -4346 26642 -4340 26650
rect -4332 26639 -4330 26650
rect -4318 26642 -4312 26650
rect -4308 26639 -4306 26650
rect -4260 26639 -4258 26789
rect -4241 26785 -4234 26833
rect -4232 26785 -4223 26837
rect -4212 26833 -4210 26939
rect -4186 26934 -4184 26939
rect -4174 26934 -4172 26939
rect -4172 26929 -4164 26934
rect -4118 26931 -4111 26957
rect -4162 26924 -4154 26929
rect -4165 26883 -4159 26909
rect -4140 26908 -4138 26911
rect -4222 26789 -4216 26833
rect -4214 26785 -4207 26833
rect -4205 26789 -4196 26843
rect -4184 26819 -4179 26847
rect -4136 26839 -4131 26841
rect -4166 26829 -4162 26837
rect -4183 26789 -4179 26819
rect -4178 26789 -4167 26829
rect -4165 26789 -4162 26829
rect -4231 26781 -4224 26785
rect -4212 26658 -4210 26785
rect -4183 26781 -4180 26789
rect -4156 26667 -4152 26789
rect -4136 26667 -4130 26839
rect -4116 26829 -4114 26931
rect -4092 26901 -4090 26961
rect -4020 26969 -4015 26979
rect -4020 26953 -4017 26969
rect -4016 26967 -4015 26969
rect -4016 26953 -4008 26967
rect -4092 26885 -4084 26901
rect -4092 26861 -4083 26885
rect -4103 26841 -4100 26851
rect -4092 26841 -4090 26861
rect -4111 26839 -4104 26841
rect -4111 26829 -4103 26839
rect -4093 26829 -4090 26841
rect -4129 26793 -4120 26829
rect -4118 26793 -4113 26829
rect -4109 26793 -4103 26829
rect -4102 26793 -4086 26829
rect -4118 26785 -4111 26793
rect -4092 26785 -4086 26793
rect -4116 26658 -4114 26785
rect -4092 26658 -4090 26785
rect -4082 26667 -4076 26839
rect -4072 26833 -4066 26841
rect -4060 26793 -4054 26833
rect -4060 26667 -4056 26793
rect -4020 26658 -4018 26953
rect -4015 26919 -4008 26953
rect -3916 26911 -3914 26969
rect -3900 26933 -3897 26959
rect -3909 26919 -3897 26933
rect -3900 26911 -3897 26919
rect -3887 26900 -3884 26910
rect -3876 26900 -3874 26979
rect -3830 26911 -3818 26914
rect -3877 26886 -3874 26900
rect -3824 26888 -3818 26911
rect -3989 26667 -3980 26843
rect -3906 26771 -3897 26781
rect -3896 26755 -3887 26771
rect -3898 26745 -3897 26755
rect -3888 26667 -3887 26745
rect -4242 26650 -4236 26658
rect -4214 26650 -4208 26658
rect -4182 26650 -4174 26658
rect -4154 26650 -4140 26658
rect -4124 26650 -4112 26658
rect -4096 26650 -4084 26658
rect -4026 26650 -4018 26658
rect -3998 26650 -3992 26658
rect -3966 26650 -3958 26658
rect -3910 26650 -3909 26661
rect -3882 26650 -3881 26661
rect -3876 26650 -3874 26886
rect -3834 26805 -3830 26815
rect -3815 26805 -3808 26979
rect -3804 26919 -3802 26979
rect -3785 26919 -3778 26979
rect -3744 26956 -3740 26966
rect -3732 26956 -3730 26979
rect -3734 26942 -3730 26956
rect -3644 26948 -3635 26979
rect -3588 26971 -3586 26979
rect -3589 26961 -3584 26971
rect -3568 26961 -3562 26979
rect -3588 26957 -3584 26961
rect -3804 26908 -3790 26919
rect -3804 26904 -3786 26908
rect -3804 26892 -3798 26904
rect -3790 26903 -3786 26904
rect -3778 26903 -3774 26906
rect -3766 26903 -3764 26929
rect -3732 26905 -3730 26942
rect -3658 26934 -3656 26939
rect -3646 26934 -3644 26939
rect -3644 26929 -3636 26934
rect -3590 26931 -3583 26957
rect -3634 26924 -3626 26929
rect -3724 26911 -3722 26921
rect -3712 26919 -3688 26921
rect -3712 26916 -3696 26919
rect -3714 26910 -3712 26911
rect -3824 26789 -3820 26805
rect -3815 26763 -3808 26789
rect -3804 26755 -3802 26892
rect -3785 26824 -3778 26903
rect -3732 26881 -3728 26905
rect -3714 26895 -3712 26896
rect -3637 26883 -3631 26909
rect -3612 26908 -3610 26911
rect -3732 26837 -3730 26881
rect -3793 26776 -3786 26824
rect -3766 26776 -3760 26824
rect -3732 26816 -3727 26837
rect -3706 26826 -3702 26837
rect -3706 26816 -3701 26826
rect -3732 26789 -3715 26816
rect -3713 26789 -3711 26816
rect -3709 26789 -3706 26816
rect -3853 26737 -3844 26745
rect -3840 26737 -3834 26755
rect -3813 26751 -3793 26755
rect -3813 26748 -3802 26751
rect -3817 26747 -3802 26748
rect -3822 26745 -3820 26747
rect -3815 26745 -3808 26747
rect -3804 26745 -3802 26747
rect -3785 26745 -3778 26776
rect -3824 26742 -3815 26745
rect -3808 26742 -3799 26745
rect -3843 26697 -3834 26737
rect -3833 26697 -3827 26737
rect -3824 26697 -3817 26742
rect -3804 26737 -3802 26742
rect -3794 26737 -3786 26745
rect -3767 26737 -3760 26747
rect -3754 26745 -3750 26751
rect -3812 26697 -3808 26737
rect -3843 26689 -3827 26697
rect -3815 26689 -3808 26697
rect -3804 26697 -3796 26737
rect -3793 26697 -3787 26737
rect -3804 26661 -3802 26697
rect -3785 26689 -3778 26737
rect -3776 26697 -3768 26737
rect -3766 26697 -3760 26737
rect -3757 26689 -3750 26697
rect -3781 26677 -3780 26689
rect -3732 26677 -3730 26789
rect -3713 26781 -3709 26789
rect -3704 26768 -3701 26816
rect -3700 26789 -3688 26816
rect -3686 26781 -3684 26816
rect -3677 26789 -3674 26826
rect -3656 26819 -3651 26847
rect -3608 26839 -3603 26841
rect -3638 26829 -3634 26837
rect -3655 26789 -3651 26819
rect -3650 26789 -3639 26829
rect -3637 26789 -3634 26829
rect -3655 26781 -3652 26789
rect -3704 26689 -3701 26747
rect -3781 26669 -3776 26677
rect -3760 26669 -3714 26677
rect -3845 26653 -3836 26661
rect -3833 26653 -3824 26661
rect -3817 26653 -3808 26661
rect -3805 26653 -3796 26661
rect -3788 26653 -3780 26661
rect -3776 26653 -3768 26661
rect -3760 26653 -3752 26661
rect -3732 26658 -3730 26669
rect -3628 26667 -3624 26789
rect -3608 26667 -3602 26839
rect -3588 26829 -3586 26931
rect -3564 26901 -3562 26961
rect -3526 26915 -3523 26925
rect -3516 26917 -3514 26979
rect -3503 26977 -3498 26979
rect -3494 26953 -3487 26979
rect -3564 26885 -3556 26901
rect -3516 26893 -3512 26917
rect -3564 26861 -3555 26885
rect -3575 26841 -3572 26851
rect -3564 26841 -3562 26861
rect -3583 26839 -3576 26841
rect -3583 26829 -3575 26839
rect -3565 26829 -3562 26841
rect -3601 26793 -3592 26829
rect -3590 26793 -3585 26829
rect -3581 26793 -3575 26829
rect -3574 26793 -3558 26829
rect -3590 26785 -3583 26793
rect -3564 26785 -3558 26793
rect -3588 26658 -3586 26785
rect -3564 26658 -3562 26785
rect -3554 26667 -3548 26839
rect -3544 26833 -3538 26841
rect -3532 26793 -3526 26833
rect -3532 26667 -3528 26793
rect -3732 26653 -3720 26658
rect -3714 26653 -3704 26658
rect -3702 26653 -3692 26658
rect -3686 26653 -3676 26658
rect -3833 26652 -3817 26653
rect -3805 26652 -3789 26653
rect -3776 26652 -3760 26653
rect -3748 26652 -3740 26653
rect -3732 26652 -3714 26653
rect -3702 26652 -3686 26653
rect -3674 26652 -3664 26658
rect -4252 26642 -4242 26650
rect -4224 26642 -4214 26650
rect -4212 26639 -4210 26650
rect -4174 26642 -4166 26650
rect -4140 26642 -4138 26650
rect -4126 26642 -4124 26650
rect -4116 26639 -4114 26650
rect -4112 26642 -4110 26650
rect -4098 26642 -4096 26650
rect -4092 26639 -4090 26650
rect -4084 26642 -4082 26650
rect -4036 26642 -4026 26650
rect -4020 26639 -4018 26650
rect -4008 26642 -3998 26650
rect -3958 26642 -3950 26650
rect -3909 26645 -3894 26650
rect -3881 26645 -3866 26650
rect -3824 26645 -3817 26652
rect -3876 26639 -3874 26645
rect -3804 26639 -3802 26652
rect -3796 26645 -3789 26652
rect -3768 26645 -3760 26652
rect -3732 26639 -3730 26652
rect -3720 26642 -3714 26652
rect -3692 26642 -3686 26652
rect -3654 26650 -3646 26658
rect -3626 26650 -3612 26658
rect -3596 26650 -3584 26658
rect -3568 26650 -3556 26658
rect -3646 26642 -3638 26650
rect -3612 26642 -3610 26650
rect -3598 26642 -3596 26650
rect -3588 26639 -3586 26650
rect -3584 26642 -3582 26650
rect -3570 26642 -3568 26650
rect -3564 26639 -3562 26650
rect -3556 26642 -3554 26650
rect -3516 26639 -3514 26893
rect -3512 26667 -3506 26841
rect -3492 26833 -3490 26953
rect -3479 26841 -3476 26851
rect -3468 26841 -3466 26979
rect -3420 26917 -3418 26979
rect -3417 26953 -3401 26964
rect -3417 26917 -3411 26953
rect -3420 26916 -3411 26917
rect -3391 26916 -3389 26964
rect -3420 26893 -3416 26916
rect -3487 26833 -3479 26841
rect -3469 26833 -3466 26841
rect -3505 26793 -3496 26833
rect -3494 26793 -3489 26833
rect -3485 26793 -3479 26833
rect -3478 26793 -3462 26833
rect -3494 26785 -3487 26793
rect -3468 26785 -3462 26793
rect -3492 26658 -3490 26785
rect -3468 26658 -3466 26785
rect -3458 26667 -3452 26841
rect -3448 26833 -3442 26841
rect -3436 26793 -3430 26833
rect -3436 26667 -3432 26793
rect -3500 26650 -3490 26658
rect -3472 26650 -3464 26658
rect -3508 26642 -3500 26650
rect -3492 26639 -3490 26650
rect -3480 26642 -3472 26650
rect -3468 26639 -3466 26650
rect -3420 26639 -3418 26893
rect -3372 26658 -3370 26979
rect -3341 26916 -3329 26956
rect -3286 26916 -3279 26964
rect -3277 26916 -3271 26956
rect -3269 26908 -3262 26956
rect -3252 26658 -3250 26979
rect -3157 26972 -3154 26979
rect -3156 26956 -3154 26972
rect -3132 26966 -3130 26979
rect -3221 26916 -3209 26956
rect -3159 26908 -3154 26956
rect -3143 26953 -3140 26963
rect -3134 26953 -3133 26956
rect -3132 26953 -3123 26966
rect -3072 26956 -3068 26966
rect -3060 26956 -3058 26979
rect -3134 26937 -3130 26953
rect -3062 26942 -3058 26956
rect -3056 26945 -3048 26956
rect -3057 26942 -3048 26945
rect -3134 26908 -3133 26937
rect -3156 26849 -3154 26908
rect -3157 26791 -3153 26849
rect -3156 26658 -3154 26791
rect -3132 26658 -3130 26937
rect -3117 26895 -3115 26899
rect -3125 26791 -3123 26889
rect -3107 26881 -3105 26895
rect -3103 26791 -3099 26849
rect -3086 26831 -3082 26839
rect -3060 26837 -3058 26942
rect -3050 26932 -3041 26942
rect -3031 26932 -3024 26979
rect -3022 26977 -3020 26979
rect -3023 26955 -3020 26965
rect -3012 26955 -3010 26979
rect -3013 26939 -3010 26955
rect -2972 26948 -2963 26979
rect -2916 26971 -2914 26979
rect -2917 26961 -2912 26971
rect -2896 26961 -2890 26979
rect -2916 26957 -2912 26961
rect -3040 26929 -3031 26932
rect -3049 26847 -3040 26881
rect -3049 26837 -3039 26847
rect -3031 26837 -3024 26916
rect -3070 26831 -3051 26837
rect -3098 26791 -3087 26831
rect -3085 26791 -3082 26831
rect -3060 26827 -3051 26831
rect -3103 26783 -3100 26791
rect -3076 26667 -3072 26791
rect -3060 26789 -3050 26827
rect -3049 26789 -3043 26831
rect -3406 26650 -3396 26658
rect -3378 26650 -3368 26658
rect -3346 26650 -3338 26658
rect -3318 26650 -3302 26658
rect -3286 26650 -3274 26658
rect -3258 26650 -3246 26658
rect -3226 26650 -3218 26658
rect -3198 26650 -3182 26658
rect -3166 26650 -3154 26658
rect -3138 26650 -3126 26658
rect -3106 26650 -3098 26658
rect -3412 26642 -3406 26650
rect -3384 26642 -3378 26650
rect -3372 26639 -3370 26650
rect -3338 26642 -3330 26650
rect -3290 26642 -3286 26650
rect -3262 26642 -3258 26650
rect -3252 26639 -3250 26650
rect -3218 26642 -3210 26650
rect -3170 26642 -3166 26650
rect -3156 26639 -3154 26650
rect -3142 26642 -3138 26650
rect -3132 26639 -3130 26650
rect -3098 26642 -3090 26650
rect -3060 26639 -3058 26789
rect -3041 26783 -3034 26831
rect -3032 26783 -3023 26837
rect -3012 26831 -3010 26939
rect -2986 26934 -2984 26939
rect -2974 26934 -2972 26939
rect -2972 26929 -2964 26934
rect -2918 26931 -2911 26957
rect -2962 26924 -2954 26929
rect -2965 26883 -2959 26909
rect -2940 26908 -2938 26911
rect -3022 26789 -3016 26831
rect -3014 26783 -3007 26831
rect -3005 26789 -2996 26841
rect -2984 26819 -2979 26847
rect -2936 26839 -2931 26841
rect -2966 26829 -2962 26837
rect -2983 26789 -2979 26819
rect -2978 26789 -2967 26829
rect -2965 26789 -2962 26829
rect -3031 26781 -3024 26783
rect -3012 26658 -3010 26783
rect -2983 26781 -2980 26789
rect -2956 26667 -2952 26789
rect -2936 26667 -2930 26839
rect -2916 26829 -2914 26931
rect -2892 26901 -2890 26961
rect -2854 26915 -2851 26925
rect -2844 26917 -2842 26979
rect -2831 26977 -2826 26979
rect -2822 26953 -2815 26979
rect -2892 26885 -2884 26901
rect -2844 26893 -2840 26917
rect -2892 26861 -2883 26885
rect -2903 26841 -2900 26851
rect -2892 26841 -2890 26861
rect -2911 26839 -2904 26841
rect -2911 26829 -2903 26839
rect -2893 26829 -2890 26841
rect -2929 26793 -2920 26829
rect -2918 26793 -2913 26829
rect -2909 26793 -2903 26829
rect -2902 26793 -2886 26829
rect -2918 26785 -2911 26793
rect -2892 26785 -2886 26793
rect -2916 26658 -2914 26785
rect -2892 26658 -2890 26785
rect -2882 26667 -2876 26839
rect -2872 26833 -2866 26841
rect -2860 26793 -2854 26833
rect -2860 26667 -2856 26793
rect -3042 26650 -3034 26658
rect -3014 26650 -3006 26658
rect -2982 26650 -2974 26658
rect -2954 26650 -2940 26658
rect -2924 26650 -2912 26658
rect -2896 26650 -2884 26658
rect -3050 26642 -3042 26650
rect -3022 26642 -3014 26650
rect -3012 26639 -3010 26650
rect -2974 26642 -2966 26650
rect -2940 26642 -2938 26650
rect -2926 26642 -2924 26650
rect -2916 26639 -2914 26650
rect -2912 26642 -2910 26650
rect -2898 26642 -2896 26650
rect -2892 26639 -2890 26650
rect -2884 26642 -2882 26650
rect -2844 26639 -2842 26893
rect -2840 26667 -2834 26841
rect -2820 26833 -2818 26953
rect -2807 26841 -2804 26851
rect -2796 26841 -2794 26979
rect -2760 26956 -2755 26966
rect -2748 26956 -2745 26979
rect -2750 26953 -2736 26956
rect -2750 26942 -2745 26953
rect -2748 26917 -2745 26942
rect -2719 26932 -2712 26979
rect -2711 26955 -2708 26965
rect -2700 26955 -2698 26979
rect -2701 26939 -2698 26955
rect -2660 26948 -2651 26979
rect -2604 26971 -2602 26979
rect -2605 26961 -2600 26971
rect -2584 26961 -2578 26979
rect -2604 26957 -2600 26961
rect -2748 26893 -2744 26917
rect -2815 26833 -2807 26841
rect -2797 26833 -2794 26841
rect -2833 26793 -2824 26833
rect -2822 26793 -2817 26833
rect -2813 26793 -2807 26833
rect -2806 26793 -2790 26833
rect -2822 26785 -2815 26793
rect -2796 26785 -2790 26793
rect -2820 26658 -2818 26785
rect -2796 26658 -2794 26785
rect -2786 26667 -2780 26841
rect -2776 26833 -2770 26841
rect -2748 26837 -2746 26893
rect -2731 26847 -2728 26893
rect -2731 26837 -2721 26847
rect -2719 26837 -2712 26916
rect -2758 26833 -2739 26837
rect -2764 26793 -2758 26833
rect -2748 26827 -2739 26833
rect -2764 26667 -2760 26793
rect -2748 26789 -2738 26827
rect -2737 26789 -2731 26833
rect -2828 26650 -2818 26658
rect -2800 26650 -2792 26658
rect -2836 26642 -2828 26650
rect -2820 26639 -2818 26650
rect -2808 26642 -2800 26650
rect -2796 26639 -2794 26650
rect -2748 26639 -2746 26789
rect -2729 26785 -2722 26833
rect -2720 26785 -2711 26837
rect -2700 26833 -2698 26939
rect -2674 26934 -2672 26939
rect -2662 26934 -2660 26939
rect -2660 26929 -2652 26934
rect -2606 26931 -2599 26957
rect -2650 26924 -2642 26929
rect -2653 26883 -2647 26909
rect -2628 26908 -2626 26911
rect -2710 26789 -2704 26833
rect -2702 26785 -2695 26833
rect -2693 26789 -2684 26843
rect -2672 26819 -2667 26847
rect -2624 26839 -2619 26841
rect -2654 26829 -2650 26837
rect -2671 26789 -2667 26819
rect -2666 26789 -2655 26829
rect -2653 26789 -2650 26829
rect -2719 26781 -2712 26785
rect -2700 26658 -2698 26785
rect -2671 26781 -2668 26789
rect -2644 26667 -2640 26789
rect -2624 26667 -2618 26839
rect -2604 26829 -2602 26931
rect -2580 26901 -2578 26961
rect -2508 26969 -2503 26979
rect -2508 26953 -2505 26969
rect -2504 26967 -2503 26969
rect -2412 26969 -2408 26979
rect -2504 26953 -2496 26967
rect -2580 26885 -2572 26901
rect -2580 26861 -2571 26885
rect -2591 26841 -2588 26851
rect -2580 26841 -2578 26861
rect -2599 26839 -2592 26841
rect -2599 26829 -2591 26839
rect -2581 26829 -2578 26841
rect -2617 26793 -2608 26829
rect -2606 26793 -2601 26829
rect -2597 26793 -2591 26829
rect -2590 26793 -2574 26829
rect -2606 26785 -2599 26793
rect -2580 26785 -2574 26793
rect -2604 26658 -2602 26785
rect -2580 26658 -2578 26785
rect -2570 26667 -2564 26839
rect -2560 26833 -2554 26841
rect -2548 26793 -2542 26833
rect -2548 26667 -2544 26793
rect -2508 26658 -2506 26953
rect -2503 26919 -2496 26953
rect -2412 26959 -2402 26969
rect -2412 26913 -2410 26959
rect -2425 26911 -2410 26913
rect -2425 26903 -2420 26911
rect -2412 26903 -2410 26911
rect -2401 26911 -2386 26959
rect -2375 26953 -2372 26963
rect -2364 26953 -2362 26979
rect -2365 26937 -2362 26953
rect -2401 26903 -2392 26911
rect -2415 26889 -2410 26903
rect -2477 26667 -2468 26843
rect -2730 26650 -2724 26658
rect -2702 26650 -2696 26658
rect -2670 26650 -2662 26658
rect -2642 26650 -2628 26658
rect -2612 26650 -2600 26658
rect -2584 26650 -2572 26658
rect -2514 26650 -2506 26658
rect -2486 26650 -2480 26658
rect -2454 26650 -2446 26658
rect -2426 26650 -2414 26658
rect -2412 26650 -2410 26889
rect -2394 26839 -2385 26849
rect -2384 26667 -2375 26839
rect -2364 26658 -2362 26937
rect -2349 26895 -2347 26899
rect -2339 26881 -2337 26895
rect -2335 26791 -2331 26849
rect -2318 26831 -2314 26839
rect -2330 26791 -2319 26831
rect -2317 26791 -2314 26831
rect -2335 26783 -2332 26791
rect -2308 26667 -2304 26791
rect -2398 26650 -2386 26658
rect -2370 26650 -2358 26658
rect -2338 26650 -2330 26658
rect -2740 26642 -2730 26650
rect -2712 26642 -2702 26650
rect -2700 26639 -2698 26650
rect -2662 26642 -2654 26650
rect -2628 26642 -2626 26650
rect -2614 26642 -2612 26650
rect -2604 26639 -2602 26650
rect -2600 26642 -2598 26650
rect -2586 26642 -2584 26650
rect -2580 26639 -2578 26650
rect -2572 26642 -2570 26650
rect -2524 26642 -2514 26650
rect -2508 26639 -2506 26650
rect -2496 26642 -2486 26650
rect -2446 26642 -2438 26650
rect -2414 26642 -2410 26650
rect -2386 26642 -2382 26650
rect -2412 26639 -2410 26642
rect -2364 26639 -2362 26650
rect -2358 26642 -2354 26650
rect -2330 26642 -2322 26650
rect -2292 26639 -2290 26979
rect -2268 26977 -2254 26979
rect -2268 26969 -2266 26977
rect -2269 26961 -2264 26969
rect -2268 26955 -2264 26961
rect -2270 26929 -2263 26955
rect -2288 26667 -2282 26841
rect -2268 26831 -2266 26929
rect -2255 26841 -2252 26851
rect -2244 26841 -2242 26979
rect -2206 26915 -2203 26925
rect -2196 26917 -2194 26979
rect -2183 26977 -2178 26979
rect -2174 26953 -2167 26979
rect -2196 26893 -2192 26917
rect -2263 26831 -2255 26841
rect -2245 26831 -2242 26841
rect -2281 26793 -2272 26831
rect -2270 26793 -2265 26831
rect -2261 26793 -2255 26831
rect -2254 26793 -2238 26831
rect -2270 26785 -2263 26793
rect -2244 26785 -2238 26793
rect -2268 26658 -2266 26785
rect -2244 26658 -2242 26785
rect -2234 26667 -2228 26841
rect -2224 26833 -2218 26841
rect -2212 26793 -2206 26833
rect -2212 26667 -2208 26793
rect -2276 26650 -2266 26658
rect -2248 26650 -2238 26658
rect -2282 26642 -2276 26650
rect -2268 26639 -2266 26650
rect -2254 26642 -2248 26650
rect -2244 26639 -2242 26650
rect -2196 26639 -2194 26893
rect -2192 26667 -2186 26841
rect -2172 26833 -2170 26953
rect -2159 26841 -2156 26851
rect -2148 26841 -2146 26979
rect -2110 26915 -2107 26925
rect -2100 26917 -2098 26979
rect -2087 26977 -2082 26979
rect -2078 26953 -2071 26979
rect -2100 26893 -2096 26917
rect -2167 26833 -2159 26841
rect -2149 26833 -2146 26841
rect -2185 26793 -2176 26833
rect -2174 26793 -2169 26833
rect -2165 26793 -2159 26833
rect -2158 26793 -2142 26833
rect -2174 26785 -2167 26793
rect -2148 26785 -2142 26793
rect -2172 26658 -2170 26785
rect -2148 26658 -2146 26785
rect -2138 26667 -2132 26841
rect -2128 26833 -2122 26841
rect -2116 26793 -2110 26833
rect -2116 26667 -2112 26793
rect -2180 26650 -2170 26658
rect -2152 26650 -2144 26658
rect -2188 26642 -2180 26650
rect -2172 26639 -2170 26650
rect -2160 26642 -2152 26650
rect -2148 26639 -2146 26650
rect -2100 26639 -2098 26893
rect -2096 26667 -2090 26841
rect -2076 26833 -2074 26953
rect -2063 26841 -2060 26851
rect -2052 26841 -2050 26979
rect -1980 26969 -1975 26979
rect -1980 26953 -1977 26969
rect -1976 26967 -1975 26969
rect -1976 26953 -1968 26967
rect -2071 26833 -2063 26841
rect -2053 26833 -2050 26841
rect -2089 26793 -2080 26833
rect -2078 26793 -2073 26833
rect -2069 26793 -2063 26833
rect -2062 26793 -2046 26833
rect -2078 26785 -2071 26793
rect -2052 26785 -2046 26793
rect -2076 26658 -2074 26785
rect -2052 26658 -2050 26785
rect -2042 26667 -2036 26841
rect -2032 26833 -2026 26841
rect -2020 26793 -2014 26833
rect -2020 26667 -2016 26793
rect -1980 26658 -1978 26953
rect -1975 26919 -1968 26953
rect -1949 26667 -1940 26843
rect -2084 26650 -2074 26658
rect -2056 26650 -2048 26658
rect -1986 26650 -1978 26658
rect -1958 26650 -1952 26658
rect -1926 26650 -1918 26658
rect -1898 26650 -1886 26658
rect -1884 26650 -1882 26979
rect -1876 26964 -1874 26969
rect -1881 26916 -1874 26964
rect -1873 26916 -1857 26959
rect -1858 26911 -1857 26916
rect -1836 26658 -1834 26979
rect -1805 26916 -1793 26956
rect -1750 26916 -1743 26964
rect -1741 26916 -1735 26956
rect -1733 26908 -1726 26956
rect -1716 26658 -1714 26979
rect -1685 26916 -1673 26956
rect -1630 26916 -1623 26964
rect -1621 26916 -1615 26956
rect -1613 26908 -1606 26956
rect -1596 26658 -1594 26979
rect -1565 26916 -1553 26956
rect -1510 26916 -1503 26964
rect -1501 26916 -1495 26956
rect -1493 26908 -1486 26956
rect -1476 26658 -1474 26979
rect -1382 26977 -1375 26979
rect -1382 26966 -1373 26977
rect -1382 26961 -1365 26966
rect -1445 26916 -1433 26956
rect -1382 26900 -1375 26961
rect -1360 26908 -1357 26956
rect -1380 26851 -1378 26900
rect -1381 26667 -1374 26851
rect -1367 26841 -1364 26851
rect -1356 26841 -1354 26979
rect -1308 26917 -1306 26979
rect -1305 26953 -1289 26964
rect -1305 26917 -1299 26953
rect -1308 26916 -1299 26917
rect -1279 26916 -1277 26964
rect -1308 26893 -1304 26916
rect -1357 26793 -1354 26841
rect -1336 26833 -1330 26841
rect -1380 26658 -1378 26667
rect -1356 26658 -1354 26793
rect -1324 26793 -1318 26833
rect -1324 26667 -1320 26793
rect -1870 26650 -1858 26658
rect -1842 26650 -1830 26658
rect -1810 26650 -1802 26658
rect -1782 26650 -1766 26658
rect -1750 26650 -1738 26658
rect -1722 26650 -1710 26658
rect -1690 26650 -1682 26658
rect -1662 26650 -1646 26658
rect -1630 26650 -1618 26658
rect -1602 26650 -1590 26658
rect -1570 26650 -1562 26658
rect -1542 26650 -1526 26658
rect -1510 26650 -1498 26658
rect -1482 26650 -1470 26658
rect -1450 26650 -1442 26658
rect -1388 26650 -1378 26658
rect -1360 26650 -1350 26658
rect -2092 26642 -2084 26650
rect -2076 26639 -2074 26650
rect -2064 26642 -2056 26650
rect -2052 26639 -2050 26650
rect -1996 26642 -1986 26650
rect -1980 26639 -1978 26650
rect -1968 26642 -1958 26650
rect -1918 26642 -1910 26650
rect -1886 26642 -1882 26650
rect -1858 26642 -1854 26650
rect -1884 26639 -1882 26642
rect -1836 26639 -1834 26650
rect -1830 26642 -1826 26650
rect -1802 26642 -1794 26650
rect -1754 26642 -1750 26650
rect -1726 26642 -1722 26650
rect -1716 26639 -1714 26650
rect -1682 26642 -1674 26650
rect -1634 26642 -1630 26650
rect -1606 26642 -1602 26650
rect -1596 26639 -1594 26650
rect -1562 26642 -1554 26650
rect -1514 26642 -1510 26650
rect -1486 26642 -1482 26650
rect -1476 26639 -1474 26650
rect -1442 26642 -1434 26650
rect -1394 26642 -1388 26650
rect -1380 26639 -1378 26650
rect -1366 26642 -1360 26650
rect -1356 26639 -1354 26650
rect -1308 26639 -1306 26893
rect -1260 26658 -1258 26979
rect -1166 26977 -1159 26979
rect -1166 26966 -1157 26977
rect -1166 26961 -1149 26966
rect -1229 26916 -1217 26956
rect -1166 26900 -1159 26961
rect -1144 26908 -1141 26956
rect -1164 26851 -1162 26900
rect -1165 26667 -1158 26851
rect -1151 26841 -1148 26851
rect -1140 26841 -1138 26979
rect -1068 26969 -1063 26979
rect -1068 26953 -1065 26969
rect -1064 26967 -1063 26969
rect -944 26967 -935 26969
rect -1064 26953 -1056 26967
rect -1141 26793 -1138 26841
rect -1120 26833 -1114 26841
rect -1164 26658 -1162 26667
rect -1140 26658 -1138 26793
rect -1108 26793 -1102 26833
rect -1108 26667 -1104 26793
rect -1068 26658 -1066 26953
rect -1063 26919 -1056 26953
rect -944 26919 -933 26967
rect -852 26921 -850 26979
rect -849 26969 -848 26979
rect -849 26921 -842 26969
rect -829 26961 -815 26969
rect -852 26915 -842 26921
rect -1037 26667 -1028 26843
rect -852 26658 -850 26915
rect -841 26911 -838 26915
rect -830 26911 -825 26959
rect -831 26841 -825 26851
rect -815 26841 -812 26851
rect -804 26841 -802 26979
rect -768 26956 -763 26966
rect -756 26956 -753 26979
rect -758 26953 -744 26956
rect -758 26942 -753 26953
rect -756 26917 -753 26942
rect -727 26932 -720 26979
rect -719 26955 -716 26965
rect -708 26955 -706 26979
rect -709 26939 -706 26955
rect -668 26948 -659 26979
rect -612 26971 -610 26979
rect -613 26961 -608 26971
rect -592 26961 -586 26979
rect -612 26957 -608 26961
rect -756 26893 -752 26917
rect -821 26793 -815 26841
rect -805 26793 -802 26841
rect -784 26833 -778 26841
rect -756 26837 -754 26893
rect -739 26847 -736 26893
rect -739 26837 -729 26847
rect -727 26837 -720 26916
rect -766 26833 -747 26837
rect -804 26658 -802 26793
rect -772 26793 -766 26833
rect -756 26827 -747 26833
rect -772 26667 -768 26793
rect -756 26789 -746 26827
rect -745 26789 -739 26833
rect -1294 26650 -1284 26658
rect -1266 26650 -1256 26658
rect -1234 26650 -1226 26658
rect -1172 26650 -1162 26658
rect -1144 26650 -1134 26658
rect -1074 26650 -1066 26658
rect -1046 26650 -1040 26658
rect -1014 26650 -1006 26658
rect -986 26650 -970 26658
rect -954 26650 -942 26658
rect -926 26650 -914 26658
rect -894 26650 -886 26658
rect -866 26650 -850 26658
rect -836 26650 -824 26658
rect -808 26650 -796 26658
rect -1300 26642 -1294 26650
rect -1272 26642 -1266 26650
rect -1260 26639 -1258 26650
rect -1226 26642 -1218 26650
rect -1178 26642 -1172 26650
rect -1164 26639 -1162 26650
rect -1150 26642 -1144 26650
rect -1140 26639 -1138 26650
rect -1084 26642 -1074 26650
rect -1068 26639 -1066 26650
rect -1056 26642 -1046 26650
rect -1006 26642 -998 26650
rect -958 26642 -954 26650
rect -930 26642 -926 26650
rect -886 26642 -878 26650
rect -852 26639 -850 26650
rect -838 26642 -836 26650
rect -824 26642 -822 26650
rect -810 26642 -808 26650
rect -804 26639 -802 26650
rect -796 26642 -794 26650
rect -756 26639 -754 26789
rect -737 26785 -730 26833
rect -728 26785 -719 26837
rect -708 26833 -706 26939
rect -682 26934 -680 26939
rect -670 26934 -668 26939
rect -668 26929 -660 26934
rect -614 26931 -607 26957
rect -658 26924 -650 26929
rect -661 26883 -655 26909
rect -636 26908 -634 26911
rect -718 26789 -712 26833
rect -710 26785 -703 26833
rect -701 26789 -692 26843
rect -680 26819 -675 26847
rect -632 26839 -627 26841
rect -662 26829 -658 26837
rect -679 26789 -675 26819
rect -674 26789 -663 26829
rect -661 26789 -658 26829
rect -727 26781 -720 26785
rect -708 26658 -706 26785
rect -679 26781 -676 26789
rect -652 26667 -648 26789
rect -632 26667 -626 26839
rect -612 26829 -610 26931
rect -588 26901 -586 26961
rect -550 26915 -547 26925
rect -540 26917 -538 26979
rect -527 26977 -522 26979
rect -518 26953 -511 26979
rect -588 26885 -580 26901
rect -540 26893 -536 26917
rect -588 26861 -579 26885
rect -599 26841 -596 26851
rect -588 26841 -586 26861
rect -607 26839 -600 26841
rect -607 26829 -599 26839
rect -589 26829 -586 26841
rect -625 26793 -616 26829
rect -614 26793 -609 26829
rect -605 26793 -599 26829
rect -598 26793 -582 26829
rect -614 26785 -607 26793
rect -588 26785 -582 26793
rect -612 26658 -610 26785
rect -588 26658 -586 26785
rect -578 26667 -572 26839
rect -568 26833 -562 26841
rect -556 26793 -550 26833
rect -556 26667 -552 26793
rect -738 26650 -732 26658
rect -710 26650 -704 26658
rect -678 26650 -670 26658
rect -650 26650 -636 26658
rect -620 26650 -608 26658
rect -592 26650 -580 26658
rect -748 26642 -738 26650
rect -720 26642 -710 26650
rect -708 26639 -706 26650
rect -670 26642 -662 26650
rect -636 26642 -634 26650
rect -622 26642 -620 26650
rect -612 26639 -610 26650
rect -608 26642 -606 26650
rect -594 26642 -592 26650
rect -588 26639 -586 26650
rect -580 26642 -578 26650
rect -540 26639 -538 26893
rect -536 26667 -530 26841
rect -516 26833 -514 26953
rect -503 26841 -500 26851
rect -492 26841 -490 26979
rect -456 26956 -451 26966
rect -444 26956 -441 26979
rect -446 26953 -432 26956
rect -446 26942 -441 26953
rect -444 26917 -441 26942
rect -415 26932 -408 26979
rect -407 26955 -404 26965
rect -396 26955 -394 26979
rect -397 26939 -394 26955
rect -356 26948 -347 26979
rect -300 26971 -298 26979
rect -301 26961 -296 26971
rect -280 26961 -274 26979
rect -300 26957 -296 26961
rect -444 26893 -440 26917
rect -511 26833 -503 26841
rect -493 26833 -490 26841
rect -529 26793 -520 26833
rect -518 26793 -513 26833
rect -509 26793 -503 26833
rect -502 26793 -486 26833
rect -518 26785 -511 26793
rect -492 26785 -486 26793
rect -516 26658 -514 26785
rect -492 26658 -490 26785
rect -482 26667 -476 26841
rect -472 26833 -466 26841
rect -444 26837 -442 26893
rect -427 26847 -424 26893
rect -427 26837 -417 26847
rect -415 26837 -408 26916
rect -454 26833 -435 26837
rect -460 26793 -454 26833
rect -444 26827 -435 26833
rect -460 26667 -456 26793
rect -444 26789 -434 26827
rect -433 26789 -427 26833
rect -524 26650 -514 26658
rect -496 26650 -488 26658
rect -532 26642 -524 26650
rect -516 26639 -514 26650
rect -504 26642 -496 26650
rect -492 26639 -490 26650
rect -444 26639 -442 26789
rect -425 26785 -418 26833
rect -416 26785 -407 26837
rect -396 26833 -394 26939
rect -370 26934 -368 26939
rect -358 26934 -356 26939
rect -356 26929 -348 26934
rect -302 26931 -295 26957
rect -346 26924 -338 26929
rect -349 26883 -343 26909
rect -324 26908 -322 26911
rect -406 26789 -400 26833
rect -398 26785 -391 26833
rect -389 26789 -380 26843
rect -368 26819 -363 26847
rect -320 26839 -315 26841
rect -350 26829 -346 26837
rect -367 26789 -363 26819
rect -362 26789 -351 26829
rect -349 26789 -346 26829
rect -415 26781 -408 26785
rect -396 26658 -394 26785
rect -367 26781 -364 26789
rect -340 26667 -336 26789
rect -320 26667 -314 26839
rect -300 26829 -298 26931
rect -276 26901 -274 26961
rect -204 26969 -199 26979
rect -204 26953 -201 26969
rect -200 26967 -199 26969
rect -200 26953 -192 26967
rect -276 26885 -268 26901
rect -276 26861 -267 26885
rect -287 26841 -284 26851
rect -276 26841 -274 26861
rect -295 26839 -288 26841
rect -295 26829 -287 26839
rect -277 26829 -274 26841
rect -313 26793 -304 26829
rect -302 26793 -297 26829
rect -293 26793 -287 26829
rect -286 26793 -270 26829
rect -302 26785 -295 26793
rect -276 26785 -270 26793
rect -300 26658 -298 26785
rect -276 26658 -274 26785
rect -266 26667 -260 26839
rect -256 26833 -250 26841
rect -244 26793 -238 26833
rect -244 26667 -240 26793
rect -204 26658 -202 26953
rect -199 26919 -192 26953
rect -108 26921 -106 26979
rect -105 26969 -104 26979
rect -105 26921 -98 26969
rect -85 26961 -71 26969
rect -108 26915 -98 26921
rect -173 26667 -164 26843
rect -108 26658 -106 26915
rect -97 26911 -94 26915
rect -86 26911 -81 26959
rect -87 26841 -81 26851
rect -71 26841 -68 26851
rect -60 26841 -58 26979
rect 12 26969 17 26979
rect 12 26953 15 26969
rect 16 26967 17 26969
rect 16 26953 24 26967
rect -77 26793 -71 26841
rect -61 26793 -58 26841
rect -40 26833 -34 26841
rect -60 26658 -58 26793
rect -28 26793 -22 26833
rect -28 26667 -24 26793
rect 12 26658 14 26953
rect 17 26919 24 26953
rect 108 26921 110 26979
rect 111 26969 112 26979
rect 111 26921 118 26969
rect 131 26961 145 26969
rect 108 26915 118 26921
rect 43 26667 52 26843
rect 108 26658 110 26915
rect 119 26911 122 26915
rect 130 26911 135 26959
rect 129 26841 135 26851
rect 145 26841 148 26851
rect 156 26841 158 26979
rect 194 26915 197 26925
rect 204 26917 206 26979
rect 217 26977 222 26979
rect 226 26953 233 26979
rect 204 26893 208 26917
rect 139 26793 145 26841
rect 155 26793 158 26841
rect 176 26833 182 26841
rect 156 26658 158 26793
rect 188 26793 194 26833
rect 188 26667 192 26793
rect -426 26650 -420 26658
rect -398 26650 -392 26658
rect -366 26650 -358 26658
rect -338 26650 -324 26658
rect -308 26650 -296 26658
rect -280 26650 -268 26658
rect -210 26650 -202 26658
rect -182 26650 -176 26658
rect -150 26650 -142 26658
rect -122 26650 -106 26658
rect -92 26650 -80 26658
rect -64 26650 -52 26658
rect 6 26650 14 26658
rect 34 26650 40 26658
rect 66 26650 74 26658
rect 94 26650 110 26658
rect 124 26650 136 26658
rect 152 26650 164 26658
rect -436 26642 -426 26650
rect -408 26642 -398 26650
rect -396 26639 -394 26650
rect -358 26642 -350 26650
rect -324 26642 -322 26650
rect -310 26642 -308 26650
rect -300 26639 -298 26650
rect -296 26642 -294 26650
rect -282 26642 -280 26650
rect -276 26639 -274 26650
rect -268 26642 -266 26650
rect -220 26642 -210 26650
rect -204 26639 -202 26650
rect -192 26642 -182 26650
rect -142 26642 -134 26650
rect -108 26639 -106 26650
rect -94 26642 -92 26650
rect -80 26642 -78 26650
rect -66 26642 -64 26650
rect -60 26639 -58 26650
rect -52 26642 -50 26650
rect -4 26642 6 26650
rect 12 26639 14 26650
rect 24 26642 34 26650
rect 74 26642 82 26650
rect 108 26639 110 26650
rect 122 26642 124 26650
rect 136 26642 138 26650
rect 150 26642 152 26650
rect 156 26639 158 26650
rect 164 26642 166 26650
rect 204 26639 206 26893
rect 208 26667 214 26841
rect 228 26833 230 26953
rect 241 26841 244 26851
rect 252 26841 254 26979
rect 300 26917 302 26979
rect 303 26953 319 26964
rect 303 26917 309 26953
rect 300 26916 309 26917
rect 329 26916 331 26964
rect 300 26893 304 26916
rect 233 26833 241 26841
rect 251 26833 254 26841
rect 215 26793 224 26833
rect 226 26793 231 26833
rect 235 26793 241 26833
rect 242 26793 258 26833
rect 226 26785 233 26793
rect 252 26785 258 26793
rect 228 26658 230 26785
rect 252 26658 254 26785
rect 262 26667 268 26841
rect 272 26833 278 26841
rect 284 26793 290 26833
rect 284 26667 288 26793
rect 220 26650 230 26658
rect 248 26650 256 26658
rect 212 26642 220 26650
rect 228 26639 230 26650
rect 240 26642 248 26650
rect 252 26639 254 26650
rect 300 26639 302 26893
rect 348 26658 350 26979
rect 379 26916 391 26956
rect 434 26916 441 26964
rect 443 26916 449 26956
rect 451 26908 458 26956
rect 468 26658 470 26979
rect 562 26977 569 26979
rect 562 26966 571 26977
rect 562 26961 579 26966
rect 499 26916 511 26956
rect 562 26900 569 26961
rect 584 26908 587 26956
rect 564 26851 566 26900
rect 563 26667 570 26851
rect 577 26841 580 26851
rect 588 26841 590 26979
rect 626 26915 629 26925
rect 636 26917 638 26979
rect 649 26977 654 26979
rect 658 26953 665 26979
rect 636 26893 640 26917
rect 587 26793 590 26841
rect 608 26833 614 26841
rect 564 26658 566 26667
rect 588 26658 590 26793
rect 620 26793 626 26833
rect 620 26667 624 26793
rect 314 26650 324 26658
rect 342 26650 352 26658
rect 374 26650 382 26658
rect 402 26650 418 26658
rect 434 26650 446 26658
rect 462 26650 474 26658
rect 494 26650 502 26658
rect 556 26650 566 26658
rect 584 26650 594 26658
rect 308 26642 314 26650
rect 336 26642 342 26650
rect 348 26639 350 26650
rect 382 26642 390 26650
rect 430 26642 434 26650
rect 458 26642 462 26650
rect 468 26639 470 26650
rect 502 26642 510 26650
rect 550 26642 556 26650
rect 564 26639 566 26650
rect 578 26642 584 26650
rect 588 26639 590 26650
rect 636 26639 638 26893
rect 640 26667 646 26841
rect 660 26833 662 26953
rect 673 26841 676 26851
rect 684 26841 686 26979
rect 732 26917 735 26979
rect 752 26972 761 26979
rect 756 26969 760 26972
rect 756 26953 759 26969
rect 719 26907 724 26913
rect 719 26903 726 26907
rect 732 26903 736 26917
rect 729 26893 736 26903
rect 729 26889 734 26893
rect 732 26843 734 26889
rect 749 26849 753 26889
rect 756 26849 758 26953
rect 665 26833 673 26841
rect 683 26833 686 26841
rect 647 26793 656 26833
rect 658 26793 663 26833
rect 667 26793 673 26833
rect 674 26793 690 26833
rect 658 26785 665 26793
rect 684 26785 690 26793
rect 660 26658 662 26785
rect 684 26658 686 26785
rect 694 26667 700 26841
rect 704 26833 710 26841
rect 716 26793 722 26833
rect 716 26667 720 26793
rect 732 26791 742 26843
rect 749 26839 759 26849
rect 761 26839 768 26972
rect 769 26953 772 26963
rect 780 26953 782 26979
rect 779 26937 782 26953
rect 756 26833 758 26839
rect 743 26791 749 26833
rect 652 26650 662 26658
rect 680 26650 688 26658
rect 644 26642 652 26650
rect 660 26639 662 26650
rect 672 26642 680 26650
rect 684 26639 686 26650
rect 732 26639 734 26791
rect 751 26785 758 26833
rect 760 26785 769 26839
rect 780 26833 782 26937
rect 876 26969 878 26979
rect 876 26955 880 26969
rect 881 26955 888 26967
rect 876 26945 888 26955
rect 795 26895 797 26899
rect 805 26881 807 26895
rect 770 26791 776 26833
rect 778 26785 785 26833
rect 787 26791 796 26843
rect 809 26791 813 26849
rect 826 26831 830 26839
rect 814 26791 825 26831
rect 827 26791 830 26831
rect 756 26658 758 26785
rect 761 26783 768 26785
rect 780 26658 782 26785
rect 809 26783 812 26791
rect 836 26667 840 26791
rect 876 26658 878 26945
rect 880 26929 888 26945
rect 881 26919 888 26929
rect 972 26921 974 26979
rect 975 26969 976 26979
rect 975 26921 982 26969
rect 995 26961 1009 26969
rect 972 26915 982 26921
rect 907 26667 916 26841
rect 972 26658 974 26915
rect 983 26911 986 26915
rect 994 26911 999 26959
rect 993 26841 999 26851
rect 1009 26841 1012 26851
rect 1020 26841 1022 26979
rect 1058 26915 1061 26925
rect 1068 26917 1070 26979
rect 1081 26977 1086 26979
rect 1090 26953 1097 26979
rect 1068 26893 1072 26917
rect 1003 26793 1009 26841
rect 1019 26793 1022 26841
rect 1040 26833 1046 26841
rect 1020 26658 1022 26793
rect 1052 26793 1058 26833
rect 1052 26667 1056 26793
rect 746 26650 758 26658
rect 774 26650 784 26658
rect 806 26650 814 26658
rect 870 26650 878 26658
rect 898 26650 906 26658
rect 930 26650 938 26658
rect 958 26650 974 26658
rect 988 26650 1000 26658
rect 1016 26650 1028 26658
rect 740 26642 746 26650
rect 756 26639 758 26650
rect 768 26642 774 26650
rect 780 26639 782 26650
rect 814 26642 822 26650
rect 862 26642 870 26650
rect 876 26639 878 26650
rect 890 26642 898 26650
rect 938 26642 946 26650
rect 972 26639 974 26650
rect 986 26642 988 26650
rect 1000 26642 1002 26650
rect 1014 26642 1016 26650
rect 1020 26639 1022 26650
rect 1028 26642 1030 26650
rect 1068 26639 1070 26893
rect 1072 26667 1078 26841
rect 1092 26833 1094 26953
rect 1105 26841 1108 26851
rect 1116 26841 1118 26979
rect 1152 26956 1157 26966
rect 1164 26956 1167 26979
rect 1162 26953 1176 26956
rect 1162 26942 1167 26953
rect 1164 26917 1167 26942
rect 1193 26932 1200 26979
rect 1201 26955 1204 26965
rect 1212 26955 1214 26979
rect 1211 26939 1214 26955
rect 1252 26948 1261 26979
rect 1308 26971 1310 26979
rect 1307 26961 1312 26971
rect 1328 26961 1334 26979
rect 1308 26957 1312 26961
rect 1164 26893 1168 26917
rect 1097 26833 1105 26841
rect 1115 26833 1118 26841
rect 1079 26793 1088 26833
rect 1090 26793 1095 26833
rect 1099 26793 1105 26833
rect 1106 26793 1122 26833
rect 1090 26785 1097 26793
rect 1116 26785 1122 26793
rect 1092 26658 1094 26785
rect 1116 26658 1118 26785
rect 1126 26667 1132 26841
rect 1136 26833 1142 26841
rect 1164 26837 1166 26893
rect 1181 26847 1184 26893
rect 1181 26837 1191 26847
rect 1193 26837 1200 26916
rect 1154 26833 1173 26837
rect 1148 26793 1154 26833
rect 1164 26827 1173 26833
rect 1148 26667 1152 26793
rect 1164 26789 1174 26827
rect 1175 26789 1181 26833
rect 1084 26650 1094 26658
rect 1112 26650 1120 26658
rect 1076 26642 1084 26650
rect 1092 26639 1094 26650
rect 1104 26642 1112 26650
rect 1116 26639 1118 26650
rect 1164 26639 1166 26789
rect 1183 26785 1190 26833
rect 1192 26785 1201 26837
rect 1212 26833 1214 26939
rect 1238 26934 1240 26939
rect 1250 26934 1252 26939
rect 1252 26929 1260 26934
rect 1306 26931 1313 26957
rect 1262 26924 1270 26929
rect 1259 26883 1265 26909
rect 1284 26908 1286 26911
rect 1202 26789 1208 26833
rect 1210 26785 1217 26833
rect 1219 26789 1228 26843
rect 1240 26819 1245 26847
rect 1288 26839 1293 26841
rect 1258 26829 1262 26837
rect 1241 26789 1245 26819
rect 1246 26789 1257 26829
rect 1259 26789 1262 26829
rect 1193 26781 1200 26785
rect 1212 26658 1214 26785
rect 1241 26781 1244 26789
rect 1268 26667 1272 26789
rect 1288 26667 1294 26839
rect 1308 26829 1310 26931
rect 1332 26901 1334 26961
rect 1380 26917 1382 26979
rect 1383 26953 1399 26964
rect 1383 26917 1389 26953
rect 1380 26916 1389 26917
rect 1409 26916 1411 26964
rect 1332 26885 1340 26901
rect 1380 26893 1384 26916
rect 1332 26861 1341 26885
rect 1321 26841 1324 26851
rect 1332 26841 1334 26861
rect 1313 26839 1320 26841
rect 1313 26829 1321 26839
rect 1331 26829 1334 26841
rect 1295 26793 1304 26829
rect 1306 26793 1311 26829
rect 1315 26793 1321 26829
rect 1322 26793 1338 26829
rect 1306 26785 1313 26793
rect 1332 26785 1338 26793
rect 1308 26658 1310 26785
rect 1332 26658 1334 26785
rect 1342 26667 1348 26839
rect 1352 26833 1358 26841
rect 1364 26793 1370 26833
rect 1364 26667 1368 26793
rect 1182 26650 1188 26658
rect 1210 26650 1216 26658
rect 1242 26650 1250 26658
rect 1270 26650 1284 26658
rect 1300 26650 1312 26658
rect 1328 26650 1340 26658
rect 1172 26642 1182 26650
rect 1200 26642 1210 26650
rect 1212 26639 1214 26650
rect 1250 26642 1258 26650
rect 1284 26642 1286 26650
rect 1298 26642 1300 26650
rect 1308 26639 1310 26650
rect 1312 26642 1314 26650
rect 1326 26642 1328 26650
rect 1332 26639 1334 26650
rect 1340 26642 1342 26650
rect 1380 26639 1382 26893
rect 1428 26658 1430 26979
rect 1522 26977 1529 26979
rect 1522 26966 1531 26977
rect 1522 26961 1539 26966
rect 1459 26916 1471 26956
rect 1522 26900 1529 26961
rect 1544 26908 1547 26956
rect 1524 26851 1526 26900
rect 1523 26667 1530 26851
rect 1537 26841 1540 26851
rect 1548 26841 1550 26979
rect 1586 26915 1589 26925
rect 1596 26917 1598 26979
rect 1609 26977 1614 26979
rect 1618 26953 1625 26979
rect 1596 26893 1600 26917
rect 1547 26793 1550 26841
rect 1568 26833 1574 26841
rect 1524 26658 1526 26667
rect 1548 26658 1550 26793
rect 1580 26793 1586 26833
rect 1580 26667 1584 26793
rect 1394 26650 1404 26658
rect 1422 26650 1432 26658
rect 1454 26650 1462 26658
rect 1516 26650 1526 26658
rect 1544 26650 1554 26658
rect 1388 26642 1394 26650
rect 1416 26642 1422 26650
rect 1428 26639 1430 26650
rect 1462 26642 1470 26650
rect 1510 26642 1516 26650
rect 1524 26639 1526 26650
rect 1538 26642 1544 26650
rect 1548 26639 1550 26650
rect 1596 26639 1598 26893
rect 1600 26667 1606 26841
rect 1620 26833 1622 26953
rect 1633 26841 1636 26851
rect 1644 26841 1646 26979
rect 1682 26915 1685 26925
rect 1692 26917 1694 26979
rect 1705 26977 1710 26979
rect 1714 26953 1721 26979
rect 1692 26893 1696 26917
rect 1625 26833 1633 26841
rect 1643 26833 1646 26841
rect 1607 26793 1616 26833
rect 1618 26793 1623 26833
rect 1627 26793 1633 26833
rect 1634 26793 1650 26833
rect 1618 26785 1625 26793
rect 1644 26785 1650 26793
rect 1620 26658 1622 26785
rect 1644 26658 1646 26785
rect 1654 26667 1660 26841
rect 1664 26833 1670 26841
rect 1676 26793 1682 26833
rect 1676 26667 1680 26793
rect 1612 26650 1622 26658
rect 1640 26650 1648 26658
rect 1604 26642 1612 26650
rect 1620 26639 1622 26650
rect 1632 26642 1640 26650
rect 1644 26639 1646 26650
rect 1692 26639 1694 26893
rect 1696 26667 1702 26841
rect 1716 26833 1718 26953
rect 1729 26841 1732 26851
rect 1740 26841 1742 26979
rect 1778 26915 1781 26925
rect 1788 26917 1790 26979
rect 1801 26977 1806 26979
rect 1810 26953 1817 26979
rect 1788 26893 1792 26917
rect 1721 26833 1729 26841
rect 1739 26833 1742 26841
rect 1703 26793 1712 26833
rect 1714 26793 1719 26833
rect 1723 26793 1729 26833
rect 1730 26793 1746 26833
rect 1714 26785 1721 26793
rect 1740 26785 1746 26793
rect 1716 26658 1718 26785
rect 1740 26658 1742 26785
rect 1750 26667 1756 26841
rect 1760 26833 1766 26841
rect 1772 26793 1778 26833
rect 1772 26667 1776 26793
rect 1708 26650 1718 26658
rect 1736 26650 1744 26658
rect 1700 26642 1708 26650
rect 1716 26639 1718 26650
rect 1728 26642 1736 26650
rect 1740 26639 1742 26650
rect 1788 26639 1790 26893
rect 1792 26667 1798 26841
rect 1812 26833 1814 26953
rect 1825 26841 1828 26851
rect 1836 26841 1838 26979
rect 1874 26915 1877 26925
rect 1884 26917 1886 26979
rect 1897 26977 1902 26979
rect 1906 26953 1913 26979
rect 1884 26893 1888 26917
rect 1817 26833 1825 26841
rect 1835 26833 1838 26841
rect 1799 26793 1808 26833
rect 1810 26793 1815 26833
rect 1819 26793 1825 26833
rect 1826 26793 1842 26833
rect 1810 26785 1817 26793
rect 1836 26785 1842 26793
rect 1812 26658 1814 26785
rect 1836 26658 1838 26785
rect 1846 26667 1852 26841
rect 1856 26833 1862 26841
rect 1868 26793 1874 26833
rect 1868 26667 1872 26793
rect 1804 26650 1814 26658
rect 1832 26650 1840 26658
rect 1796 26642 1804 26650
rect 1812 26639 1814 26650
rect 1824 26642 1832 26650
rect 1836 26639 1838 26650
rect 1884 26639 1886 26893
rect 1888 26667 1894 26841
rect 1908 26833 1910 26953
rect 1921 26841 1924 26851
rect 1932 26841 1934 26979
rect 1970 26915 1973 26925
rect 1980 26917 1982 26979
rect 1993 26977 1998 26979
rect 2002 26953 2009 26979
rect 1980 26893 1984 26917
rect 1913 26833 1921 26841
rect 1931 26833 1934 26841
rect 1895 26793 1904 26833
rect 1906 26793 1911 26833
rect 1915 26793 1921 26833
rect 1922 26793 1938 26833
rect 1906 26785 1913 26793
rect 1932 26785 1938 26793
rect 1908 26658 1910 26785
rect 1932 26658 1934 26785
rect 1942 26667 1948 26841
rect 1952 26833 1958 26841
rect 1964 26793 1970 26833
rect 1964 26667 1968 26793
rect 1900 26650 1910 26658
rect 1928 26650 1936 26658
rect 1892 26642 1900 26650
rect 1908 26639 1910 26650
rect 1920 26642 1928 26650
rect 1932 26639 1934 26650
rect 1980 26639 1982 26893
rect 1984 26667 1990 26841
rect 2004 26833 2006 26953
rect 2017 26841 2020 26851
rect 2028 26841 2030 26979
rect 2066 26915 2069 26925
rect 2076 26917 2078 26979
rect 2089 26977 2094 26979
rect 2098 26953 2105 26979
rect 2076 26893 2080 26917
rect 2009 26833 2017 26841
rect 2027 26833 2030 26841
rect 1991 26793 2000 26833
rect 2002 26793 2007 26833
rect 2011 26793 2017 26833
rect 2018 26793 2034 26833
rect 2002 26785 2009 26793
rect 2028 26785 2034 26793
rect 2004 26658 2006 26785
rect 2028 26658 2030 26785
rect 2038 26667 2044 26841
rect 2048 26833 2054 26841
rect 2060 26793 2066 26833
rect 2060 26667 2064 26793
rect 1996 26650 2006 26658
rect 2024 26650 2032 26658
rect 1988 26642 1996 26650
rect 2004 26639 2006 26650
rect 2016 26642 2024 26650
rect 2028 26639 2030 26650
rect 2076 26639 2078 26893
rect 2080 26667 2086 26841
rect 2100 26833 2102 26953
rect 2113 26841 2116 26851
rect 2124 26841 2126 26979
rect 2162 26915 2165 26925
rect 2172 26917 2174 26979
rect 2185 26977 2190 26979
rect 2194 26953 2201 26979
rect 2172 26893 2176 26917
rect 2105 26833 2113 26841
rect 2123 26833 2126 26841
rect 2087 26793 2096 26833
rect 2098 26793 2103 26833
rect 2107 26793 2113 26833
rect 2114 26793 2130 26833
rect 2098 26785 2105 26793
rect 2124 26785 2130 26793
rect 2100 26658 2102 26785
rect 2124 26658 2126 26785
rect 2134 26667 2140 26841
rect 2144 26833 2150 26841
rect 2156 26793 2162 26833
rect 2156 26667 2160 26793
rect 2092 26650 2102 26658
rect 2120 26650 2128 26658
rect 2084 26642 2092 26650
rect 2100 26639 2102 26650
rect 2112 26642 2120 26650
rect 2124 26639 2126 26650
rect 2172 26639 2174 26893
rect 2176 26667 2182 26841
rect 2196 26833 2198 26953
rect 2209 26841 2212 26851
rect 2220 26841 2222 26979
rect 2258 26915 2261 26925
rect 2268 26917 2270 26979
rect 2281 26977 2286 26979
rect 2290 26953 2297 26979
rect 2268 26893 2272 26917
rect 2201 26833 2209 26841
rect 2219 26833 2222 26841
rect 2183 26793 2192 26833
rect 2194 26793 2199 26833
rect 2203 26793 2209 26833
rect 2210 26793 2226 26833
rect 2194 26785 2201 26793
rect 2220 26785 2226 26793
rect 2196 26658 2198 26785
rect 2220 26658 2222 26785
rect 2230 26667 2236 26841
rect 2240 26833 2246 26841
rect 2252 26793 2258 26833
rect 2252 26667 2256 26793
rect 2188 26650 2198 26658
rect 2216 26650 2224 26658
rect 2180 26642 2188 26650
rect 2196 26639 2198 26650
rect 2208 26642 2216 26650
rect 2220 26639 2222 26650
rect 2268 26639 2270 26893
rect 2272 26667 2278 26841
rect 2292 26833 2294 26953
rect 2305 26841 2308 26851
rect 2316 26841 2318 26979
rect 2354 26915 2357 26925
rect 2364 26917 2366 26979
rect 2377 26977 2382 26979
rect 2386 26953 2393 26979
rect 2364 26893 2368 26917
rect 2297 26833 2305 26841
rect 2315 26833 2318 26841
rect 2279 26793 2288 26833
rect 2290 26793 2295 26833
rect 2299 26793 2305 26833
rect 2306 26793 2322 26833
rect 2290 26785 2297 26793
rect 2316 26785 2322 26793
rect 2292 26658 2294 26785
rect 2316 26658 2318 26785
rect 2326 26667 2332 26841
rect 2336 26833 2342 26841
rect 2348 26793 2354 26833
rect 2348 26667 2352 26793
rect 2284 26650 2294 26658
rect 2312 26650 2320 26658
rect 2276 26642 2284 26650
rect 2292 26639 2294 26650
rect 2304 26642 2312 26650
rect 2316 26639 2318 26650
rect 2364 26639 2366 26893
rect 2368 26667 2374 26841
rect 2388 26833 2390 26953
rect 2401 26841 2404 26851
rect 2412 26841 2414 26979
rect 2450 26915 2453 26925
rect 2460 26917 2462 26979
rect 2473 26977 2478 26979
rect 2482 26953 2489 26979
rect 2460 26893 2464 26917
rect 2393 26833 2401 26841
rect 2411 26833 2414 26841
rect 2375 26793 2384 26833
rect 2386 26793 2391 26833
rect 2395 26793 2401 26833
rect 2402 26793 2418 26833
rect 2386 26785 2393 26793
rect 2412 26785 2418 26793
rect 2388 26658 2390 26785
rect 2412 26658 2414 26785
rect 2422 26667 2428 26841
rect 2432 26833 2438 26841
rect 2444 26793 2450 26833
rect 2444 26667 2448 26793
rect 2380 26650 2390 26658
rect 2408 26650 2416 26658
rect 2372 26642 2380 26650
rect 2388 26639 2390 26650
rect 2400 26642 2408 26650
rect 2412 26639 2414 26650
rect 2460 26639 2462 26893
rect 2464 26667 2470 26841
rect 2484 26833 2486 26953
rect 2497 26841 2500 26851
rect 2508 26841 2510 26979
rect 2546 26915 2549 26925
rect 2556 26917 2558 26979
rect 2569 26977 2574 26979
rect 2578 26953 2585 26979
rect 2556 26893 2560 26917
rect 2489 26833 2497 26841
rect 2507 26833 2510 26841
rect 2471 26793 2480 26833
rect 2482 26793 2487 26833
rect 2491 26793 2497 26833
rect 2498 26793 2514 26833
rect 2482 26785 2489 26793
rect 2508 26785 2514 26793
rect 2484 26658 2486 26785
rect 2508 26658 2510 26785
rect 2518 26667 2524 26841
rect 2528 26833 2534 26841
rect 2540 26793 2546 26833
rect 2540 26667 2544 26793
rect 2476 26650 2486 26658
rect 2504 26650 2512 26658
rect 2468 26642 2476 26650
rect 2484 26639 2486 26650
rect 2496 26642 2504 26650
rect 2508 26639 2510 26650
rect 2556 26639 2558 26893
rect 2560 26667 2566 26841
rect 2580 26833 2582 26953
rect 2593 26841 2596 26851
rect 2604 26841 2606 26979
rect 2642 26915 2645 26925
rect 2652 26917 2654 26979
rect 2665 26977 2670 26979
rect 2674 26953 2681 26979
rect 2652 26893 2656 26917
rect 2585 26833 2593 26841
rect 2603 26833 2606 26841
rect 2567 26793 2576 26833
rect 2578 26793 2583 26833
rect 2587 26793 2593 26833
rect 2594 26793 2610 26833
rect 2578 26785 2585 26793
rect 2604 26785 2610 26793
rect 2580 26658 2582 26785
rect 2604 26658 2606 26785
rect 2614 26667 2620 26841
rect 2624 26833 2630 26841
rect 2636 26793 2642 26833
rect 2636 26667 2640 26793
rect 2572 26650 2582 26658
rect 2600 26650 2608 26658
rect 2564 26642 2572 26650
rect 2580 26639 2582 26650
rect 2592 26642 2600 26650
rect 2604 26639 2606 26650
rect 2652 26639 2654 26893
rect 2656 26667 2662 26841
rect 2676 26833 2678 26953
rect 2689 26841 2692 26851
rect 2700 26841 2702 26979
rect 2738 26915 2741 26925
rect 2748 26917 2750 26979
rect 2761 26977 2766 26979
rect 2770 26953 2777 26979
rect 2748 26893 2752 26917
rect 2681 26833 2689 26841
rect 2699 26833 2702 26841
rect 2663 26793 2672 26833
rect 2674 26793 2679 26833
rect 2683 26793 2689 26833
rect 2690 26793 2706 26833
rect 2674 26785 2681 26793
rect 2700 26785 2706 26793
rect 2676 26658 2678 26785
rect 2700 26658 2702 26785
rect 2710 26667 2716 26841
rect 2720 26833 2726 26841
rect 2732 26793 2738 26833
rect 2732 26667 2736 26793
rect 2668 26650 2678 26658
rect 2696 26650 2704 26658
rect 2660 26642 2668 26650
rect 2676 26639 2678 26650
rect 2688 26642 2696 26650
rect 2700 26639 2702 26650
rect 2748 26639 2750 26893
rect 2752 26667 2758 26841
rect 2772 26833 2774 26953
rect 2785 26841 2788 26851
rect 2796 26841 2798 26979
rect 2841 26917 2847 26979
rect 2860 26969 2863 26979
rect 2868 26969 2872 26979
rect 2868 26953 2871 26969
rect 2831 26907 2836 26913
rect 2831 26903 2838 26907
rect 2841 26893 2848 26917
rect 2841 26889 2846 26893
rect 2844 26841 2846 26889
rect 2860 26891 2863 26953
rect 2860 26889 2865 26891
rect 2860 26851 2863 26889
rect 2868 26851 2870 26953
rect 2857 26841 2870 26851
rect 2777 26833 2785 26841
rect 2795 26833 2798 26841
rect 2759 26793 2768 26833
rect 2770 26793 2775 26833
rect 2779 26793 2785 26833
rect 2786 26793 2802 26833
rect 2770 26785 2777 26793
rect 2796 26785 2802 26793
rect 2772 26658 2774 26785
rect 2796 26658 2798 26785
rect 2806 26667 2812 26841
rect 2816 26833 2822 26841
rect 2844 26833 2853 26841
rect 2861 26833 2870 26841
rect 2873 26841 2877 26979
rect 2887 26841 2890 26979
rect 2828 26793 2834 26833
rect 2842 26793 2853 26833
rect 2855 26793 2858 26833
rect 2860 26793 2871 26833
rect 2873 26793 2880 26841
rect 2892 26833 2894 26979
rect 2936 26978 2942 26979
rect 2929 26841 2932 26851
rect 2940 26841 2942 26978
rect 2908 26833 2912 26841
rect 2936 26833 2942 26841
rect 2962 26833 2966 26841
rect 2882 26793 2885 26833
rect 2828 26667 2832 26793
rect 2764 26650 2774 26658
rect 2792 26650 2800 26658
rect 2824 26650 2840 26658
rect 2756 26642 2764 26650
rect 2772 26639 2774 26650
rect 2784 26642 2792 26650
rect 2796 26639 2798 26650
rect 2844 26639 2846 26793
rect 2860 26785 2867 26793
rect 2868 26658 2870 26793
rect 2887 26785 2894 26833
rect 2896 26793 2898 26833
rect 2892 26658 2894 26785
rect 2918 26667 2922 26833
rect 2923 26793 2934 26833
rect 2936 26793 2943 26833
rect 2945 26793 2948 26833
rect 2950 26793 2961 26833
rect 2963 26793 2966 26833
rect 2856 26650 2870 26658
rect 2884 26650 2896 26658
rect 2916 26650 2924 26658
rect 2852 26642 2856 26650
rect 2868 26639 2870 26650
rect 2880 26642 2884 26650
rect 2892 26639 2894 26650
rect 2924 26642 2932 26650
rect 2940 26639 2942 26793
rect 2943 26785 2948 26793
rect 2972 26667 2976 26793
rect 3012 26658 3014 26979
rect 3016 26970 3017 26979
rect 3108 26969 3112 26979
rect 3017 26919 3024 26967
rect 3108 26959 3118 26969
rect 3108 26913 3110 26959
rect 3095 26911 3110 26913
rect 3095 26903 3100 26911
rect 3108 26903 3110 26911
rect 3119 26911 3134 26959
rect 3145 26953 3148 26963
rect 3156 26953 3158 26979
rect 3155 26937 3158 26953
rect 3119 26903 3128 26911
rect 3105 26889 3110 26903
rect 3043 26667 3052 26843
rect 2944 26650 2952 26658
rect 3006 26650 3016 26658
rect 3034 26650 3044 26658
rect 3066 26650 3074 26658
rect 3094 26650 3106 26658
rect 3108 26650 3110 26889
rect 3126 26839 3135 26849
rect 3136 26667 3145 26839
rect 3156 26658 3158 26937
rect 3252 26969 3254 26979
rect 3348 26969 3352 26979
rect 3252 26955 3256 26969
rect 3257 26955 3264 26967
rect 3252 26945 3264 26955
rect 3171 26895 3173 26899
rect 3181 26881 3183 26895
rect 3185 26791 3189 26849
rect 3202 26831 3206 26839
rect 3190 26791 3201 26831
rect 3203 26791 3206 26831
rect 3185 26783 3188 26791
rect 3212 26667 3216 26791
rect 3252 26658 3254 26945
rect 3256 26929 3264 26945
rect 3257 26919 3264 26929
rect 3348 26959 3358 26969
rect 3348 26913 3350 26959
rect 3335 26911 3350 26913
rect 3335 26903 3340 26911
rect 3348 26903 3350 26911
rect 3359 26911 3374 26959
rect 3385 26953 3388 26963
rect 3396 26953 3398 26979
rect 3395 26937 3398 26953
rect 3359 26903 3368 26911
rect 3345 26889 3350 26903
rect 3283 26667 3292 26841
rect 3122 26650 3134 26658
rect 3150 26650 3162 26658
rect 3182 26650 3190 26658
rect 3246 26650 3254 26658
rect 3274 26650 3282 26658
rect 3306 26650 3314 26658
rect 3334 26650 3346 26658
rect 3348 26650 3350 26889
rect 3366 26839 3375 26849
rect 3376 26667 3385 26839
rect 3396 26658 3398 26937
rect 3455 26903 3460 26913
rect 3468 26903 3470 26979
rect 3491 26977 3504 26979
rect 3491 26972 3494 26977
rect 3411 26895 3413 26899
rect 3421 26881 3423 26895
rect 3465 26889 3470 26903
rect 3425 26791 3429 26849
rect 3468 26841 3470 26889
rect 3492 26969 3494 26972
rect 3492 26945 3496 26969
rect 3442 26831 3446 26839
rect 3430 26791 3441 26831
rect 3443 26791 3446 26831
rect 3468 26791 3478 26841
rect 3486 26839 3489 26849
rect 3492 26831 3494 26945
rect 3497 26839 3504 26972
rect 3505 26953 3508 26963
rect 3516 26953 3518 26979
rect 3515 26937 3518 26953
rect 3479 26791 3485 26831
rect 3425 26783 3428 26791
rect 3452 26667 3456 26791
rect 3362 26650 3374 26658
rect 3390 26650 3402 26658
rect 3422 26650 3430 26658
rect 3450 26650 3466 26658
rect 2952 26642 2960 26650
rect 3000 26642 3006 26650
rect 3012 26639 3014 26650
rect 3028 26642 3034 26650
rect 3074 26642 3082 26650
rect 3106 26642 3110 26650
rect 3134 26642 3138 26650
rect 3108 26639 3110 26642
rect 3156 26639 3158 26650
rect 3162 26642 3166 26650
rect 3190 26642 3198 26650
rect 3238 26642 3246 26650
rect 3252 26639 3254 26650
rect 3266 26642 3274 26650
rect 3314 26642 3322 26650
rect 3346 26642 3350 26650
rect 3374 26642 3378 26650
rect 3348 26639 3350 26642
rect 3396 26639 3398 26650
rect 3402 26642 3406 26650
rect 3430 26642 3438 26650
rect 3468 26639 3470 26791
rect 3487 26783 3494 26831
rect 3496 26783 3505 26839
rect 3516 26831 3518 26937
rect 3575 26903 3580 26913
rect 3588 26903 3590 26979
rect 3611 26977 3624 26979
rect 3611 26972 3614 26977
rect 3531 26895 3533 26899
rect 3541 26881 3543 26895
rect 3585 26889 3590 26903
rect 3506 26791 3512 26831
rect 3514 26783 3521 26831
rect 3523 26791 3532 26841
rect 3545 26791 3549 26849
rect 3588 26841 3590 26889
rect 3612 26969 3614 26972
rect 3612 26945 3616 26969
rect 3562 26831 3566 26839
rect 3550 26791 3561 26831
rect 3563 26791 3566 26831
rect 3588 26791 3598 26841
rect 3606 26839 3609 26849
rect 3612 26831 3614 26945
rect 3617 26839 3624 26972
rect 3625 26953 3628 26963
rect 3636 26953 3638 26979
rect 3635 26937 3638 26953
rect 3599 26791 3605 26831
rect 3545 26783 3548 26791
rect 3492 26658 3494 26783
rect 3516 26658 3518 26783
rect 3572 26667 3576 26791
rect 3482 26650 3494 26658
rect 3510 26650 3522 26658
rect 3542 26650 3550 26658
rect 3570 26650 3586 26658
rect 3478 26642 3482 26650
rect 3492 26639 3494 26650
rect 3506 26642 3510 26650
rect 3516 26639 3518 26650
rect 3550 26642 3558 26650
rect 3588 26639 3590 26791
rect 3607 26783 3614 26831
rect 3616 26783 3625 26839
rect 3636 26831 3638 26937
rect 3651 26895 3653 26899
rect 3661 26881 3663 26895
rect 3626 26791 3632 26831
rect 3634 26783 3641 26831
rect 3643 26791 3652 26841
rect 3665 26791 3669 26849
rect 3682 26831 3686 26839
rect 3670 26791 3681 26831
rect 3683 26791 3686 26831
rect 3665 26783 3668 26791
rect 3612 26658 3614 26783
rect 3636 26658 3638 26783
rect 3692 26667 3696 26791
rect 3602 26650 3614 26658
rect 3630 26650 3642 26658
rect 3662 26650 3670 26658
rect 3598 26642 3602 26650
rect 3612 26639 3614 26650
rect 3626 26642 3630 26650
rect 3636 26639 3638 26650
rect 3670 26642 3678 26650
rect 3708 26639 3710 26979
rect 3732 26977 3746 26979
rect 3732 26969 3734 26977
rect 3731 26961 3736 26969
rect 3732 26955 3736 26961
rect 3730 26929 3737 26955
rect 3712 26667 3718 26841
rect 3732 26831 3734 26929
rect 3745 26841 3748 26851
rect 3756 26841 3758 26979
rect 3794 26915 3797 26925
rect 3804 26917 3806 26979
rect 3817 26977 3822 26979
rect 3826 26953 3833 26979
rect 3804 26893 3808 26917
rect 3737 26831 3745 26841
rect 3755 26831 3758 26841
rect 3719 26793 3728 26831
rect 3730 26793 3735 26831
rect 3739 26793 3745 26831
rect 3746 26793 3762 26831
rect 3730 26785 3737 26793
rect 3756 26785 3762 26793
rect 3732 26658 3734 26785
rect 3756 26658 3758 26785
rect 3766 26667 3772 26841
rect 3776 26833 3782 26841
rect 3788 26793 3794 26833
rect 3788 26667 3792 26793
rect 3724 26650 3734 26658
rect 3752 26650 3762 26658
rect 3718 26642 3724 26650
rect 3732 26639 3734 26650
rect 3746 26642 3752 26650
rect 3756 26639 3758 26650
rect 3804 26639 3806 26893
rect 3808 26667 3814 26841
rect 3828 26833 3830 26953
rect 3841 26841 3844 26851
rect 3852 26841 3854 26979
rect 3890 26915 3893 26925
rect 3900 26917 3902 26979
rect 3913 26977 3918 26979
rect 3922 26953 3929 26979
rect 3900 26893 3904 26917
rect 3833 26833 3841 26841
rect 3851 26833 3854 26841
rect 3815 26793 3824 26833
rect 3826 26793 3831 26833
rect 3835 26793 3841 26833
rect 3842 26793 3858 26833
rect 3826 26785 3833 26793
rect 3852 26785 3858 26793
rect 3828 26658 3830 26785
rect 3852 26658 3854 26785
rect 3862 26667 3868 26841
rect 3872 26833 3878 26841
rect 3884 26793 3890 26833
rect 3884 26667 3888 26793
rect 3820 26650 3830 26658
rect 3848 26650 3856 26658
rect 3812 26642 3820 26650
rect 3828 26639 3830 26650
rect 3840 26642 3848 26650
rect 3852 26639 3854 26650
rect 3900 26639 3902 26893
rect 3904 26667 3910 26841
rect 3924 26833 3926 26953
rect 3937 26841 3940 26851
rect 3948 26841 3950 26979
rect 3986 26915 3989 26925
rect 3996 26917 3998 26979
rect 4009 26977 4014 26979
rect 4018 26953 4025 26979
rect 3996 26893 4000 26917
rect 3929 26833 3937 26841
rect 3947 26833 3950 26841
rect 3911 26793 3920 26833
rect 3922 26793 3927 26833
rect 3931 26793 3937 26833
rect 3938 26793 3954 26833
rect 3922 26785 3929 26793
rect 3948 26785 3954 26793
rect 3924 26658 3926 26785
rect 3948 26658 3950 26785
rect 3958 26667 3964 26841
rect 3968 26833 3974 26841
rect 3980 26793 3986 26833
rect 3980 26667 3984 26793
rect 3916 26650 3926 26658
rect 3944 26650 3952 26658
rect 3908 26642 3916 26650
rect 3924 26639 3926 26650
rect 3936 26642 3944 26650
rect 3948 26639 3950 26650
rect 3996 26639 3998 26893
rect 4000 26667 4006 26841
rect 4020 26833 4022 26953
rect 4033 26841 4036 26851
rect 4044 26841 4046 26979
rect 4082 26915 4085 26925
rect 4092 26917 4094 26979
rect 4105 26977 4110 26979
rect 4114 26953 4121 26979
rect 4092 26893 4096 26917
rect 4025 26833 4033 26841
rect 4043 26833 4046 26841
rect 4007 26793 4016 26833
rect 4018 26793 4023 26833
rect 4027 26793 4033 26833
rect 4034 26793 4050 26833
rect 4018 26785 4025 26793
rect 4044 26785 4050 26793
rect 4020 26658 4022 26785
rect 4044 26658 4046 26785
rect 4054 26667 4060 26841
rect 4064 26833 4070 26841
rect 4076 26793 4082 26833
rect 4076 26667 4080 26793
rect 4012 26650 4022 26658
rect 4040 26650 4048 26658
rect 4004 26642 4012 26650
rect 4020 26639 4022 26650
rect 4032 26642 4040 26650
rect 4044 26639 4046 26650
rect 4092 26639 4094 26893
rect 4096 26667 4102 26841
rect 4116 26833 4118 26953
rect 4129 26841 4132 26851
rect 4140 26841 4142 26979
rect 4178 26915 4181 26925
rect 4188 26917 4190 26979
rect 4201 26977 4206 26979
rect 4210 26953 4217 26979
rect 4188 26893 4192 26917
rect 4121 26833 4129 26841
rect 4139 26833 4142 26841
rect 4103 26793 4112 26833
rect 4114 26793 4119 26833
rect 4123 26793 4129 26833
rect 4130 26793 4146 26833
rect 4114 26785 4121 26793
rect 4140 26785 4146 26793
rect 4116 26658 4118 26785
rect 4140 26658 4142 26785
rect 4150 26667 4156 26841
rect 4160 26833 4166 26841
rect 4172 26793 4178 26833
rect 4172 26667 4176 26793
rect 4108 26650 4118 26658
rect 4136 26650 4144 26658
rect 4100 26642 4108 26650
rect 4116 26639 4118 26650
rect 4128 26642 4136 26650
rect 4140 26639 4142 26650
rect 4188 26639 4190 26893
rect 4192 26667 4198 26841
rect 4212 26833 4214 26953
rect 4225 26841 4228 26851
rect 4236 26841 4238 26979
rect 4274 26915 4277 26925
rect 4284 26917 4286 26979
rect 4297 26977 4302 26979
rect 4306 26953 4313 26979
rect 4284 26893 4288 26917
rect 4217 26833 4225 26841
rect 4235 26833 4238 26841
rect 4199 26793 4208 26833
rect 4210 26793 4215 26833
rect 4219 26793 4225 26833
rect 4226 26793 4242 26833
rect 4210 26785 4217 26793
rect 4236 26785 4242 26793
rect 4212 26658 4214 26785
rect 4236 26658 4238 26785
rect 4246 26667 4252 26841
rect 4256 26833 4262 26841
rect 4268 26793 4274 26833
rect 4268 26667 4272 26793
rect 4204 26650 4214 26658
rect 4232 26650 4240 26658
rect 4196 26642 4204 26650
rect 4212 26639 4214 26650
rect 4224 26642 4232 26650
rect 4236 26639 4238 26650
rect 4284 26639 4286 26893
rect 4288 26667 4294 26841
rect 4308 26833 4310 26953
rect 4321 26841 4324 26851
rect 4332 26841 4334 26979
rect 4370 26915 4373 26925
rect 4380 26917 4382 26979
rect 4393 26977 4398 26979
rect 4402 26953 4409 26979
rect 4380 26893 4384 26917
rect 4313 26833 4321 26841
rect 4331 26833 4334 26841
rect 4295 26793 4304 26833
rect 4306 26793 4311 26833
rect 4315 26793 4321 26833
rect 4322 26793 4338 26833
rect 4306 26785 4313 26793
rect 4332 26785 4338 26793
rect 4308 26658 4310 26785
rect 4332 26658 4334 26785
rect 4342 26667 4348 26841
rect 4352 26833 4358 26841
rect 4364 26793 4370 26833
rect 4364 26667 4368 26793
rect 4300 26650 4310 26658
rect 4328 26650 4336 26658
rect 4292 26642 4300 26650
rect 4308 26639 4310 26650
rect 4320 26642 4328 26650
rect 4332 26639 4334 26650
rect 4380 26639 4382 26893
rect 4384 26667 4390 26841
rect 4404 26833 4406 26953
rect 4417 26841 4420 26851
rect 4428 26841 4430 26979
rect 4466 26915 4469 26925
rect 4476 26917 4478 26979
rect 4489 26977 4494 26979
rect 4498 26953 4505 26979
rect 4476 26893 4480 26917
rect 4409 26833 4417 26841
rect 4427 26833 4430 26841
rect 4391 26793 4400 26833
rect 4402 26793 4407 26833
rect 4411 26793 4417 26833
rect 4418 26793 4434 26833
rect 4402 26785 4409 26793
rect 4428 26785 4434 26793
rect 4404 26658 4406 26785
rect 4428 26658 4430 26785
rect 4438 26667 4444 26841
rect 4448 26833 4454 26841
rect 4460 26793 4466 26833
rect 4460 26667 4464 26793
rect 4396 26650 4406 26658
rect 4424 26650 4432 26658
rect 4388 26642 4396 26650
rect 4404 26639 4406 26650
rect 4416 26642 4424 26650
rect 4428 26639 4430 26650
rect 4476 26639 4478 26893
rect 4480 26667 4486 26841
rect 4500 26833 4502 26953
rect 4513 26841 4516 26851
rect 4524 26841 4526 26979
rect 4596 26969 4601 26979
rect 4809 26969 4816 26979
rect 4596 26953 4599 26969
rect 4600 26967 4601 26969
rect 4720 26967 4729 26969
rect 4600 26953 4608 26967
rect 4505 26833 4513 26841
rect 4523 26833 4526 26841
rect 4487 26793 4496 26833
rect 4498 26793 4503 26833
rect 4507 26793 4513 26833
rect 4514 26793 4530 26833
rect 4498 26785 4505 26793
rect 4524 26785 4530 26793
rect 4500 26658 4502 26785
rect 4524 26658 4526 26785
rect 4534 26667 4540 26841
rect 4544 26833 4550 26841
rect 4556 26793 4562 26833
rect 4556 26667 4560 26793
rect 4596 26658 4598 26953
rect 4601 26919 4608 26953
rect 4720 26919 4731 26967
rect 4809 26959 4819 26969
rect 4828 26959 4831 26979
rect 4799 26903 4804 26913
rect 4812 26903 4814 26959
rect 4823 26911 4835 26959
rect 4823 26903 4831 26911
rect 4809 26889 4814 26903
rect 4627 26667 4636 26843
rect 4492 26650 4502 26658
rect 4520 26650 4528 26658
rect 4590 26650 4598 26658
rect 4618 26650 4624 26658
rect 4650 26650 4658 26658
rect 4678 26650 4694 26658
rect 4710 26650 4722 26658
rect 4738 26650 4750 26658
rect 4770 26650 4778 26658
rect 4798 26650 4808 26658
rect 4812 26650 4814 26889
rect 4860 26658 4862 26979
rect 4904 26978 4910 26979
rect 4897 26841 4900 26851
rect 4908 26841 4910 26978
rect 4943 26903 4948 26913
rect 4956 26903 4958 26979
rect 4976 26972 4985 26979
rect 4953 26889 4958 26903
rect 4956 26843 4958 26889
rect 4876 26833 4880 26841
rect 4904 26833 4910 26841
rect 4930 26833 4934 26841
rect 4886 26667 4890 26833
rect 4891 26793 4902 26833
rect 4904 26793 4911 26833
rect 4913 26793 4916 26833
rect 4918 26793 4929 26833
rect 4931 26793 4934 26833
rect 4826 26650 4836 26658
rect 4854 26650 4864 26658
rect 4884 26650 4892 26658
rect 4484 26642 4492 26650
rect 4500 26639 4502 26650
rect 4512 26642 4520 26650
rect 4524 26639 4526 26650
rect 4580 26642 4590 26650
rect 4596 26639 4598 26650
rect 4608 26642 4618 26650
rect 4658 26642 4666 26650
rect 4706 26642 4710 26650
rect 4734 26642 4738 26650
rect 4778 26642 4786 26650
rect 4808 26642 4814 26650
rect 4836 26642 4842 26650
rect 4812 26639 4814 26642
rect 4860 26639 4862 26650
rect 4864 26642 4870 26650
rect 4892 26642 4900 26650
rect 4908 26639 4910 26793
rect 4911 26785 4916 26793
rect 4940 26667 4944 26793
rect 4956 26791 4966 26843
rect 4974 26839 4977 26849
rect 4980 26833 4982 26972
rect 4985 26839 4992 26972
rect 4993 26953 4996 26963
rect 5004 26953 5006 26979
rect 5003 26937 5006 26953
rect 4967 26791 4973 26833
rect 4912 26650 4920 26658
rect 4940 26650 4954 26658
rect 4956 26650 4958 26791
rect 4975 26785 4982 26833
rect 4984 26785 4993 26839
rect 5004 26833 5006 26937
rect 5019 26895 5021 26899
rect 5029 26881 5031 26895
rect 4994 26791 5000 26833
rect 5002 26785 5009 26833
rect 5011 26791 5020 26843
rect 5033 26791 5037 26849
rect 5050 26831 5054 26839
rect 5038 26791 5049 26831
rect 5051 26791 5054 26831
rect 4980 26658 4982 26785
rect 4985 26783 4992 26785
rect 5004 26658 5006 26785
rect 5033 26783 5036 26791
rect 5060 26667 5064 26791
rect 4970 26650 4982 26658
rect 4998 26650 5010 26658
rect 5030 26650 5038 26658
rect 4920 26642 4928 26650
rect 4954 26642 4958 26650
rect 4968 26642 4970 26650
rect 4980 26642 4984 26650
rect 4996 26642 4998 26650
rect 4956 26639 4958 26642
rect 4980 26639 4982 26642
rect 5004 26639 5006 26650
rect 5010 26642 5012 26650
rect 5038 26642 5046 26650
rect 5076 26639 5078 26979
rect 5100 26977 5114 26979
rect 5100 26969 5102 26977
rect 5099 26961 5104 26969
rect 5100 26955 5104 26961
rect 5098 26929 5105 26955
rect 5080 26667 5086 26841
rect 5100 26831 5102 26929
rect 5113 26841 5116 26851
rect 5124 26841 5126 26979
rect 5162 26915 5165 26925
rect 5172 26917 5174 26979
rect 5185 26977 5190 26979
rect 5194 26953 5201 26979
rect 5172 26893 5176 26917
rect 5105 26831 5113 26841
rect 5123 26831 5126 26841
rect 5087 26793 5096 26831
rect 5098 26793 5103 26831
rect 5107 26793 5113 26831
rect 5114 26793 5130 26831
rect 5098 26785 5105 26793
rect 5124 26785 5130 26793
rect 5100 26658 5102 26785
rect 5124 26658 5126 26785
rect 5134 26667 5140 26841
rect 5144 26833 5150 26841
rect 5156 26793 5162 26833
rect 5156 26667 5160 26793
rect 5092 26650 5102 26658
rect 5120 26650 5130 26658
rect 5086 26642 5092 26650
rect 5100 26639 5102 26650
rect 5114 26642 5120 26650
rect 5124 26639 5126 26650
rect 5172 26639 5174 26893
rect 5176 26667 5182 26841
rect 5196 26833 5198 26953
rect 5209 26841 5212 26851
rect 5220 26841 5222 26979
rect 5268 26917 5271 26979
rect 5288 26972 5297 26979
rect 5292 26969 5296 26972
rect 5292 26953 5295 26969
rect 5255 26907 5260 26913
rect 5255 26903 5262 26907
rect 5268 26903 5272 26917
rect 5265 26893 5272 26903
rect 5265 26889 5270 26893
rect 5268 26843 5270 26889
rect 5285 26849 5289 26889
rect 5292 26849 5294 26953
rect 5201 26833 5209 26841
rect 5219 26833 5222 26841
rect 5183 26793 5192 26833
rect 5194 26793 5199 26833
rect 5203 26793 5209 26833
rect 5210 26793 5226 26833
rect 5194 26785 5201 26793
rect 5220 26785 5226 26793
rect 5196 26658 5198 26785
rect 5220 26658 5222 26785
rect 5230 26667 5236 26841
rect 5240 26833 5246 26841
rect 5252 26793 5258 26833
rect 5252 26667 5256 26793
rect 5268 26791 5278 26843
rect 5285 26839 5295 26849
rect 5297 26839 5304 26972
rect 5305 26953 5308 26963
rect 5316 26953 5318 26979
rect 5315 26937 5318 26953
rect 5292 26833 5294 26839
rect 5279 26791 5285 26833
rect 5188 26650 5198 26658
rect 5216 26650 5224 26658
rect 5180 26642 5188 26650
rect 5196 26639 5198 26650
rect 5208 26642 5216 26650
rect 5220 26639 5222 26650
rect 5268 26639 5270 26791
rect 5287 26785 5294 26833
rect 5296 26785 5305 26839
rect 5316 26833 5318 26937
rect 5331 26895 5333 26899
rect 5341 26881 5343 26895
rect 5306 26791 5312 26833
rect 5314 26785 5321 26833
rect 5323 26791 5332 26843
rect 5345 26791 5349 26849
rect 5362 26831 5366 26839
rect 5350 26791 5361 26831
rect 5363 26791 5366 26831
rect 5292 26658 5294 26785
rect 5297 26783 5304 26785
rect 5316 26658 5318 26785
rect 5345 26783 5348 26791
rect 5372 26667 5376 26791
rect 5282 26650 5294 26658
rect 5310 26650 5320 26658
rect 5342 26650 5350 26658
rect 5276 26642 5282 26650
rect 5292 26639 5294 26650
rect 5304 26642 5310 26650
rect 5316 26639 5318 26650
rect 5350 26642 5358 26650
rect 5388 26639 5390 26979
rect 5412 26977 5426 26979
rect 5412 26969 5414 26977
rect 5411 26961 5416 26969
rect 5412 26955 5416 26961
rect 5410 26929 5417 26955
rect 5392 26667 5398 26841
rect 5412 26831 5414 26929
rect 5425 26841 5428 26851
rect 5436 26841 5438 26979
rect 5474 26915 5477 26925
rect 5484 26917 5486 26979
rect 5497 26977 5502 26979
rect 5506 26953 5513 26979
rect 5484 26893 5488 26917
rect 5417 26831 5425 26841
rect 5435 26831 5438 26841
rect 5399 26793 5408 26831
rect 5410 26793 5415 26831
rect 5419 26793 5425 26831
rect 5426 26793 5442 26831
rect 5410 26785 5417 26793
rect 5436 26785 5442 26793
rect 5412 26658 5414 26785
rect 5436 26658 5438 26785
rect 5446 26667 5452 26841
rect 5456 26833 5462 26841
rect 5468 26793 5474 26833
rect 5468 26667 5472 26793
rect 5404 26650 5414 26658
rect 5432 26650 5442 26658
rect 5398 26642 5404 26650
rect 5412 26639 5414 26650
rect 5426 26642 5432 26650
rect 5436 26639 5438 26650
rect 5484 26639 5486 26893
rect 5488 26667 5494 26841
rect 5508 26833 5510 26953
rect 5521 26841 5524 26851
rect 5532 26841 5534 26979
rect 5580 26917 5582 26979
rect 5583 26953 5599 26964
rect 5583 26917 5589 26953
rect 5580 26916 5589 26917
rect 5609 26916 5611 26964
rect 5580 26893 5584 26916
rect 5513 26833 5521 26841
rect 5531 26833 5534 26841
rect 5495 26793 5504 26833
rect 5506 26793 5511 26833
rect 5515 26793 5521 26833
rect 5522 26793 5538 26833
rect 5506 26785 5513 26793
rect 5532 26785 5538 26793
rect 5508 26658 5510 26785
rect 5532 26658 5534 26785
rect 5542 26667 5548 26841
rect 5552 26833 5558 26841
rect 5564 26793 5570 26833
rect 5564 26667 5568 26793
rect 5500 26650 5510 26658
rect 5528 26650 5536 26658
rect 5492 26642 5500 26650
rect 5508 26639 5510 26650
rect 5520 26642 5528 26650
rect 5532 26639 5534 26650
rect 5580 26639 5582 26893
rect 5628 26658 5630 26979
rect 5722 26977 5729 26979
rect 5722 26966 5731 26977
rect 5722 26961 5739 26966
rect 5659 26916 5671 26956
rect 5722 26900 5729 26961
rect 5744 26908 5747 26956
rect 5724 26851 5726 26900
rect 5723 26667 5730 26851
rect 5737 26841 5740 26851
rect 5748 26841 5750 26979
rect 5786 26915 5789 26925
rect 5796 26917 5798 26979
rect 5809 26977 5814 26979
rect 5818 26953 5825 26979
rect 5796 26893 5800 26917
rect 5747 26793 5750 26841
rect 5768 26833 5774 26841
rect 5724 26658 5726 26667
rect 5748 26658 5750 26793
rect 5780 26793 5786 26833
rect 5780 26667 5784 26793
rect 5594 26650 5604 26658
rect 5622 26650 5632 26658
rect 5654 26650 5662 26658
rect 5716 26650 5726 26658
rect 5744 26650 5754 26658
rect 5588 26642 5594 26650
rect 5616 26642 5622 26650
rect 5628 26639 5630 26650
rect 5662 26642 5670 26650
rect 5710 26642 5716 26650
rect 5724 26639 5726 26650
rect 5738 26642 5744 26650
rect 5748 26639 5750 26650
rect 5796 26639 5798 26893
rect 5800 26667 5806 26841
rect 5820 26833 5822 26953
rect 5833 26841 5836 26851
rect 5844 26841 5846 26979
rect 5916 26969 5921 26979
rect 5916 26953 5919 26969
rect 5920 26967 5921 26969
rect 6040 26967 6049 26969
rect 5920 26953 5928 26967
rect 5825 26833 5833 26841
rect 5843 26833 5846 26841
rect 5807 26793 5816 26833
rect 5818 26793 5823 26833
rect 5827 26793 5833 26833
rect 5834 26793 5850 26833
rect 5818 26785 5825 26793
rect 5844 26785 5850 26793
rect 5820 26658 5822 26785
rect 5844 26658 5846 26785
rect 5854 26667 5860 26841
rect 5864 26833 5870 26841
rect 5876 26793 5882 26833
rect 5876 26667 5880 26793
rect 5916 26658 5918 26953
rect 5921 26919 5928 26953
rect 6040 26919 6051 26967
rect 6132 26921 6134 26979
rect 6135 26969 6136 26979
rect 6135 26921 6142 26969
rect 6155 26961 6169 26969
rect 6132 26915 6142 26921
rect 5947 26667 5956 26843
rect 6132 26658 6134 26915
rect 6143 26911 6146 26915
rect 6154 26911 6159 26959
rect 6153 26841 6159 26851
rect 6169 26841 6172 26851
rect 6180 26841 6182 26979
rect 6218 26915 6221 26925
rect 6228 26917 6230 26979
rect 6241 26977 6246 26979
rect 6250 26953 6257 26979
rect 6228 26893 6232 26917
rect 6163 26793 6169 26841
rect 6179 26793 6182 26841
rect 6200 26833 6206 26841
rect 6180 26658 6182 26793
rect 6212 26793 6218 26833
rect 6212 26667 6216 26793
rect 5812 26650 5822 26658
rect 5840 26650 5848 26658
rect 5910 26650 5918 26658
rect 5938 26650 5944 26658
rect 5970 26650 5978 26658
rect 5998 26650 6014 26658
rect 6030 26650 6042 26658
rect 6058 26650 6070 26658
rect 6090 26650 6098 26658
rect 6118 26650 6134 26658
rect 6148 26650 6160 26658
rect 6176 26650 6188 26658
rect 5804 26642 5812 26650
rect 5820 26639 5822 26650
rect 5832 26642 5840 26650
rect 5844 26639 5846 26650
rect 5900 26642 5910 26650
rect 5916 26639 5918 26650
rect 5928 26642 5938 26650
rect 5978 26642 5986 26650
rect 6026 26642 6030 26650
rect 6054 26642 6058 26650
rect 6098 26642 6106 26650
rect 6132 26639 6134 26650
rect 6146 26642 6148 26650
rect 6160 26642 6162 26650
rect 6174 26642 6176 26650
rect 6180 26639 6182 26650
rect 6188 26642 6190 26650
rect 6228 26639 6230 26893
rect 6232 26667 6238 26841
rect 6252 26833 6254 26953
rect 6265 26841 6268 26851
rect 6276 26841 6278 26979
rect 6324 26917 6326 26979
rect 6327 26953 6343 26964
rect 6327 26917 6333 26953
rect 6324 26916 6333 26917
rect 6353 26916 6355 26964
rect 6324 26893 6328 26916
rect 6257 26833 6265 26841
rect 6275 26833 6278 26841
rect 6239 26793 6248 26833
rect 6250 26793 6255 26833
rect 6259 26793 6265 26833
rect 6266 26793 6282 26833
rect 6250 26785 6257 26793
rect 6276 26785 6282 26793
rect 6252 26658 6254 26785
rect 6276 26658 6278 26785
rect 6286 26667 6292 26841
rect 6296 26833 6302 26841
rect 6308 26793 6314 26833
rect 6308 26667 6312 26793
rect 6244 26650 6254 26658
rect 6272 26650 6280 26658
rect 6236 26642 6244 26650
rect 6252 26639 6254 26650
rect 6264 26642 6272 26650
rect 6276 26639 6278 26650
rect 6324 26639 6326 26893
rect 6372 26658 6374 26979
rect 6467 26972 6470 26979
rect 6468 26956 6470 26972
rect 6492 26966 6494 26979
rect 6403 26916 6415 26956
rect 6465 26908 6470 26956
rect 6481 26953 6484 26963
rect 6490 26953 6491 26956
rect 6492 26953 6501 26966
rect 6490 26937 6494 26953
rect 6490 26908 6491 26937
rect 6468 26849 6470 26908
rect 6467 26791 6471 26849
rect 6468 26658 6470 26791
rect 6492 26658 6494 26937
rect 6507 26895 6509 26899
rect 6499 26791 6501 26889
rect 6517 26881 6519 26895
rect 6521 26791 6525 26849
rect 6538 26831 6542 26839
rect 6526 26791 6537 26831
rect 6539 26791 6542 26831
rect 6521 26783 6524 26791
rect 6548 26667 6552 26791
rect 6338 26650 6348 26658
rect 6366 26650 6376 26658
rect 6398 26650 6406 26658
rect 6426 26650 6442 26658
rect 6458 26650 6470 26658
rect 6486 26650 6498 26658
rect 6518 26650 6526 26658
rect 6332 26642 6338 26650
rect 6360 26642 6366 26650
rect 6372 26639 6374 26650
rect 6406 26642 6414 26650
rect 6454 26642 6458 26650
rect 6468 26639 6470 26650
rect 6482 26642 6486 26650
rect 6492 26639 6494 26650
rect 6526 26642 6534 26650
rect 6564 26639 6566 26979
rect 6588 26977 6602 26979
rect 6588 26969 6590 26977
rect 6587 26961 6592 26969
rect 6588 26955 6592 26961
rect 6586 26929 6593 26955
rect 6568 26667 6574 26841
rect 6588 26831 6590 26929
rect 6601 26841 6604 26851
rect 6612 26841 6614 26979
rect 6660 26917 6663 26979
rect 6680 26972 6689 26979
rect 6684 26969 6688 26972
rect 6684 26953 6687 26969
rect 6647 26907 6652 26913
rect 6647 26903 6654 26907
rect 6660 26903 6664 26917
rect 6657 26893 6664 26903
rect 6657 26889 6662 26893
rect 6660 26843 6662 26889
rect 6677 26849 6681 26889
rect 6684 26849 6686 26953
rect 6593 26831 6601 26841
rect 6611 26831 6614 26841
rect 6575 26793 6584 26831
rect 6586 26793 6591 26831
rect 6595 26793 6601 26831
rect 6602 26793 6618 26831
rect 6586 26785 6593 26793
rect 6612 26785 6618 26793
rect 6588 26658 6590 26785
rect 6612 26658 6614 26785
rect 6622 26667 6628 26841
rect 6632 26833 6638 26841
rect 6644 26793 6650 26833
rect 6644 26667 6648 26793
rect 6660 26791 6670 26843
rect 6677 26839 6687 26849
rect 6689 26839 6696 26972
rect 6697 26953 6700 26963
rect 6708 26953 6710 26979
rect 6707 26937 6710 26953
rect 6684 26833 6686 26839
rect 6671 26791 6677 26833
rect 6580 26650 6590 26658
rect 6608 26650 6618 26658
rect 6574 26642 6580 26650
rect 6588 26639 6590 26650
rect 6602 26642 6608 26650
rect 6612 26639 6614 26650
rect 6660 26639 6662 26791
rect 6679 26785 6686 26833
rect 6688 26785 6697 26839
rect 6708 26833 6710 26937
rect 6723 26895 6725 26899
rect 6733 26881 6735 26895
rect 6698 26791 6704 26833
rect 6706 26785 6713 26833
rect 6715 26791 6724 26843
rect 6737 26791 6741 26849
rect 6754 26831 6758 26839
rect 6742 26791 6753 26831
rect 6755 26791 6758 26831
rect 6684 26658 6686 26785
rect 6689 26783 6696 26785
rect 6708 26658 6710 26785
rect 6737 26783 6740 26791
rect 6764 26667 6768 26791
rect 6674 26650 6686 26658
rect 6702 26650 6712 26658
rect 6734 26650 6742 26658
rect 6668 26642 6674 26650
rect 6684 26639 6686 26650
rect 6696 26642 6702 26650
rect 6708 26639 6710 26650
rect 6742 26642 6750 26650
rect 6780 26639 6782 26979
rect 6804 26977 6818 26979
rect 6804 26969 6806 26977
rect 6803 26961 6808 26969
rect 6804 26955 6808 26961
rect 6802 26929 6809 26955
rect 6784 26667 6790 26841
rect 6804 26831 6806 26929
rect 6817 26841 6820 26851
rect 6828 26841 6830 26979
rect 6866 26915 6869 26925
rect 6876 26917 6878 26979
rect 6889 26977 6894 26979
rect 6898 26953 6905 26979
rect 6876 26893 6880 26917
rect 6809 26831 6817 26841
rect 6827 26831 6830 26841
rect 6791 26793 6800 26831
rect 6802 26793 6807 26831
rect 6811 26793 6817 26831
rect 6818 26793 6834 26831
rect 6802 26785 6809 26793
rect 6828 26785 6834 26793
rect 6804 26658 6806 26785
rect 6828 26658 6830 26785
rect 6838 26667 6844 26841
rect 6848 26833 6854 26841
rect 6860 26793 6866 26833
rect 6860 26667 6864 26793
rect 6796 26650 6806 26658
rect 6824 26650 6834 26658
rect 6790 26642 6796 26650
rect 6804 26639 6806 26650
rect 6818 26642 6824 26650
rect 6828 26639 6830 26650
rect 6876 26639 6878 26893
rect 6880 26667 6886 26841
rect 6900 26833 6902 26953
rect 6913 26841 6916 26851
rect 6924 26841 6926 26979
rect 6972 26917 6974 26979
rect 6975 26953 6991 26964
rect 6975 26917 6981 26953
rect 6972 26916 6981 26917
rect 7001 26916 7003 26964
rect 6972 26893 6976 26916
rect 6905 26833 6913 26841
rect 6923 26833 6926 26841
rect 6887 26793 6896 26833
rect 6898 26793 6903 26833
rect 6907 26793 6913 26833
rect 6914 26793 6930 26833
rect 6898 26785 6905 26793
rect 6924 26785 6930 26793
rect 6900 26658 6902 26785
rect 6924 26658 6926 26785
rect 6934 26667 6940 26841
rect 6944 26833 6950 26841
rect 6956 26793 6962 26833
rect 6956 26667 6960 26793
rect 6892 26650 6902 26658
rect 6920 26650 6928 26658
rect 6884 26642 6892 26650
rect 6900 26639 6902 26650
rect 6912 26642 6920 26650
rect 6924 26639 6926 26650
rect 6972 26639 6974 26893
rect 7020 26658 7022 26979
rect 7051 26916 7063 26956
rect 7106 26916 7113 26964
rect 7115 26916 7121 26956
rect 7123 26908 7130 26956
rect 7140 26658 7142 26979
rect 7235 26972 7238 26979
rect 7236 26956 7238 26972
rect 7260 26966 7262 26979
rect 7171 26916 7183 26956
rect 7233 26908 7238 26956
rect 7249 26953 7252 26963
rect 7258 26953 7259 26956
rect 7260 26953 7269 26966
rect 7258 26937 7262 26953
rect 7258 26908 7259 26937
rect 7236 26849 7238 26908
rect 7235 26791 7239 26849
rect 7236 26658 7238 26791
rect 7260 26658 7262 26937
rect 7275 26895 7277 26899
rect 7267 26791 7269 26889
rect 7285 26881 7287 26895
rect 7289 26791 7293 26849
rect 7306 26831 7310 26839
rect 7294 26791 7305 26831
rect 7307 26791 7310 26831
rect 7289 26783 7292 26791
rect 7316 26667 7320 26791
rect 6986 26650 6996 26658
rect 7014 26650 7024 26658
rect 7046 26650 7054 26658
rect 7074 26650 7090 26658
rect 7106 26650 7118 26658
rect 7134 26650 7146 26658
rect 7166 26650 7174 26658
rect 7194 26650 7210 26658
rect 7226 26650 7238 26658
rect 7254 26650 7266 26658
rect 7286 26650 7294 26658
rect 6980 26642 6986 26650
rect 7008 26642 7014 26650
rect 7020 26639 7022 26650
rect 7054 26642 7062 26650
rect 7102 26642 7106 26650
rect 7130 26642 7134 26650
rect 7140 26639 7142 26650
rect 7174 26642 7182 26650
rect 7222 26642 7226 26650
rect 7236 26639 7238 26650
rect 7250 26642 7254 26650
rect 7260 26639 7262 26650
rect 7294 26642 7302 26650
rect 7332 26639 7334 26979
rect 7356 26977 7370 26979
rect 7356 26969 7358 26977
rect 7355 26961 7360 26969
rect 7356 26955 7360 26961
rect 7354 26929 7361 26955
rect 7336 26667 7342 26841
rect 7356 26831 7358 26929
rect 7369 26841 7372 26851
rect 7380 26841 7382 26979
rect 7418 26915 7421 26925
rect 7428 26917 7430 26979
rect 7441 26977 7446 26979
rect 7450 26953 7457 26979
rect 7428 26893 7432 26917
rect 7361 26831 7369 26841
rect 7379 26831 7382 26841
rect 7343 26793 7352 26831
rect 7354 26793 7359 26831
rect 7363 26793 7369 26831
rect 7370 26793 7386 26831
rect 7354 26785 7361 26793
rect 7380 26785 7386 26793
rect 7356 26658 7358 26785
rect 7380 26658 7382 26785
rect 7390 26667 7396 26841
rect 7400 26833 7406 26841
rect 7412 26793 7418 26833
rect 7412 26667 7416 26793
rect 7348 26650 7358 26658
rect 7376 26650 7386 26658
rect 7342 26642 7348 26650
rect 7356 26639 7358 26650
rect 7370 26642 7376 26650
rect 7380 26639 7382 26650
rect 7428 26639 7430 26893
rect 7432 26667 7438 26841
rect 7452 26833 7454 26953
rect 7465 26841 7468 26851
rect 7476 26841 7478 26979
rect 7514 26915 7517 26925
rect 7524 26917 7526 26979
rect 7537 26977 7542 26979
rect 7546 26953 7553 26979
rect 7524 26893 7528 26917
rect 7457 26833 7465 26841
rect 7475 26833 7478 26841
rect 7439 26793 7448 26833
rect 7450 26793 7455 26833
rect 7459 26793 7465 26833
rect 7466 26793 7482 26833
rect 7450 26785 7457 26793
rect 7476 26785 7482 26793
rect 7452 26658 7454 26785
rect 7476 26658 7478 26785
rect 7486 26667 7492 26841
rect 7496 26833 7502 26841
rect 7508 26793 7514 26833
rect 7508 26667 7512 26793
rect 7444 26650 7454 26658
rect 7472 26650 7480 26658
rect 7436 26642 7444 26650
rect 7452 26639 7454 26650
rect 7464 26642 7472 26650
rect 7476 26639 7478 26650
rect 7524 26639 7526 26893
rect 7528 26667 7534 26841
rect 7548 26833 7550 26953
rect 7561 26841 7564 26851
rect 7572 26841 7574 26979
rect 7610 26915 7613 26925
rect 7620 26917 7622 26979
rect 7633 26977 7638 26979
rect 7642 26953 7649 26979
rect 7620 26893 7624 26917
rect 7553 26833 7561 26841
rect 7571 26833 7574 26841
rect 7535 26793 7544 26833
rect 7546 26793 7551 26833
rect 7555 26793 7561 26833
rect 7562 26793 7578 26833
rect 7546 26785 7553 26793
rect 7572 26785 7578 26793
rect 7548 26658 7550 26785
rect 7572 26658 7574 26785
rect 7582 26667 7588 26841
rect 7592 26833 7598 26841
rect 7604 26793 7610 26833
rect 7604 26667 7608 26793
rect 7540 26650 7550 26658
rect 7568 26650 7576 26658
rect 7532 26642 7540 26650
rect 7548 26639 7550 26650
rect 7560 26642 7568 26650
rect 7572 26639 7574 26650
rect 7620 26639 7622 26893
rect 7624 26667 7630 26841
rect 7644 26833 7646 26953
rect 7657 26841 7660 26851
rect 7668 26841 7670 26979
rect 7716 26917 7719 26979
rect 7736 26972 7745 26979
rect 7740 26969 7744 26972
rect 7740 26953 7743 26969
rect 7703 26907 7708 26913
rect 7703 26903 7710 26907
rect 7716 26903 7720 26917
rect 7713 26893 7720 26903
rect 7713 26889 7718 26893
rect 7716 26843 7718 26889
rect 7733 26849 7737 26889
rect 7740 26849 7742 26953
rect 7649 26833 7657 26841
rect 7667 26833 7670 26841
rect 7631 26793 7640 26833
rect 7642 26793 7647 26833
rect 7651 26793 7657 26833
rect 7658 26793 7674 26833
rect 7642 26785 7649 26793
rect 7668 26785 7674 26793
rect 7644 26658 7646 26785
rect 7668 26658 7670 26785
rect 7678 26667 7684 26841
rect 7688 26833 7694 26841
rect 7700 26793 7706 26833
rect 7700 26667 7704 26793
rect 7716 26791 7726 26843
rect 7733 26839 7743 26849
rect 7745 26839 7752 26972
rect 7753 26953 7756 26963
rect 7764 26953 7766 26979
rect 7763 26937 7766 26953
rect 7740 26833 7742 26839
rect 7727 26791 7733 26833
rect 7636 26650 7646 26658
rect 7664 26650 7672 26658
rect 7628 26642 7636 26650
rect 7644 26639 7646 26650
rect 7656 26642 7664 26650
rect 7668 26639 7670 26650
rect 7716 26639 7718 26791
rect 7735 26785 7742 26833
rect 7744 26785 7753 26839
rect 7764 26833 7766 26937
rect 7779 26895 7781 26899
rect 7789 26881 7791 26895
rect 7754 26791 7760 26833
rect 7762 26785 7769 26833
rect 7771 26791 7780 26843
rect 7793 26791 7797 26849
rect 7810 26831 7814 26839
rect 7798 26791 7809 26831
rect 7811 26791 7814 26831
rect 7740 26658 7742 26785
rect 7745 26783 7752 26785
rect 7764 26658 7766 26785
rect 7793 26783 7796 26791
rect 7820 26667 7824 26791
rect 7730 26650 7742 26658
rect 7758 26650 7768 26658
rect 7790 26650 7798 26658
rect 7724 26642 7730 26650
rect 7740 26639 7742 26650
rect 7752 26642 7758 26650
rect 7764 26639 7766 26650
rect 7798 26642 7806 26650
rect 7836 26639 7838 26979
rect 7860 26977 7874 26979
rect 7860 26969 7862 26977
rect 7859 26961 7864 26969
rect 7860 26955 7864 26961
rect 7858 26929 7865 26955
rect 7840 26667 7846 26841
rect 7860 26831 7862 26929
rect 7873 26841 7876 26851
rect 7884 26841 7886 26979
rect 7922 26915 7925 26925
rect 7932 26917 7934 26979
rect 7945 26977 7950 26979
rect 7954 26953 7961 26979
rect 7932 26893 7936 26917
rect 7865 26831 7873 26841
rect 7883 26831 7886 26841
rect 7847 26793 7856 26831
rect 7858 26793 7863 26831
rect 7867 26793 7873 26831
rect 7874 26793 7890 26831
rect 7858 26785 7865 26793
rect 7884 26785 7890 26793
rect 7860 26658 7862 26785
rect 7884 26658 7886 26785
rect 7894 26667 7900 26841
rect 7904 26833 7910 26841
rect 7916 26793 7922 26833
rect 7916 26667 7920 26793
rect 7852 26650 7862 26658
rect 7880 26650 7890 26658
rect 7846 26642 7852 26650
rect 7860 26639 7862 26650
rect 7874 26642 7880 26650
rect 7884 26639 7886 26650
rect 7932 26639 7934 26893
rect 7936 26667 7942 26841
rect 7956 26833 7958 26953
rect 7969 26841 7972 26851
rect 7980 26841 7982 26979
rect 8052 26969 8057 26979
rect 8052 26953 8055 26969
rect 8056 26967 8057 26969
rect 8056 26953 8064 26967
rect 7961 26833 7969 26841
rect 7979 26833 7982 26841
rect 7943 26793 7952 26833
rect 7954 26793 7959 26833
rect 7963 26793 7969 26833
rect 7970 26793 7986 26833
rect 7954 26785 7961 26793
rect 7980 26785 7986 26793
rect 7956 26658 7958 26785
rect 7980 26658 7982 26785
rect 7990 26667 7996 26841
rect 8000 26833 8006 26841
rect 8012 26793 8018 26833
rect 8012 26667 8016 26793
rect 8052 26658 8054 26953
rect 8057 26919 8064 26953
rect 8148 26921 8150 26979
rect 8151 26969 8152 26979
rect 8151 26921 8158 26969
rect 8171 26961 8185 26969
rect 8148 26915 8158 26921
rect 8083 26667 8092 26843
rect 8148 26658 8150 26915
rect 8159 26911 8162 26915
rect 8170 26911 8175 26959
rect 8169 26841 8175 26851
rect 8185 26841 8188 26851
rect 8196 26841 8198 26979
rect 8234 26915 8237 26925
rect 8244 26917 8246 26979
rect 8257 26977 8262 26979
rect 8266 26953 8273 26979
rect 8244 26893 8248 26917
rect 8179 26793 8185 26841
rect 8195 26793 8198 26841
rect 8216 26833 8222 26841
rect 8196 26658 8198 26793
rect 8228 26793 8234 26833
rect 8228 26667 8232 26793
rect 7948 26650 7958 26658
rect 7976 26650 7984 26658
rect 8046 26650 8054 26658
rect 8074 26650 8080 26658
rect 8106 26650 8114 26658
rect 8134 26650 8150 26658
rect 8164 26650 8176 26658
rect 8192 26650 8204 26658
rect 7940 26642 7948 26650
rect 7956 26639 7958 26650
rect 7968 26642 7976 26650
rect 7980 26639 7982 26650
rect 8036 26642 8046 26650
rect 8052 26639 8054 26650
rect 8064 26642 8074 26650
rect 8114 26642 8122 26650
rect 8148 26639 8150 26650
rect 8162 26642 8164 26650
rect 8176 26642 8178 26650
rect 8190 26642 8192 26650
rect 8196 26639 8198 26650
rect 8204 26642 8206 26650
rect 8244 26639 8246 26893
rect 8248 26667 8254 26841
rect 8268 26833 8270 26953
rect 8281 26841 8284 26851
rect 8292 26841 8294 26979
rect 8330 26915 8333 26925
rect 8340 26917 8342 26979
rect 8353 26977 8358 26979
rect 8362 26953 8369 26979
rect 8340 26893 8344 26917
rect 8273 26833 8281 26841
rect 8291 26833 8294 26841
rect 8255 26793 8264 26833
rect 8266 26793 8271 26833
rect 8275 26793 8281 26833
rect 8282 26793 8298 26833
rect 8266 26785 8273 26793
rect 8292 26785 8298 26793
rect 8268 26658 8270 26785
rect 8292 26658 8294 26785
rect 8302 26667 8308 26841
rect 8312 26833 8318 26841
rect 8324 26793 8330 26833
rect 8324 26667 8328 26793
rect 8260 26650 8270 26658
rect 8288 26650 8296 26658
rect 8252 26642 8260 26650
rect 8268 26639 8270 26650
rect 8280 26642 8288 26650
rect 8292 26639 8294 26650
rect 8340 26639 8342 26893
rect 8344 26667 8350 26841
rect 8364 26833 8366 26953
rect 8377 26841 8380 26851
rect 8388 26841 8390 26979
rect 8436 26917 8439 26979
rect 8456 26972 8465 26979
rect 8460 26969 8464 26972
rect 8460 26953 8463 26969
rect 8423 26907 8428 26913
rect 8423 26903 8430 26907
rect 8436 26903 8440 26917
rect 8433 26893 8440 26903
rect 8433 26889 8438 26893
rect 8436 26843 8438 26889
rect 8453 26849 8457 26889
rect 8460 26849 8462 26953
rect 8369 26833 8377 26841
rect 8387 26833 8390 26841
rect 8351 26793 8360 26833
rect 8362 26793 8367 26833
rect 8371 26793 8377 26833
rect 8378 26793 8394 26833
rect 8362 26785 8369 26793
rect 8388 26785 8394 26793
rect 8364 26658 8366 26785
rect 8388 26658 8390 26785
rect 8398 26667 8404 26841
rect 8408 26833 8414 26841
rect 8420 26793 8426 26833
rect 8420 26667 8424 26793
rect 8436 26791 8446 26843
rect 8453 26839 8463 26849
rect 8465 26839 8472 26972
rect 8473 26953 8476 26963
rect 8484 26953 8486 26979
rect 8483 26937 8486 26953
rect 8460 26833 8462 26839
rect 8447 26791 8453 26833
rect 8356 26650 8366 26658
rect 8384 26650 8392 26658
rect 8348 26642 8356 26650
rect 8364 26639 8366 26650
rect 8376 26642 8384 26650
rect 8388 26639 8390 26650
rect 8436 26639 8438 26791
rect 8455 26785 8462 26833
rect 8464 26785 8473 26839
rect 8484 26833 8486 26937
rect 8543 26903 8548 26913
rect 8556 26903 8558 26979
rect 8579 26977 8592 26979
rect 8579 26972 8582 26977
rect 8499 26895 8501 26899
rect 8509 26881 8511 26895
rect 8553 26889 8558 26903
rect 8474 26791 8480 26833
rect 8482 26785 8489 26833
rect 8491 26791 8500 26843
rect 8513 26791 8517 26849
rect 8556 26841 8558 26889
rect 8580 26969 8582 26972
rect 8580 26945 8584 26969
rect 8530 26831 8534 26839
rect 8518 26791 8529 26831
rect 8531 26791 8534 26831
rect 8556 26791 8566 26841
rect 8574 26839 8577 26849
rect 8580 26831 8582 26945
rect 8585 26839 8592 26972
rect 8593 26953 8596 26963
rect 8604 26953 8606 26979
rect 8673 26964 8678 26979
rect 8603 26937 8606 26953
rect 8567 26791 8573 26831
rect 8460 26658 8462 26785
rect 8465 26783 8472 26785
rect 8484 26658 8486 26785
rect 8513 26783 8516 26791
rect 8540 26667 8544 26791
rect 8450 26650 8462 26658
rect 8478 26650 8488 26658
rect 8510 26650 8518 26658
rect 8538 26650 8554 26658
rect 8444 26642 8450 26650
rect 8460 26639 8462 26650
rect 8472 26642 8478 26650
rect 8484 26639 8486 26650
rect 8518 26642 8526 26650
rect 8556 26639 8558 26791
rect 8575 26783 8582 26831
rect 8584 26783 8593 26839
rect 8604 26831 8606 26937
rect 8663 26903 8668 26913
rect 8676 26903 8678 26964
rect 8692 26945 8695 26979
rect 8700 26969 8702 26979
rect 8700 26945 8704 26969
rect 8619 26895 8621 26899
rect 8629 26881 8631 26895
rect 8673 26889 8678 26903
rect 8594 26791 8600 26831
rect 8602 26783 8609 26831
rect 8611 26791 8620 26841
rect 8633 26791 8637 26849
rect 8676 26841 8678 26889
rect 8692 26851 8695 26929
rect 8689 26841 8695 26851
rect 8700 26891 8702 26945
rect 8705 26891 8709 26979
rect 8700 26841 8709 26891
rect 8719 26841 8722 26979
rect 8650 26831 8654 26839
rect 8676 26831 8685 26841
rect 8699 26831 8712 26841
rect 8724 26831 8726 26979
rect 8768 26978 8774 26979
rect 8761 26841 8764 26851
rect 8772 26841 8774 26978
rect 8820 26903 8822 26979
rect 8833 26977 8839 26979
rect 8842 26970 8849 26979
rect 8844 26903 8846 26970
rect 8820 26901 8851 26903
rect 8740 26833 8744 26841
rect 8768 26833 8774 26841
rect 8794 26833 8798 26841
rect 8638 26791 8649 26831
rect 8651 26791 8654 26831
rect 8674 26793 8685 26831
rect 8687 26793 8690 26831
rect 8692 26793 8703 26831
rect 8705 26793 8712 26831
rect 8714 26793 8717 26831
rect 8633 26783 8636 26791
rect 8580 26658 8582 26783
rect 8604 26658 8606 26783
rect 8660 26667 8664 26791
rect 8570 26650 8582 26658
rect 8598 26650 8610 26658
rect 8630 26650 8638 26658
rect 8658 26650 8672 26658
rect 8566 26642 8570 26650
rect 8580 26639 8582 26650
rect 8594 26642 8598 26650
rect 8604 26639 8606 26650
rect 8638 26642 8646 26650
rect 8672 26642 8674 26650
rect 8676 26639 8678 26793
rect 8692 26785 8699 26793
rect 8700 26658 8702 26793
rect 8719 26785 8726 26831
rect 8728 26793 8730 26831
rect 8724 26658 8726 26785
rect 8750 26667 8754 26833
rect 8755 26793 8766 26833
rect 8768 26793 8775 26833
rect 8777 26793 8780 26833
rect 8782 26793 8793 26833
rect 8795 26793 8798 26833
rect 8688 26650 8702 26658
rect 8716 26650 8728 26658
rect 8748 26650 8756 26658
rect 8686 26642 8688 26650
rect 8700 26639 8702 26650
rect 8714 26642 8716 26650
rect 8724 26639 8726 26650
rect 8728 26642 8730 26650
rect 8756 26642 8764 26650
rect 8772 26639 8774 26793
rect 8775 26785 8780 26793
rect 8804 26667 8808 26793
rect 8820 26658 8822 26901
rect 8824 26667 8830 26841
rect 8844 26833 8846 26901
rect 8857 26841 8860 26851
rect 8868 26841 8870 26979
rect 8914 26893 8933 26902
rect 9026 26882 9033 26979
rect 9076 26976 9079 26979
rect 9152 26968 9155 26979
rect 9193 26970 9196 26979
rect 9211 26978 9297 26979
rect 9246 26960 9249 26961
rect 9056 26952 9062 26960
rect 9069 26952 9083 26960
rect 9143 26952 9152 26953
rect 9212 26952 9214 26960
rect 9221 26952 9255 26960
rect 9076 26950 9079 26952
rect 9152 26950 9155 26952
rect 9062 26902 9069 26950
rect 9072 26902 9073 26942
rect 9057 26894 9066 26902
rect 9076 26894 9083 26942
rect 9094 26902 9101 26950
rect 9145 26947 9159 26950
rect 9152 26942 9159 26947
rect 9133 26902 9136 26942
rect 9088 26894 9133 26902
rect 9138 26894 9145 26942
rect 9153 26894 9159 26942
rect 9210 26902 9212 26942
rect 9214 26902 9221 26950
rect 9241 26947 9262 26950
rect 9255 26942 9262 26947
rect 9308 26942 9312 26978
rect 9229 26902 9230 26942
rect 9179 26894 9186 26902
rect 9232 26894 9239 26942
rect 9243 26902 9247 26942
rect 9255 26902 9259 26942
rect 9286 26902 9287 26942
rect 9262 26894 9269 26902
rect 9295 26894 9302 26942
rect 9076 26882 9079 26894
rect 9152 26892 9159 26894
rect 9152 26882 9155 26892
rect 9016 26874 9088 26882
rect 9133 26874 9210 26882
rect 9026 26872 9033 26874
rect 9036 26856 9040 26862
rect 8849 26833 8857 26841
rect 8867 26833 8870 26841
rect 8831 26793 8840 26833
rect 8842 26793 8847 26833
rect 8851 26793 8857 26833
rect 8858 26793 8874 26833
rect 8842 26785 8849 26793
rect 8868 26785 8874 26793
rect 8844 26658 8846 26785
rect 8868 26658 8870 26785
rect 8878 26667 8884 26841
rect 8888 26833 8894 26841
rect 8900 26793 8906 26833
rect 8900 26667 8904 26793
rect 8924 26667 8926 26843
rect 8952 26824 8957 26833
rect 8927 26785 8940 26824
rect 8950 26785 8952 26824
rect 8954 26785 8957 26824
rect 8960 26785 8970 26824
rect 9026 26816 9033 26856
rect 9076 26841 9079 26874
rect 9080 26864 9083 26874
rect 9090 26854 9093 26864
rect 9090 26848 9106 26854
rect 9134 26848 9146 26854
rect 9048 26824 9052 26834
rect 9062 26826 9084 26834
rect 9062 26825 9078 26826
rect 9152 26824 9155 26874
rect 9178 26854 9300 26859
rect 9204 26839 9222 26846
rect 9159 26826 9179 26834
rect 9308 26826 9312 26894
rect 9058 26820 9076 26824
rect 8945 26777 8950 26785
rect 9018 26768 9025 26816
rect 9058 26776 9064 26820
rect 9094 26776 9101 26824
rect 9152 26816 9160 26824
rect 9214 26816 9221 26824
rect 9134 26776 9136 26816
rect 9036 26768 9052 26775
rect 9058 26768 9062 26776
rect 9138 26768 9145 26816
rect 9153 26768 9160 26816
rect 9196 26777 9204 26816
rect 9196 26776 9212 26777
rect 9026 26705 9033 26768
rect 9152 26765 9160 26768
rect 9179 26765 9186 26776
rect 9204 26768 9212 26776
rect 9232 26768 9239 26816
rect 9241 26776 9245 26816
rect 9255 26776 9257 26824
rect 9262 26768 9269 26816
rect 9274 26778 9280 26816
rect 9308 26778 9315 26826
rect 9317 26778 9321 26816
rect 9295 26768 9302 26778
rect 9378 26771 9382 26818
rect 9451 26815 9454 26841
rect 9462 26815 9468 26979
rect 9492 26824 9499 26979
rect 9396 26783 9397 26813
rect 9443 26805 9445 26815
rect 9462 26805 9469 26815
rect 9482 26805 9489 26824
rect 9505 26823 9517 26824
rect 9504 26807 9517 26823
rect 9453 26789 9455 26805
rect 9472 26789 9489 26805
rect 9378 26770 9395 26771
rect 9264 26767 9267 26768
rect 9308 26767 9312 26768
rect 9040 26747 9076 26755
rect 9152 26753 9155 26765
rect 9462 26763 9468 26789
rect 9474 26776 9489 26789
rect 9509 26776 9516 26807
rect 9541 26791 9545 26839
rect 9568 26826 9575 26972
rect 9603 26895 9605 26899
rect 9613 26881 9615 26895
rect 9550 26791 9557 26816
rect 9559 26783 9566 26816
rect 9128 26747 9176 26753
rect 9234 26747 9245 26755
rect 9075 26737 9076 26747
rect 9100 26745 9101 26747
rect 9094 26737 9101 26745
rect 9152 26743 9155 26747
rect 9026 26697 9042 26705
rect 9016 26685 9024 26695
rect 9026 26689 9035 26697
rect 9050 26687 9052 26715
rect 9075 26689 9083 26737
rect 9100 26697 9101 26737
rect 9121 26689 9128 26737
rect 9138 26727 9154 26737
rect 9214 26735 9221 26745
rect 9264 26735 9270 26755
rect 9278 26737 9287 26745
rect 9290 26737 9297 26755
rect 9342 26747 9359 26755
rect 9369 26747 9382 26755
rect 9380 26746 9382 26747
rect 9214 26719 9230 26735
rect 9192 26693 9198 26699
rect 9290 26697 9299 26737
rect 9352 26697 9363 26737
rect 9381 26697 9382 26746
rect 9435 26737 9441 26755
rect 9447 26747 9455 26759
rect 9492 26755 9499 26776
rect 9568 26768 9576 26826
rect 9577 26791 9584 26816
rect 9586 26783 9593 26816
rect 9595 26791 9603 26826
rect 9617 26791 9621 26849
rect 9634 26831 9638 26839
rect 9622 26791 9633 26831
rect 9635 26791 9638 26831
rect 9617 26783 9620 26791
rect 9458 26751 9482 26755
rect 9489 26751 9500 26755
rect 9458 26747 9471 26751
rect 9447 26745 9457 26747
rect 9462 26745 9468 26747
rect 9492 26745 9499 26751
rect 9510 26745 9517 26747
rect 9451 26742 9462 26745
rect 9469 26742 9476 26745
rect 9451 26737 9460 26742
rect 9481 26737 9490 26745
rect 9509 26737 9517 26745
rect 9523 26737 9527 26751
rect 9428 26697 9431 26737
rect 9433 26697 9440 26737
rect 9444 26697 9448 26737
rect 9451 26697 9458 26737
rect 9463 26697 9470 26737
rect 9474 26697 9479 26737
rect 9482 26697 9489 26737
rect 9491 26697 9500 26737
rect 9501 26697 9507 26737
rect 9509 26697 9516 26737
rect 9188 26689 9192 26693
rect 9254 26685 9260 26695
rect 9290 26689 9297 26697
rect 9428 26689 9448 26697
rect 9462 26689 9469 26697
rect 9491 26689 9499 26697
rect 9520 26689 9527 26737
rect 9568 26689 9576 26747
rect 9026 26677 9034 26685
rect 9264 26677 9270 26685
rect 9494 26677 9497 26689
rect 9026 26669 9142 26677
rect 9264 26669 9271 26677
rect 9287 26669 9305 26677
rect 9321 26669 9336 26677
rect 9494 26669 9501 26677
rect 9517 26669 9563 26677
rect 9568 26669 9573 26689
rect 9644 26667 9648 26791
rect 8776 26650 8784 26658
rect 8804 26650 8822 26658
rect 8836 26650 8848 26658
rect 8864 26650 8876 26658
rect 8934 26650 8940 26658
rect 8962 26650 8968 26658
rect 8994 26650 9002 26658
rect 9022 26650 9030 26658
rect 9050 26650 9058 26658
rect 9078 26650 9086 26658
rect 9089 26656 9102 26658
rect 9106 26650 9114 26658
rect 9134 26650 9142 26658
rect 9147 26656 9158 26658
rect 9162 26650 9170 26658
rect 9190 26650 9198 26658
rect 9218 26650 9226 26658
rect 9246 26650 9254 26658
rect 9274 26650 9282 26658
rect 9302 26656 9320 26658
rect 9302 26650 9310 26656
rect 9358 26650 9364 26661
rect 9386 26650 9392 26661
rect 9428 26653 9436 26661
rect 9440 26653 9448 26661
rect 9456 26653 9464 26661
rect 9468 26653 9476 26661
rect 9484 26653 9492 26661
rect 9496 26653 9504 26661
rect 9512 26653 9520 26661
rect 9524 26653 9538 26658
rect 9554 26653 9566 26658
rect 9582 26653 9594 26658
rect 9440 26652 9456 26653
rect 9468 26652 9484 26653
rect 9496 26652 9512 26653
rect 9524 26652 9532 26653
rect 8784 26642 8792 26650
rect 8820 26639 8822 26650
rect 8832 26642 8836 26650
rect 8844 26639 8846 26650
rect 8860 26642 8864 26650
rect 8868 26639 8870 26650
rect 8924 26642 8934 26650
rect 8952 26642 8962 26650
rect 9002 26642 9010 26650
rect 9030 26642 9038 26650
rect 9058 26642 9066 26650
rect 9086 26642 9094 26650
rect 9114 26642 9122 26650
rect 9142 26642 9150 26650
rect 9170 26642 9178 26650
rect 9198 26642 9206 26650
rect 9226 26642 9234 26650
rect 9254 26642 9262 26650
rect 9282 26642 9290 26650
rect 9310 26642 9318 26650
rect 9364 26645 9374 26650
rect 9392 26645 9402 26650
rect 9448 26645 9456 26652
rect 9476 26645 9484 26652
rect 9504 26645 9512 26652
rect 9538 26642 9540 26653
rect 9552 26642 9554 26653
rect 9566 26642 9568 26653
rect 9580 26642 9582 26653
rect 9594 26642 9596 26653
rect 9614 26650 9622 26658
rect 9622 26642 9630 26650
rect 9000 26639 9036 26642
rect 9386 26639 9420 26641
rect 9660 26639 9662 26979
rect 9684 26977 9698 26979
rect 9684 26969 9686 26977
rect 9683 26961 9688 26969
rect 9684 26955 9688 26961
rect 9682 26929 9689 26955
rect 9664 26667 9670 26841
rect 9684 26831 9686 26929
rect 9697 26841 9700 26851
rect 9708 26841 9710 26979
rect 9746 26915 9749 26925
rect 9756 26917 9758 26979
rect 9769 26977 9774 26979
rect 9778 26953 9785 26979
rect 9756 26893 9760 26917
rect 9689 26831 9697 26841
rect 9707 26831 9710 26841
rect 9671 26793 9680 26831
rect 9682 26793 9687 26831
rect 9691 26793 9697 26831
rect 9698 26793 9714 26831
rect 9682 26785 9689 26793
rect 9708 26785 9714 26793
rect 9684 26658 9686 26785
rect 9708 26658 9710 26785
rect 9718 26667 9724 26841
rect 9728 26833 9734 26841
rect 9740 26793 9746 26833
rect 9740 26667 9744 26793
rect 9676 26650 9686 26658
rect 9704 26650 9714 26658
rect 9670 26642 9676 26650
rect 9684 26639 9686 26650
rect 9698 26642 9704 26650
rect 9708 26639 9710 26650
rect 9756 26639 9758 26893
rect 9760 26667 9766 26841
rect 9780 26833 9782 26953
rect 9793 26841 9796 26851
rect 9804 26841 9806 26979
rect 9842 26915 9845 26925
rect 9852 26917 9854 26979
rect 9865 26977 9870 26979
rect 9874 26953 9881 26979
rect 9852 26893 9856 26917
rect 9785 26833 9793 26841
rect 9803 26833 9806 26841
rect 9767 26793 9776 26833
rect 9778 26793 9783 26833
rect 9787 26793 9793 26833
rect 9794 26793 9810 26833
rect 9778 26785 9785 26793
rect 9804 26785 9810 26793
rect 9780 26658 9782 26785
rect 9804 26658 9806 26785
rect 9814 26667 9820 26841
rect 9824 26833 9830 26841
rect 9836 26793 9842 26833
rect 9836 26667 9840 26793
rect 9772 26650 9782 26658
rect 9800 26650 9808 26658
rect 9764 26642 9772 26650
rect 9780 26639 9782 26650
rect 9792 26642 9800 26650
rect 9804 26639 9806 26650
rect 9852 26639 9854 26893
rect 9856 26667 9862 26841
rect 9876 26833 9878 26953
rect 9889 26841 9892 26851
rect 9900 26841 9902 26979
rect 9948 26917 9951 26979
rect 9968 26972 9977 26979
rect 9972 26969 9976 26972
rect 9972 26953 9975 26969
rect 9935 26907 9940 26913
rect 9935 26903 9942 26907
rect 9948 26903 9952 26917
rect 9945 26893 9952 26903
rect 9945 26889 9950 26893
rect 9948 26843 9950 26889
rect 9965 26849 9969 26889
rect 9972 26849 9974 26953
rect 9881 26833 9889 26841
rect 9899 26833 9902 26841
rect 9863 26793 9872 26833
rect 9874 26793 9879 26833
rect 9883 26793 9889 26833
rect 9890 26793 9906 26833
rect 9874 26785 9881 26793
rect 9900 26785 9906 26793
rect 9876 26658 9878 26785
rect 9900 26658 9902 26785
rect 9910 26667 9916 26841
rect 9920 26833 9926 26841
rect 9932 26793 9938 26833
rect 9932 26667 9936 26793
rect 9948 26791 9958 26843
rect 9965 26839 9975 26849
rect 9977 26839 9984 26972
rect 9985 26953 9988 26963
rect 9996 26953 9998 26979
rect 9995 26937 9998 26953
rect 9972 26833 9974 26839
rect 9959 26791 9965 26833
rect 9868 26650 9878 26658
rect 9896 26650 9904 26658
rect 9860 26642 9868 26650
rect 9876 26639 9878 26650
rect 9888 26642 9896 26650
rect 9900 26639 9902 26650
rect 9948 26639 9950 26791
rect 9967 26785 9974 26833
rect 9976 26785 9985 26839
rect 9996 26833 9998 26937
rect 10011 26895 10013 26899
rect 10021 26881 10023 26895
rect 9986 26791 9992 26833
rect 9994 26785 10001 26833
rect 10003 26791 10012 26843
rect 10025 26791 10029 26849
rect 10042 26831 10046 26839
rect 10030 26791 10041 26831
rect 10043 26791 10046 26831
rect 9972 26658 9974 26785
rect 9977 26783 9984 26785
rect 9996 26658 9998 26785
rect 10025 26783 10028 26791
rect 10052 26667 10056 26791
rect 9962 26650 9974 26658
rect 9990 26650 10000 26658
rect 10022 26650 10030 26658
rect 9956 26642 9962 26650
rect 9972 26639 9974 26650
rect 9984 26642 9990 26650
rect 9996 26639 9998 26650
rect 10030 26642 10038 26650
rect 10068 26639 10070 26979
rect 10092 26977 10106 26979
rect 10092 26969 10094 26977
rect 10091 26961 10096 26969
rect 10092 26955 10096 26961
rect 10090 26929 10097 26955
rect 10072 26667 10078 26841
rect 10092 26831 10094 26929
rect 10105 26841 10108 26851
rect 10116 26841 10118 26979
rect 10154 26915 10157 26925
rect 10164 26917 10166 26979
rect 10177 26977 10182 26979
rect 10186 26953 10193 26979
rect 10164 26893 10168 26917
rect 10097 26831 10105 26841
rect 10115 26831 10118 26841
rect 10079 26793 10088 26831
rect 10090 26793 10095 26831
rect 10099 26793 10105 26831
rect 10106 26793 10122 26831
rect 10090 26785 10097 26793
rect 10116 26785 10122 26793
rect 10092 26658 10094 26785
rect 10116 26658 10118 26785
rect 10126 26667 10132 26841
rect 10136 26833 10142 26841
rect 10148 26793 10154 26833
rect 10148 26667 10152 26793
rect 10084 26650 10094 26658
rect 10112 26650 10122 26658
rect 10078 26642 10084 26650
rect 10092 26639 10094 26650
rect 10106 26642 10112 26650
rect 10116 26639 10118 26650
rect 10164 26639 10166 26893
rect 10168 26667 10174 26841
rect 10188 26833 10190 26953
rect 10201 26841 10204 26851
rect 10212 26841 10214 26979
rect 10260 26917 10263 26979
rect 10280 26972 10289 26979
rect 10284 26969 10288 26972
rect 10284 26953 10287 26969
rect 10247 26907 10252 26913
rect 10247 26903 10254 26907
rect 10260 26903 10264 26917
rect 10257 26893 10264 26903
rect 10257 26889 10262 26893
rect 10260 26843 10262 26889
rect 10277 26849 10281 26889
rect 10284 26849 10286 26953
rect 10193 26833 10201 26841
rect 10211 26833 10214 26841
rect 10175 26793 10184 26833
rect 10186 26793 10191 26833
rect 10195 26793 10201 26833
rect 10202 26793 10218 26833
rect 10186 26785 10193 26793
rect 10212 26785 10218 26793
rect 10188 26658 10190 26785
rect 10212 26658 10214 26785
rect 10222 26667 10228 26841
rect 10232 26833 10238 26841
rect 10244 26793 10250 26833
rect 10244 26667 10248 26793
rect 10260 26791 10270 26843
rect 10277 26839 10287 26849
rect 10289 26839 10296 26972
rect 10297 26953 10300 26963
rect 10308 26953 10310 26979
rect 10307 26937 10310 26953
rect 10284 26833 10286 26839
rect 10271 26791 10277 26833
rect 10180 26650 10190 26658
rect 10208 26650 10216 26658
rect 10172 26642 10180 26650
rect 10188 26639 10190 26650
rect 10200 26642 10208 26650
rect 10212 26639 10214 26650
rect 10260 26639 10262 26791
rect 10279 26785 10286 26833
rect 10288 26785 10297 26839
rect 10308 26833 10310 26937
rect 10323 26895 10325 26899
rect 10333 26881 10335 26895
rect 10298 26791 10304 26833
rect 10306 26785 10313 26833
rect 10315 26791 10324 26843
rect 10337 26791 10341 26849
rect 10354 26831 10358 26839
rect 10342 26791 10353 26831
rect 10355 26791 10358 26831
rect 10284 26658 10286 26785
rect 10289 26783 10296 26785
rect 10308 26658 10310 26785
rect 10337 26783 10340 26791
rect 10364 26667 10368 26791
rect 10274 26650 10286 26658
rect 10302 26650 10312 26658
rect 10334 26650 10342 26658
rect 10268 26642 10274 26650
rect 10284 26639 10286 26650
rect 10296 26642 10302 26650
rect 10308 26639 10310 26650
rect 10342 26642 10350 26650
rect 10380 26639 10382 26979
rect 10404 26977 10418 26979
rect 10404 26969 10406 26977
rect 10403 26961 10408 26969
rect 10404 26955 10408 26961
rect 10402 26929 10409 26955
rect 10384 26667 10390 26841
rect 10404 26831 10406 26929
rect 10417 26841 10420 26851
rect 10428 26841 10430 26979
rect 10466 26915 10469 26925
rect 10476 26917 10478 26979
rect 10489 26977 10494 26979
rect 10498 26953 10505 26979
rect 10476 26893 10480 26917
rect 10409 26831 10417 26841
rect 10427 26831 10430 26841
rect 10391 26793 10400 26831
rect 10402 26793 10407 26831
rect 10411 26793 10417 26831
rect 10418 26793 10434 26831
rect 10402 26785 10409 26793
rect 10428 26785 10434 26793
rect 10404 26658 10406 26785
rect 10428 26658 10430 26785
rect 10438 26667 10444 26841
rect 10448 26833 10454 26841
rect 10460 26793 10466 26833
rect 10460 26667 10464 26793
rect 10396 26650 10406 26658
rect 10424 26650 10434 26658
rect 10390 26642 10396 26650
rect 10404 26639 10406 26650
rect 10418 26642 10424 26650
rect 10428 26639 10430 26650
rect 10476 26639 10478 26893
rect 10480 26667 10486 26841
rect 10500 26833 10502 26953
rect 10513 26841 10516 26851
rect 10524 26841 10526 26979
rect 10562 26915 10565 26925
rect 10572 26917 10574 26979
rect 10585 26977 10590 26979
rect 10594 26953 10601 26979
rect 10572 26893 10576 26917
rect 10505 26833 10513 26841
rect 10523 26833 10526 26841
rect 10487 26793 10496 26833
rect 10498 26793 10503 26833
rect 10507 26793 10513 26833
rect 10514 26793 10530 26833
rect 10498 26785 10505 26793
rect 10524 26785 10530 26793
rect 10500 26658 10502 26785
rect 10524 26658 10526 26785
rect 10534 26667 10540 26841
rect 10544 26833 10550 26841
rect 10556 26793 10562 26833
rect 10556 26667 10560 26793
rect 10492 26650 10502 26658
rect 10520 26650 10528 26658
rect 10484 26642 10492 26650
rect 10500 26639 10502 26650
rect 10512 26642 10520 26650
rect 10524 26639 10526 26650
rect 10572 26639 10574 26893
rect 10576 26667 10582 26841
rect 10596 26833 10598 26953
rect 10609 26841 10612 26851
rect 10620 26841 10622 26979
rect 10668 26917 10671 26979
rect 10688 26972 10697 26979
rect 10692 26969 10696 26972
rect 10692 26953 10695 26969
rect 10655 26907 10660 26913
rect 10655 26903 10662 26907
rect 10668 26903 10672 26917
rect 10665 26893 10672 26903
rect 10665 26889 10670 26893
rect 10668 26843 10670 26889
rect 10685 26849 10689 26889
rect 10692 26849 10694 26953
rect 10601 26833 10609 26841
rect 10619 26833 10622 26841
rect 10583 26793 10592 26833
rect 10594 26793 10599 26833
rect 10603 26793 10609 26833
rect 10610 26793 10626 26833
rect 10594 26785 10601 26793
rect 10620 26785 10626 26793
rect 10596 26658 10598 26785
rect 10620 26658 10622 26785
rect 10630 26667 10636 26841
rect 10640 26833 10646 26841
rect 10652 26793 10658 26833
rect 10652 26667 10656 26793
rect 10668 26791 10678 26843
rect 10685 26839 10695 26849
rect 10697 26839 10704 26972
rect 10705 26953 10708 26963
rect 10716 26953 10718 26979
rect 10715 26937 10718 26953
rect 10692 26833 10694 26839
rect 10679 26791 10685 26833
rect 10588 26650 10598 26658
rect 10616 26650 10624 26658
rect 10580 26642 10588 26650
rect 10596 26639 10598 26650
rect 10608 26642 10616 26650
rect 10620 26639 10622 26650
rect 10668 26639 10670 26791
rect 10687 26785 10694 26833
rect 10696 26785 10705 26839
rect 10716 26833 10718 26937
rect 10731 26895 10733 26899
rect 10741 26881 10743 26895
rect 10706 26791 10712 26833
rect 10714 26785 10721 26833
rect 10723 26791 10732 26843
rect 10745 26791 10749 26849
rect 10762 26831 10766 26839
rect 10750 26791 10761 26831
rect 10763 26791 10766 26831
rect 10692 26658 10694 26785
rect 10697 26783 10704 26785
rect 10716 26658 10718 26785
rect 10745 26783 10748 26791
rect 10772 26667 10776 26791
rect 10682 26650 10694 26658
rect 10710 26650 10720 26658
rect 10742 26650 10750 26658
rect 10770 26650 10786 26658
rect 10676 26642 10682 26650
rect 10692 26639 10694 26650
rect 10704 26642 10710 26650
rect 10716 26639 10718 26650
rect 10750 26642 10758 26650
rect 10788 26639 10790 26979
rect 10814 26977 10816 26979
rect 10791 26959 10797 26964
rect 10791 26945 10806 26959
rect 10791 26929 10807 26945
rect 10791 26916 10797 26929
rect 10817 26916 10819 26964
rect 10836 26658 10838 26979
rect 10956 26966 10958 26979
rect 10867 26916 10879 26956
rect 10929 26932 10934 26956
rect 10945 26955 10948 26965
rect 10954 26955 10955 26956
rect 10956 26955 10965 26966
rect 10954 26939 10958 26955
rect 10996 26948 11005 26979
rect 11044 26947 11047 26979
rect 11052 26971 11054 26979
rect 11052 26947 11056 26971
rect 10928 26916 10944 26932
rect 10929 26908 10934 26916
rect 10954 26908 10955 26939
rect 10931 26789 10935 26847
rect 10956 26658 10958 26939
rect 10982 26934 10984 26939
rect 10994 26934 10996 26939
rect 10996 26929 11004 26934
rect 11006 26924 11014 26929
rect 11025 26921 11030 26934
rect 10963 26789 10965 26919
rect 11035 26911 11039 26913
rect 11044 26911 11047 26931
rect 11003 26883 11009 26909
rect 11025 26908 11030 26911
rect 11039 26903 11047 26911
rect 11044 26851 11047 26903
rect 10984 26819 10989 26847
rect 11041 26841 11047 26851
rect 11052 26891 11054 26947
rect 11057 26891 11061 26979
rect 11071 26891 11074 26979
rect 11052 26841 11061 26891
rect 11076 26885 11078 26979
rect 11120 26978 11126 26979
rect 11071 26841 11074 26875
rect 11076 26861 11085 26885
rect 11002 26829 11006 26837
rect 10985 26789 10989 26819
rect 10990 26789 11001 26829
rect 11003 26789 11006 26829
rect 11026 26793 11028 26829
rect 11030 26793 11037 26841
rect 11051 26829 11064 26841
rect 11076 26829 11078 26861
rect 11113 26841 11116 26851
rect 11124 26841 11126 26978
rect 11160 26956 11164 26966
rect 11172 26956 11174 26979
rect 11170 26942 11174 26956
rect 11092 26833 11096 26841
rect 11120 26833 11126 26841
rect 11146 26833 11150 26841
rect 11172 26837 11174 26942
rect 11201 26932 11208 26979
rect 11209 26955 11212 26965
rect 11220 26955 11222 26979
rect 11219 26939 11222 26955
rect 11260 26948 11269 26979
rect 11296 26947 11304 26956
rect 11295 26942 11304 26947
rect 11183 26847 11192 26883
rect 11183 26837 11193 26847
rect 11201 26837 11208 26916
rect 11162 26833 11181 26837
rect 11039 26793 11042 26829
rect 11044 26793 11055 26829
rect 11057 26793 11064 26829
rect 11066 26793 11069 26829
rect 10985 26781 10988 26789
rect 11012 26667 11016 26789
rect 11044 26785 11051 26793
rect 11052 26658 11054 26793
rect 11071 26785 11078 26829
rect 11080 26793 11082 26829
rect 11076 26658 11078 26785
rect 11102 26667 11106 26833
rect 11107 26793 11118 26833
rect 11120 26793 11127 26833
rect 11129 26793 11132 26833
rect 11134 26793 11145 26833
rect 11147 26793 11150 26833
rect 11172 26827 11181 26833
rect 10802 26650 10814 26658
rect 10830 26650 10842 26658
rect 10862 26650 10870 26658
rect 10926 26650 10934 26658
rect 10954 26650 10962 26658
rect 10986 26650 10994 26658
rect 11014 26650 11024 26658
rect 11042 26650 11054 26658
rect 11070 26650 11080 26658
rect 11100 26650 11108 26658
rect 10798 26642 10802 26650
rect 10826 26642 10830 26650
rect 10836 26639 10838 26650
rect 10870 26642 10878 26650
rect 10918 26642 10926 26650
rect 10946 26642 10954 26650
rect 10956 26639 10958 26650
rect 10994 26642 11002 26650
rect 11024 26642 11030 26650
rect 11052 26642 11058 26650
rect 11052 26639 11054 26642
rect 11076 26639 11078 26650
rect 11080 26642 11086 26650
rect 11108 26642 11116 26650
rect 11124 26639 11126 26793
rect 11127 26785 11132 26793
rect 11156 26667 11160 26793
rect 11172 26789 11182 26827
rect 11183 26789 11189 26833
rect 11128 26650 11136 26658
rect 11136 26642 11144 26650
rect 11172 26639 11174 26789
rect 11191 26785 11198 26833
rect 11200 26785 11209 26837
rect 11220 26833 11222 26939
rect 11246 26934 11248 26939
rect 11258 26934 11260 26939
rect 11260 26929 11268 26934
rect 11270 26924 11278 26929
rect 11292 26921 11294 26934
rect 11302 26932 11311 26942
rect 11321 26932 11328 26979
rect 11329 26955 11332 26965
rect 11340 26955 11342 26979
rect 11312 26931 11321 26932
rect 11336 26929 11338 26942
rect 11339 26939 11342 26955
rect 11380 26948 11389 26979
rect 11436 26971 11438 26979
rect 11456 26977 11460 26979
rect 11436 26957 11440 26971
rect 11456 26967 11466 26977
rect 11441 26957 11448 26967
rect 11436 26947 11448 26957
rect 11267 26883 11273 26909
rect 11292 26908 11294 26911
rect 11303 26847 11312 26911
rect 11210 26789 11216 26833
rect 11218 26785 11225 26833
rect 11227 26789 11236 26843
rect 11248 26819 11253 26847
rect 11303 26837 11313 26847
rect 11321 26837 11328 26916
rect 11340 26885 11342 26939
rect 11366 26934 11368 26939
rect 11378 26934 11380 26939
rect 11380 26929 11388 26934
rect 11390 26924 11398 26929
rect 11347 26911 11356 26919
rect 11347 26885 11349 26901
rect 11340 26861 11349 26885
rect 11387 26883 11393 26909
rect 11266 26829 11270 26837
rect 11282 26829 11292 26837
rect 11249 26789 11253 26819
rect 11254 26789 11265 26829
rect 11267 26789 11270 26829
rect 11294 26827 11301 26837
rect 11293 26789 11302 26827
rect 11303 26789 11309 26829
rect 11201 26781 11208 26785
rect 11220 26658 11222 26785
rect 11249 26781 11252 26789
rect 11276 26667 11280 26789
rect 11311 26781 11318 26829
rect 11320 26781 11329 26837
rect 11340 26829 11342 26861
rect 11330 26789 11336 26829
rect 11338 26781 11345 26829
rect 11347 26789 11356 26839
rect 11368 26819 11373 26847
rect 11386 26829 11390 26837
rect 11369 26789 11373 26819
rect 11374 26789 11385 26829
rect 11387 26789 11390 26829
rect 11369 26781 11372 26789
rect 11340 26658 11342 26781
rect 11396 26667 11400 26789
rect 11436 26658 11438 26947
rect 11440 26931 11448 26947
rect 11441 26919 11448 26931
rect 11467 26911 11476 26967
rect 11532 26921 11534 26979
rect 11535 26969 11536 26979
rect 11535 26921 11542 26969
rect 11555 26961 11569 26969
rect 11532 26915 11542 26921
rect 11467 26861 11469 26901
rect 11467 26667 11476 26839
rect 11532 26658 11534 26915
rect 11543 26911 11546 26915
rect 11554 26911 11559 26959
rect 11553 26841 11559 26851
rect 11569 26841 11572 26851
rect 11580 26841 11582 26979
rect 11628 26917 11631 26979
rect 11648 26972 11657 26979
rect 11652 26969 11656 26972
rect 11652 26953 11655 26969
rect 11615 26907 11620 26913
rect 11615 26903 11622 26907
rect 11628 26903 11632 26917
rect 11625 26893 11632 26903
rect 11625 26889 11630 26893
rect 11628 26843 11630 26889
rect 11645 26849 11649 26889
rect 11652 26849 11654 26953
rect 11563 26793 11569 26841
rect 11579 26793 11582 26841
rect 11600 26833 11606 26841
rect 11580 26658 11582 26793
rect 11612 26793 11618 26833
rect 11612 26667 11616 26793
rect 11628 26791 11638 26843
rect 11645 26839 11655 26849
rect 11657 26839 11664 26972
rect 11665 26953 11668 26963
rect 11676 26953 11678 26979
rect 11675 26937 11678 26953
rect 11652 26833 11654 26839
rect 11639 26791 11645 26833
rect 11190 26650 11200 26658
rect 11218 26650 11228 26658
rect 11250 26650 11258 26658
rect 11278 26650 11294 26658
rect 11310 26650 11322 26658
rect 11338 26650 11350 26658
rect 11370 26650 11378 26658
rect 11398 26650 11414 26658
rect 11430 26650 11442 26658
rect 11458 26650 11470 26658
rect 11490 26650 11498 26658
rect 11518 26650 11534 26658
rect 11548 26650 11560 26658
rect 11576 26650 11588 26658
rect 11184 26642 11190 26650
rect 11212 26642 11218 26650
rect 11220 26639 11222 26650
rect 11258 26642 11266 26650
rect 11306 26642 11310 26650
rect 11334 26642 11338 26650
rect 11340 26639 11342 26650
rect 11378 26642 11386 26650
rect 11426 26642 11430 26650
rect 11436 26639 11438 26650
rect 11454 26642 11458 26650
rect 11498 26642 11506 26650
rect 11532 26639 11534 26650
rect 11546 26642 11548 26650
rect 11560 26642 11562 26650
rect 11574 26642 11576 26650
rect 11580 26639 11582 26650
rect 11588 26642 11590 26650
rect 11628 26639 11630 26791
rect 11647 26785 11654 26833
rect 11656 26785 11665 26839
rect 11676 26833 11678 26937
rect 11691 26895 11693 26899
rect 11701 26881 11703 26895
rect 11666 26791 11672 26833
rect 11674 26785 11681 26833
rect 11683 26791 11692 26843
rect 11705 26791 11709 26849
rect 11722 26831 11726 26839
rect 11710 26791 11721 26831
rect 11723 26791 11726 26831
rect 11652 26658 11654 26785
rect 11657 26783 11664 26785
rect 11676 26658 11678 26785
rect 11705 26783 11708 26791
rect 11732 26667 11736 26791
rect 11642 26650 11654 26658
rect 11670 26650 11680 26658
rect 11702 26650 11710 26658
rect 11636 26642 11642 26650
rect 11652 26639 11654 26650
rect 11664 26642 11670 26650
rect 11676 26639 11678 26650
rect 11710 26642 11718 26650
rect 11748 26639 11750 26979
rect 11772 26977 11786 26979
rect 11772 26969 11774 26977
rect 11771 26961 11776 26969
rect 11772 26955 11776 26961
rect 11770 26929 11777 26955
rect 11752 26667 11758 26841
rect 11772 26831 11774 26929
rect 11785 26841 11788 26851
rect 11796 26841 11798 26979
rect 11832 26956 11837 26966
rect 11844 26956 11847 26979
rect 11842 26953 11856 26956
rect 11842 26942 11847 26953
rect 11844 26917 11847 26942
rect 11873 26932 11880 26979
rect 11881 26955 11884 26965
rect 11892 26955 11894 26979
rect 11891 26939 11894 26955
rect 11932 26948 11941 26979
rect 11987 26972 11990 26979
rect 12008 26972 12010 26979
rect 11988 26971 11990 26972
rect 11988 26947 11992 26971
rect 11844 26893 11848 26917
rect 11777 26831 11785 26841
rect 11795 26831 11798 26841
rect 11759 26793 11768 26831
rect 11770 26793 11775 26831
rect 11779 26793 11785 26831
rect 11786 26793 11802 26831
rect 11770 26785 11777 26793
rect 11796 26785 11802 26793
rect 11772 26658 11774 26785
rect 11796 26658 11798 26785
rect 11806 26667 11812 26841
rect 11816 26833 11822 26841
rect 11844 26837 11846 26893
rect 11861 26847 11864 26893
rect 11861 26837 11871 26847
rect 11873 26837 11880 26916
rect 11834 26833 11853 26837
rect 11828 26793 11834 26833
rect 11844 26827 11853 26833
rect 11828 26667 11832 26793
rect 11844 26789 11854 26827
rect 11855 26789 11861 26833
rect 11764 26650 11774 26658
rect 11792 26650 11802 26658
rect 11758 26642 11764 26650
rect 11772 26639 11774 26650
rect 11786 26642 11792 26650
rect 11796 26639 11798 26650
rect 11844 26639 11846 26789
rect 11863 26785 11870 26833
rect 11872 26785 11881 26837
rect 11892 26833 11894 26939
rect 11918 26934 11920 26939
rect 11930 26934 11932 26939
rect 11932 26929 11940 26934
rect 11942 26924 11950 26929
rect 11964 26921 11966 26934
rect 11951 26911 11964 26913
rect 11974 26911 11975 26913
rect 11939 26883 11945 26909
rect 11951 26908 11956 26911
rect 11964 26908 11966 26911
rect 11975 26903 11984 26911
rect 11882 26789 11888 26833
rect 11890 26785 11897 26833
rect 11899 26789 11908 26843
rect 11920 26819 11925 26847
rect 11982 26839 11985 26849
rect 11938 26829 11942 26837
rect 11921 26789 11925 26819
rect 11926 26789 11937 26829
rect 11939 26789 11942 26829
rect 11965 26791 11974 26839
rect 11988 26829 11990 26947
rect 11993 26839 12000 26972
rect 12001 26953 12004 26963
rect 12012 26953 12014 26979
rect 12072 26956 12076 26966
rect 12084 26956 12086 26979
rect 12011 26937 12014 26953
rect 12082 26942 12086 26956
rect 12088 26945 12096 26956
rect 12087 26942 12096 26945
rect 12012 26885 12014 26937
rect 12027 26895 12029 26899
rect 12019 26885 12021 26889
rect 12012 26861 12021 26885
rect 12037 26881 12039 26895
rect 11975 26791 11981 26829
rect 11873 26781 11880 26785
rect 11892 26658 11894 26785
rect 11921 26781 11924 26789
rect 11948 26667 11952 26789
rect 11983 26783 11990 26829
rect 11988 26658 11990 26783
rect 11992 26781 12001 26839
rect 12012 26829 12014 26861
rect 12002 26791 12008 26829
rect 12010 26783 12017 26829
rect 12019 26791 12028 26839
rect 12041 26791 12045 26849
rect 12058 26831 12062 26839
rect 12084 26837 12086 26942
rect 12094 26932 12103 26942
rect 12113 26932 12120 26979
rect 12122 26977 12124 26979
rect 12121 26955 12124 26965
rect 12132 26955 12134 26979
rect 12131 26939 12134 26955
rect 12172 26948 12181 26979
rect 12228 26971 12230 26979
rect 12227 26961 12232 26971
rect 12248 26961 12254 26979
rect 12228 26957 12232 26961
rect 12104 26929 12113 26932
rect 12095 26847 12104 26881
rect 12095 26837 12105 26847
rect 12113 26837 12120 26916
rect 12074 26831 12093 26837
rect 12046 26791 12057 26831
rect 12059 26791 12062 26831
rect 12084 26827 12093 26831
rect 12041 26783 12044 26791
rect 12012 26658 12014 26783
rect 12068 26667 12072 26791
rect 12084 26789 12094 26827
rect 12095 26789 12101 26831
rect 11862 26650 11868 26658
rect 11890 26650 11896 26658
rect 11922 26650 11930 26658
rect 11950 26650 11962 26658
rect 11978 26650 11990 26658
rect 12006 26650 12018 26658
rect 12038 26650 12046 26658
rect 11852 26642 11862 26650
rect 11880 26642 11890 26650
rect 11892 26639 11894 26650
rect 11930 26642 11938 26650
rect 11962 26642 11966 26650
rect 11988 26642 11994 26650
rect 11988 26639 11990 26642
rect 12012 26639 12014 26650
rect 12018 26642 12022 26650
rect 12046 26642 12054 26650
rect 12084 26639 12086 26789
rect 12103 26783 12110 26831
rect 12112 26783 12121 26837
rect 12132 26831 12134 26939
rect 12158 26934 12160 26939
rect 12170 26934 12172 26939
rect 12172 26929 12180 26934
rect 12226 26931 12233 26957
rect 12182 26924 12190 26929
rect 12179 26883 12185 26909
rect 12204 26908 12206 26911
rect 12122 26789 12128 26831
rect 12130 26783 12137 26831
rect 12139 26789 12148 26841
rect 12160 26819 12165 26847
rect 12208 26839 12213 26841
rect 12178 26829 12182 26837
rect 12161 26789 12165 26819
rect 12166 26789 12177 26829
rect 12179 26789 12182 26829
rect 12113 26781 12120 26783
rect 12132 26658 12134 26783
rect 12161 26781 12164 26789
rect 12188 26667 12192 26789
rect 12208 26667 12214 26839
rect 12228 26829 12230 26931
rect 12252 26901 12254 26961
rect 12290 26915 12293 26925
rect 12300 26917 12302 26979
rect 12313 26977 12318 26979
rect 12322 26953 12329 26979
rect 12252 26885 12260 26901
rect 12300 26893 12304 26917
rect 12252 26861 12261 26885
rect 12241 26841 12244 26851
rect 12252 26841 12254 26861
rect 12233 26839 12240 26841
rect 12233 26829 12241 26839
rect 12251 26829 12254 26841
rect 12215 26793 12224 26829
rect 12226 26793 12231 26829
rect 12235 26793 12241 26829
rect 12242 26793 12258 26829
rect 12226 26785 12233 26793
rect 12252 26785 12258 26793
rect 12228 26658 12230 26785
rect 12252 26658 12254 26785
rect 12262 26667 12268 26839
rect 12272 26833 12278 26841
rect 12284 26793 12290 26833
rect 12284 26667 12288 26793
rect 12102 26650 12110 26658
rect 12130 26650 12138 26658
rect 12162 26650 12170 26658
rect 12190 26650 12204 26658
rect 12220 26650 12232 26658
rect 12248 26650 12260 26658
rect 12094 26642 12102 26650
rect 12122 26642 12130 26650
rect 12132 26639 12134 26650
rect 12170 26642 12178 26650
rect 12204 26642 12206 26650
rect 12218 26642 12220 26650
rect 12228 26639 12230 26650
rect 12232 26642 12234 26650
rect 12246 26642 12248 26650
rect 12252 26639 12254 26650
rect 12260 26642 12262 26650
rect 12300 26639 12302 26893
rect 12304 26667 12310 26841
rect 12324 26833 12326 26953
rect 12337 26841 12340 26851
rect 12348 26841 12350 26979
rect 12386 26915 12389 26925
rect 12396 26917 12398 26979
rect 12409 26977 12414 26979
rect 12418 26953 12425 26979
rect 12396 26893 12400 26917
rect 12329 26833 12337 26841
rect 12347 26833 12350 26841
rect 12311 26793 12320 26833
rect 12322 26793 12327 26833
rect 12331 26793 12337 26833
rect 12338 26793 12354 26833
rect 12322 26785 12329 26793
rect 12348 26785 12354 26793
rect 12324 26658 12326 26785
rect 12348 26658 12350 26785
rect 12358 26667 12364 26841
rect 12368 26833 12374 26841
rect 12380 26793 12386 26833
rect 12380 26667 12384 26793
rect 12316 26650 12326 26658
rect 12344 26650 12352 26658
rect 12308 26642 12316 26650
rect 12324 26639 12326 26650
rect 12336 26642 12344 26650
rect 12348 26639 12350 26650
rect 12396 26639 12398 26893
rect 12400 26667 12406 26841
rect 12420 26833 12422 26953
rect 12433 26841 12436 26851
rect 12444 26841 12446 26979
rect 12482 26915 12485 26925
rect 12492 26917 12494 26979
rect 12505 26977 12510 26979
rect 12514 26953 12521 26979
rect 12492 26893 12496 26917
rect 12425 26833 12433 26841
rect 12443 26833 12446 26841
rect 12407 26793 12416 26833
rect 12418 26793 12423 26833
rect 12427 26793 12433 26833
rect 12434 26793 12450 26833
rect 12418 26785 12425 26793
rect 12444 26785 12450 26793
rect 12420 26658 12422 26785
rect 12444 26658 12446 26785
rect 12454 26667 12460 26841
rect 12464 26833 12470 26841
rect 12476 26793 12482 26833
rect 12476 26667 12480 26793
rect 12412 26650 12422 26658
rect 12440 26650 12448 26658
rect 12404 26642 12412 26650
rect 12420 26639 12422 26650
rect 12432 26642 12440 26650
rect 12444 26639 12446 26650
rect 12492 26639 12494 26893
rect 12496 26667 12502 26841
rect 12516 26833 12518 26953
rect 12529 26841 12532 26851
rect 12540 26841 12542 26979
rect 12588 26917 12590 26979
rect 12591 26953 12607 26964
rect 12591 26917 12597 26953
rect 12588 26916 12597 26917
rect 12617 26916 12619 26964
rect 12588 26893 12592 26916
rect 12521 26833 12529 26841
rect 12539 26833 12542 26841
rect 12503 26793 12512 26833
rect 12514 26793 12519 26833
rect 12523 26793 12529 26833
rect 12530 26793 12546 26833
rect 12514 26785 12521 26793
rect 12540 26785 12546 26793
rect 12516 26658 12518 26785
rect 12540 26658 12542 26785
rect 12550 26667 12556 26841
rect 12560 26833 12566 26841
rect 12572 26793 12578 26833
rect 12572 26667 12576 26793
rect 12508 26650 12518 26658
rect 12536 26650 12544 26658
rect 12500 26642 12508 26650
rect 12516 26639 12518 26650
rect 12528 26642 12536 26650
rect 12540 26639 12542 26650
rect 12588 26639 12590 26893
rect 12636 26658 12638 26979
rect 12730 26977 12737 26979
rect 12730 26966 12739 26977
rect 12730 26961 12747 26966
rect 12667 26916 12679 26956
rect 12730 26900 12737 26961
rect 12752 26908 12755 26956
rect 12732 26851 12734 26900
rect 12731 26667 12738 26851
rect 12745 26841 12748 26851
rect 12756 26841 12758 26979
rect 12794 26915 12797 26925
rect 12804 26917 12806 26979
rect 12817 26977 12822 26979
rect 12826 26953 12833 26979
rect 12804 26893 12808 26917
rect 12755 26793 12758 26841
rect 12776 26833 12782 26841
rect 12732 26658 12734 26667
rect 12756 26658 12758 26793
rect 12788 26793 12794 26833
rect 12788 26667 12792 26793
rect 12602 26650 12612 26658
rect 12630 26650 12640 26658
rect 12662 26650 12670 26658
rect 12724 26650 12734 26658
rect 12752 26650 12762 26658
rect 12596 26642 12602 26650
rect 12624 26642 12630 26650
rect 12636 26639 12638 26650
rect 12670 26642 12678 26650
rect 12718 26642 12724 26650
rect 12732 26639 12734 26650
rect 12746 26642 12752 26650
rect 12756 26639 12758 26650
rect 12804 26639 12806 26893
rect 12808 26667 12814 26841
rect 12828 26833 12830 26953
rect 12841 26841 12844 26851
rect 12852 26841 12854 26979
rect 12900 26917 12903 26979
rect 12920 26972 12929 26979
rect 12924 26969 12928 26972
rect 12924 26953 12927 26969
rect 12887 26907 12892 26913
rect 12887 26903 12894 26907
rect 12900 26903 12904 26917
rect 12897 26893 12904 26903
rect 12897 26889 12902 26893
rect 12900 26843 12902 26889
rect 12917 26849 12921 26889
rect 12924 26849 12926 26953
rect 12833 26833 12841 26841
rect 12851 26833 12854 26841
rect 12815 26793 12824 26833
rect 12826 26793 12831 26833
rect 12835 26793 12841 26833
rect 12842 26793 12858 26833
rect 12826 26785 12833 26793
rect 12852 26785 12858 26793
rect 12828 26658 12830 26785
rect 12852 26658 12854 26785
rect 12862 26667 12868 26841
rect 12872 26833 12878 26841
rect 12884 26793 12890 26833
rect 12884 26667 12888 26793
rect 12900 26791 12910 26843
rect 12917 26839 12927 26849
rect 12929 26839 12936 26972
rect 12937 26953 12940 26963
rect 12948 26953 12950 26979
rect 13017 26964 13022 26979
rect 12947 26937 12950 26953
rect 12924 26833 12926 26839
rect 12911 26791 12917 26833
rect 12820 26650 12830 26658
rect 12848 26650 12856 26658
rect 12812 26642 12820 26650
rect 12828 26639 12830 26650
rect 12840 26642 12848 26650
rect 12852 26639 12854 26650
rect 12900 26639 12902 26791
rect 12919 26785 12926 26833
rect 12928 26785 12937 26839
rect 12948 26833 12950 26937
rect 13007 26903 13012 26913
rect 13020 26903 13022 26964
rect 13036 26945 13039 26979
rect 13044 26969 13046 26979
rect 13044 26945 13048 26969
rect 12963 26895 12965 26899
rect 12973 26881 12975 26895
rect 13017 26889 13022 26903
rect 12938 26791 12944 26833
rect 12946 26785 12953 26833
rect 12955 26791 12964 26843
rect 12977 26791 12981 26849
rect 13020 26841 13022 26889
rect 13036 26851 13039 26929
rect 13033 26841 13039 26851
rect 13044 26891 13046 26945
rect 13049 26891 13053 26979
rect 13044 26841 13053 26891
rect 13063 26841 13066 26979
rect 12994 26831 12998 26839
rect 13020 26831 13029 26841
rect 13043 26831 13056 26841
rect 13068 26831 13070 26979
rect 13112 26978 13118 26979
rect 13105 26841 13108 26851
rect 13116 26841 13118 26978
rect 13084 26833 13088 26841
rect 13112 26833 13118 26841
rect 13138 26833 13142 26841
rect 12982 26791 12993 26831
rect 12995 26791 12998 26831
rect 13018 26793 13029 26831
rect 13031 26793 13034 26831
rect 13036 26793 13047 26831
rect 13049 26793 13056 26831
rect 13058 26793 13061 26831
rect 12924 26658 12926 26785
rect 12929 26783 12936 26785
rect 12948 26658 12950 26785
rect 12977 26783 12980 26791
rect 13004 26667 13008 26791
rect 12914 26650 12926 26658
rect 12942 26650 12952 26658
rect 12974 26650 12982 26658
rect 13002 26650 13016 26658
rect 12908 26642 12914 26650
rect 12924 26639 12926 26650
rect 12936 26642 12942 26650
rect 12948 26639 12950 26650
rect 12982 26642 12990 26650
rect 13016 26642 13018 26650
rect 13020 26639 13022 26793
rect 13036 26785 13043 26793
rect 13044 26658 13046 26793
rect 13063 26785 13070 26831
rect 13072 26793 13074 26831
rect 13068 26658 13070 26785
rect 13094 26667 13098 26833
rect 13099 26793 13110 26833
rect 13112 26793 13119 26833
rect 13121 26793 13124 26833
rect 13126 26793 13137 26833
rect 13139 26793 13142 26833
rect 13032 26650 13046 26658
rect 13060 26650 13072 26658
rect 13092 26650 13100 26658
rect 13030 26642 13032 26650
rect 13044 26639 13046 26650
rect 13058 26642 13060 26650
rect 13068 26639 13070 26650
rect 13072 26642 13074 26650
rect 13100 26642 13108 26650
rect 13116 26639 13118 26793
rect 13119 26785 13124 26793
rect 13148 26667 13152 26793
rect 13188 26658 13190 26979
rect 13192 26970 13193 26979
rect 13193 26919 13200 26967
rect 13219 26667 13228 26843
rect 13120 26650 13128 26658
rect 13182 26650 13192 26658
rect 13210 26650 13220 26658
rect 13242 26650 13250 26658
rect 13270 26650 13282 26658
rect 13284 26650 13286 26979
rect 13292 26964 13294 26969
rect 13287 26916 13294 26964
rect 13295 26916 13311 26959
rect 13310 26911 13311 26916
rect 13332 26658 13334 26979
rect 13363 26916 13375 26956
rect 13428 26658 13430 26979
rect 13524 26969 13528 26979
rect 13432 26919 13448 26956
rect 13450 26911 13451 26956
rect 13459 26667 13461 26966
rect 13524 26959 13534 26969
rect 13524 26913 13526 26959
rect 13511 26911 13526 26913
rect 13511 26903 13516 26911
rect 13524 26903 13526 26911
rect 13535 26911 13550 26959
rect 13561 26953 13564 26963
rect 13572 26953 13574 26979
rect 13571 26937 13574 26953
rect 13535 26903 13544 26911
rect 13521 26889 13526 26903
rect 13298 26650 13310 26658
rect 13326 26650 13338 26658
rect 13358 26650 13366 26658
rect 13422 26650 13430 26658
rect 13450 26650 13458 26658
rect 13482 26650 13490 26658
rect 13510 26650 13522 26658
rect 13524 26650 13526 26889
rect 13542 26839 13551 26849
rect 13552 26667 13561 26839
rect 13572 26658 13574 26937
rect 13631 26903 13636 26913
rect 13644 26903 13646 26979
rect 13667 26977 13680 26979
rect 13667 26972 13670 26977
rect 13587 26895 13589 26899
rect 13597 26881 13599 26895
rect 13641 26889 13646 26903
rect 13601 26791 13605 26849
rect 13644 26841 13646 26889
rect 13668 26969 13670 26972
rect 13668 26945 13672 26969
rect 13618 26831 13622 26839
rect 13606 26791 13617 26831
rect 13619 26791 13622 26831
rect 13644 26791 13654 26841
rect 13662 26839 13665 26849
rect 13668 26831 13670 26945
rect 13673 26839 13680 26972
rect 13681 26953 13684 26963
rect 13692 26953 13694 26979
rect 13691 26937 13694 26953
rect 13655 26791 13661 26831
rect 13601 26783 13604 26791
rect 13628 26667 13632 26791
rect 13538 26650 13550 26658
rect 13566 26650 13578 26658
rect 13598 26650 13606 26658
rect 13626 26650 13642 26658
rect 13128 26642 13136 26650
rect 13176 26642 13182 26650
rect 13188 26639 13190 26650
rect 13204 26642 13210 26650
rect 13250 26642 13258 26650
rect 13282 26642 13286 26650
rect 13310 26642 13314 26650
rect 13284 26639 13286 26642
rect 13332 26639 13334 26650
rect 13338 26642 13342 26650
rect 13366 26642 13374 26650
rect 13414 26642 13422 26650
rect 13428 26639 13430 26650
rect 13442 26642 13450 26650
rect 13490 26642 13498 26650
rect 13522 26642 13526 26650
rect 13550 26642 13554 26650
rect 13524 26639 13526 26642
rect 13572 26639 13574 26650
rect 13578 26642 13582 26650
rect 13606 26642 13614 26650
rect 13644 26639 13646 26791
rect 13663 26783 13670 26831
rect 13672 26783 13681 26839
rect 13692 26831 13694 26937
rect 13707 26895 13709 26899
rect 13717 26881 13719 26895
rect 13682 26791 13688 26831
rect 13690 26783 13697 26831
rect 13699 26791 13708 26841
rect 13721 26791 13725 26849
rect 13738 26831 13742 26839
rect 13726 26791 13737 26831
rect 13739 26791 13742 26831
rect 13721 26783 13724 26791
rect 13668 26658 13670 26783
rect 13692 26658 13694 26783
rect 13748 26667 13752 26791
rect 13658 26650 13670 26658
rect 13686 26650 13698 26658
rect 13718 26650 13726 26658
rect 13654 26642 13658 26650
rect 13668 26639 13670 26650
rect 13682 26642 13686 26650
rect 13692 26639 13694 26650
rect 13726 26642 13734 26650
rect 13764 26639 13766 26979
rect 13788 26977 13802 26979
rect 13788 26969 13790 26977
rect 13787 26961 13792 26969
rect 13788 26955 13792 26961
rect 13786 26929 13793 26955
rect 13768 26667 13774 26841
rect 13788 26831 13790 26929
rect 13801 26841 13804 26851
rect 13812 26841 13814 26979
rect 13850 26915 13853 26925
rect 13860 26917 13862 26979
rect 13873 26977 13878 26979
rect 13882 26953 13889 26979
rect 13860 26893 13864 26917
rect 13793 26831 13801 26841
rect 13811 26831 13814 26841
rect 13775 26793 13784 26831
rect 13786 26793 13791 26831
rect 13795 26793 13801 26831
rect 13802 26793 13818 26831
rect 13786 26785 13793 26793
rect 13812 26785 13818 26793
rect 13788 26658 13790 26785
rect 13812 26658 13814 26785
rect 13822 26667 13828 26841
rect 13832 26833 13838 26841
rect 13844 26793 13850 26833
rect 13844 26667 13848 26793
rect 13780 26650 13790 26658
rect 13808 26650 13818 26658
rect 13774 26642 13780 26650
rect 13788 26639 13790 26650
rect 13802 26642 13808 26650
rect 13812 26639 13814 26650
rect 13860 26639 13862 26893
rect 13864 26667 13870 26841
rect 13884 26833 13886 26953
rect 13897 26841 13900 26851
rect 13908 26841 13910 26979
rect 13956 26917 13958 26979
rect 13959 26953 13975 26964
rect 13959 26917 13965 26953
rect 13956 26916 13965 26917
rect 13985 26916 13987 26964
rect 13956 26893 13960 26916
rect 13889 26833 13897 26841
rect 13907 26833 13910 26841
rect 13871 26793 13880 26833
rect 13882 26793 13887 26833
rect 13891 26793 13897 26833
rect 13898 26793 13914 26833
rect 13882 26785 13889 26793
rect 13908 26785 13914 26793
rect 13884 26658 13886 26785
rect 13908 26658 13910 26785
rect 13918 26667 13924 26841
rect 13928 26833 13934 26841
rect 13940 26793 13946 26833
rect 13940 26667 13944 26793
rect 13876 26650 13886 26658
rect 13904 26650 13912 26658
rect 13868 26642 13876 26650
rect 13884 26639 13886 26650
rect 13896 26642 13904 26650
rect 13908 26639 13910 26650
rect 13956 26639 13958 26893
rect 14004 26658 14006 26979
rect 14035 26916 14047 26956
rect 14100 26658 14102 26979
rect 14193 26969 14200 26979
rect 14104 26919 14120 26956
rect 14122 26911 14123 26956
rect 14131 26667 14133 26966
rect 14193 26959 14203 26969
rect 14212 26959 14215 26979
rect 14183 26903 14188 26913
rect 14196 26903 14198 26959
rect 14207 26911 14219 26959
rect 14207 26903 14215 26911
rect 14193 26889 14198 26903
rect 13970 26650 13980 26658
rect 13998 26650 14008 26658
rect 14030 26650 14038 26658
rect 14094 26650 14102 26658
rect 14122 26650 14130 26658
rect 14154 26650 14162 26658
rect 14182 26650 14192 26658
rect 14196 26650 14198 26889
rect 14244 26658 14246 26979
rect 14288 26978 14294 26979
rect 14281 26841 14284 26851
rect 14292 26841 14294 26978
rect 14450 26882 14457 26979
rect 14500 26976 14503 26979
rect 14576 26968 14579 26979
rect 14617 26970 14620 26979
rect 14635 26978 14721 26979
rect 14670 26960 14673 26961
rect 14480 26952 14486 26960
rect 14493 26952 14507 26960
rect 14567 26952 14576 26953
rect 14636 26952 14638 26960
rect 14645 26952 14679 26960
rect 14500 26950 14503 26952
rect 14576 26950 14579 26952
rect 14486 26902 14493 26950
rect 14496 26902 14497 26942
rect 14481 26894 14490 26902
rect 14500 26894 14507 26942
rect 14518 26902 14525 26950
rect 14569 26947 14583 26950
rect 14576 26942 14583 26947
rect 14557 26902 14560 26942
rect 14512 26894 14557 26902
rect 14562 26894 14569 26942
rect 14577 26894 14583 26942
rect 14634 26902 14636 26942
rect 14638 26902 14645 26950
rect 14665 26947 14686 26950
rect 14679 26942 14686 26947
rect 14732 26942 14736 26978
rect 14653 26902 14654 26942
rect 14603 26894 14610 26902
rect 14656 26894 14663 26942
rect 14667 26902 14671 26942
rect 14679 26902 14683 26942
rect 14710 26902 14711 26942
rect 14686 26894 14693 26902
rect 14719 26894 14726 26942
rect 14500 26882 14503 26894
rect 14576 26892 14583 26894
rect 14576 26882 14579 26892
rect 14440 26874 14512 26882
rect 14557 26874 14634 26882
rect 14450 26872 14457 26874
rect 14460 26856 14464 26862
rect 14260 26833 14264 26841
rect 14288 26833 14294 26841
rect 14314 26833 14318 26841
rect 14270 26667 14274 26833
rect 14275 26793 14286 26833
rect 14288 26793 14295 26833
rect 14297 26793 14300 26833
rect 14302 26793 14313 26833
rect 14315 26793 14318 26833
rect 14210 26650 14220 26658
rect 14238 26650 14248 26658
rect 14268 26650 14276 26658
rect 13964 26642 13970 26650
rect 13992 26642 13998 26650
rect 14004 26639 14006 26650
rect 14038 26642 14046 26650
rect 14086 26642 14094 26650
rect 14100 26639 14102 26650
rect 14114 26642 14122 26650
rect 14162 26642 14170 26650
rect 14192 26642 14198 26650
rect 14220 26642 14226 26650
rect 14196 26639 14198 26642
rect 14244 26639 14246 26650
rect 14248 26642 14254 26650
rect 14276 26642 14284 26650
rect 14292 26639 14294 26793
rect 14295 26785 14300 26793
rect 14324 26667 14328 26793
rect 14348 26667 14350 26843
rect 14376 26824 14381 26833
rect 14351 26785 14364 26824
rect 14374 26785 14376 26824
rect 14378 26785 14381 26824
rect 14384 26785 14394 26824
rect 14450 26816 14457 26856
rect 14500 26841 14503 26874
rect 14504 26864 14507 26874
rect 14514 26854 14517 26864
rect 14514 26848 14530 26854
rect 14558 26848 14570 26854
rect 14472 26824 14476 26834
rect 14486 26826 14508 26834
rect 14486 26825 14502 26826
rect 14576 26824 14579 26874
rect 14602 26854 14724 26859
rect 14628 26839 14646 26846
rect 14583 26826 14603 26834
rect 14732 26826 14736 26894
rect 14482 26820 14500 26824
rect 14369 26777 14374 26785
rect 14442 26768 14449 26816
rect 14482 26776 14488 26820
rect 14518 26776 14525 26824
rect 14576 26816 14584 26824
rect 14638 26816 14645 26824
rect 14558 26776 14560 26816
rect 14460 26768 14476 26775
rect 14482 26768 14486 26776
rect 14562 26768 14569 26816
rect 14577 26768 14584 26816
rect 14620 26777 14628 26816
rect 14620 26776 14636 26777
rect 14450 26705 14457 26768
rect 14576 26765 14584 26768
rect 14603 26765 14610 26776
rect 14628 26768 14636 26776
rect 14656 26768 14663 26816
rect 14665 26776 14669 26816
rect 14679 26776 14681 26824
rect 14686 26768 14693 26816
rect 14698 26778 14704 26816
rect 14732 26778 14739 26826
rect 14741 26778 14745 26816
rect 14719 26768 14726 26778
rect 14802 26771 14806 26818
rect 14875 26815 14878 26841
rect 14886 26815 14892 26979
rect 14916 26824 14923 26979
rect 14992 26932 14999 26979
rect 15052 26948 15061 26979
rect 15088 26947 15096 26956
rect 15087 26942 15096 26947
rect 15038 26934 15040 26939
rect 15050 26934 15052 26939
rect 15052 26929 15060 26934
rect 15062 26924 15070 26929
rect 15084 26921 15086 26934
rect 15094 26932 15103 26942
rect 15113 26932 15120 26979
rect 15121 26955 15124 26965
rect 15132 26955 15134 26979
rect 15104 26931 15113 26932
rect 15128 26929 15130 26942
rect 15131 26939 15134 26955
rect 15172 26948 15181 26979
rect 15228 26971 15230 26979
rect 15227 26961 15232 26971
rect 15248 26961 15254 26979
rect 15228 26957 15232 26961
rect 14820 26783 14821 26813
rect 14867 26805 14869 26815
rect 14886 26805 14893 26815
rect 14906 26805 14913 26824
rect 14929 26823 14941 26824
rect 14928 26807 14941 26823
rect 14877 26789 14879 26805
rect 14896 26789 14913 26805
rect 14802 26770 14819 26771
rect 14688 26767 14691 26768
rect 14732 26767 14736 26768
rect 14464 26747 14500 26755
rect 14576 26753 14579 26765
rect 14886 26763 14892 26789
rect 14898 26776 14913 26789
rect 14933 26776 14940 26807
rect 14965 26789 14969 26837
rect 14992 26826 14999 26916
rect 15059 26883 15065 26909
rect 15084 26908 15086 26911
rect 15095 26847 15104 26911
rect 14974 26789 14981 26816
rect 14983 26781 14990 26816
rect 14552 26747 14600 26753
rect 14658 26747 14669 26755
rect 14499 26737 14500 26747
rect 14524 26745 14525 26747
rect 14518 26737 14525 26745
rect 14576 26743 14579 26747
rect 14450 26697 14466 26705
rect 14440 26685 14448 26695
rect 14450 26689 14459 26697
rect 14474 26687 14476 26715
rect 14499 26689 14507 26737
rect 14524 26697 14525 26737
rect 14545 26689 14552 26737
rect 14562 26727 14578 26737
rect 14638 26735 14645 26745
rect 14688 26735 14694 26755
rect 14702 26737 14711 26745
rect 14714 26737 14721 26755
rect 14766 26747 14783 26755
rect 14793 26747 14806 26755
rect 14804 26746 14806 26747
rect 14638 26719 14654 26735
rect 14616 26693 14622 26699
rect 14714 26697 14723 26737
rect 14776 26697 14787 26737
rect 14805 26697 14806 26746
rect 14859 26737 14865 26755
rect 14871 26747 14879 26759
rect 14916 26755 14923 26776
rect 14992 26768 15000 26826
rect 15001 26789 15008 26816
rect 15010 26781 15017 26816
rect 15019 26789 15027 26826
rect 15040 26819 15045 26847
rect 15095 26837 15105 26847
rect 15113 26837 15120 26916
rect 15132 26885 15134 26939
rect 15158 26934 15160 26939
rect 15170 26934 15172 26939
rect 15172 26929 15180 26934
rect 15226 26931 15233 26957
rect 15182 26924 15190 26929
rect 15139 26911 15148 26919
rect 15139 26885 15141 26901
rect 15132 26861 15141 26885
rect 15179 26883 15185 26909
rect 15204 26908 15206 26911
rect 15058 26829 15062 26837
rect 15074 26829 15084 26837
rect 15041 26789 15045 26819
rect 15046 26789 15057 26829
rect 15059 26789 15062 26829
rect 15086 26827 15093 26837
rect 15085 26789 15094 26827
rect 15095 26789 15101 26829
rect 15041 26781 15044 26789
rect 14882 26751 14906 26755
rect 14913 26751 14924 26755
rect 14882 26747 14895 26751
rect 14871 26745 14881 26747
rect 14886 26745 14892 26747
rect 14916 26745 14923 26751
rect 14934 26745 14941 26747
rect 14875 26742 14886 26745
rect 14893 26742 14900 26745
rect 14875 26737 14884 26742
rect 14905 26737 14914 26745
rect 14933 26737 14941 26745
rect 14947 26737 14951 26751
rect 14852 26697 14855 26737
rect 14857 26697 14864 26737
rect 14868 26697 14872 26737
rect 14875 26697 14882 26737
rect 14887 26697 14894 26737
rect 14898 26697 14903 26737
rect 14906 26697 14913 26737
rect 14915 26697 14924 26737
rect 14925 26697 14931 26737
rect 14933 26697 14940 26737
rect 14612 26689 14616 26693
rect 14678 26685 14684 26695
rect 14714 26689 14721 26697
rect 14852 26689 14872 26697
rect 14886 26689 14893 26697
rect 14915 26689 14923 26697
rect 14944 26689 14951 26737
rect 14992 26689 15000 26747
rect 14450 26677 14458 26685
rect 14688 26677 14694 26685
rect 14918 26677 14921 26689
rect 14450 26669 14566 26677
rect 14688 26669 14695 26677
rect 14711 26669 14729 26677
rect 14745 26669 14760 26677
rect 14918 26669 14925 26677
rect 14941 26669 14987 26677
rect 14992 26669 14997 26689
rect 15068 26667 15072 26789
rect 15103 26781 15110 26829
rect 15112 26781 15121 26837
rect 15132 26829 15134 26861
rect 15122 26789 15128 26829
rect 15130 26781 15137 26829
rect 15139 26789 15148 26839
rect 15160 26819 15165 26847
rect 15208 26839 15213 26841
rect 15178 26829 15182 26837
rect 15161 26789 15165 26819
rect 15166 26789 15177 26829
rect 15179 26789 15182 26829
rect 15161 26781 15164 26789
rect 14296 26650 14304 26658
rect 14358 26650 14368 26658
rect 14386 26650 14396 26658
rect 14418 26650 14426 26658
rect 14446 26650 14454 26658
rect 14474 26650 14482 26658
rect 14502 26650 14510 26658
rect 14513 26656 14526 26658
rect 14530 26650 14538 26658
rect 14558 26650 14566 26658
rect 14571 26656 14582 26658
rect 14586 26650 14594 26658
rect 14614 26650 14622 26658
rect 14642 26650 14650 26658
rect 14670 26650 14678 26658
rect 14698 26650 14706 26658
rect 14726 26656 14744 26658
rect 14726 26650 14734 26656
rect 14782 26650 14788 26661
rect 14810 26650 14816 26661
rect 14852 26653 14860 26661
rect 14864 26653 14872 26661
rect 14880 26653 14888 26661
rect 14892 26653 14900 26661
rect 14908 26653 14916 26661
rect 14920 26653 14928 26661
rect 14936 26653 14944 26661
rect 15132 26658 15134 26781
rect 15188 26667 15192 26789
rect 15208 26667 15214 26839
rect 15228 26829 15230 26931
rect 15252 26901 15254 26961
rect 15290 26915 15293 26925
rect 15300 26917 15302 26979
rect 15313 26977 15318 26979
rect 15322 26953 15329 26979
rect 15252 26885 15260 26901
rect 15300 26893 15304 26917
rect 15252 26861 15261 26885
rect 15241 26841 15244 26851
rect 15252 26841 15254 26861
rect 15233 26839 15240 26841
rect 15233 26829 15241 26839
rect 15251 26829 15254 26841
rect 15215 26793 15224 26829
rect 15226 26793 15231 26829
rect 15235 26793 15241 26829
rect 15242 26793 15258 26829
rect 15226 26785 15233 26793
rect 15252 26785 15258 26793
rect 15228 26658 15230 26785
rect 15252 26658 15254 26785
rect 15262 26667 15268 26839
rect 15272 26833 15278 26841
rect 15284 26793 15290 26833
rect 15284 26667 15288 26793
rect 14966 26653 14976 26658
rect 14982 26653 14992 26658
rect 14994 26653 15004 26658
rect 15010 26653 15020 26658
rect 14864 26652 14880 26653
rect 14892 26652 14908 26653
rect 14920 26652 14936 26653
rect 14948 26652 14956 26653
rect 14966 26652 14982 26653
rect 14994 26652 15010 26653
rect 15022 26652 15032 26658
rect 14304 26642 14312 26650
rect 14352 26642 14358 26650
rect 14380 26642 14386 26650
rect 14426 26642 14434 26650
rect 14454 26642 14462 26650
rect 14482 26642 14490 26650
rect 14510 26642 14518 26650
rect 14538 26642 14546 26650
rect 14566 26642 14574 26650
rect 14594 26642 14602 26650
rect 14622 26642 14630 26650
rect 14650 26642 14658 26650
rect 14678 26642 14686 26650
rect 14706 26642 14714 26650
rect 14734 26642 14742 26650
rect 14788 26645 14798 26650
rect 14816 26645 14826 26650
rect 14872 26645 14880 26652
rect 14900 26645 14908 26652
rect 14928 26645 14936 26652
rect 14976 26642 14982 26652
rect 15004 26642 15010 26652
rect 15042 26650 15050 26658
rect 15070 26650 15086 26658
rect 15102 26650 15114 26658
rect 15130 26650 15142 26658
rect 15162 26650 15170 26658
rect 15190 26650 15204 26658
rect 15220 26650 15232 26658
rect 15248 26650 15260 26658
rect 15050 26642 15058 26650
rect 15098 26642 15102 26650
rect 15126 26642 15130 26650
rect 14424 26639 14460 26642
rect 14810 26639 14844 26641
rect 15132 26639 15134 26650
rect 15170 26642 15178 26650
rect 15204 26642 15206 26650
rect 15218 26642 15220 26650
rect 15228 26639 15230 26650
rect 15232 26642 15234 26650
rect 15246 26642 15248 26650
rect 15252 26639 15254 26650
rect 15260 26642 15262 26650
rect 15300 26639 15302 26893
rect 15304 26667 15310 26841
rect 15324 26833 15326 26953
rect 15337 26841 15340 26851
rect 15348 26841 15350 26979
rect 15386 26915 15389 26925
rect 15396 26917 15398 26979
rect 15409 26977 15414 26979
rect 15418 26953 15425 26979
rect 15396 26893 15400 26917
rect 15329 26833 15337 26841
rect 15347 26833 15350 26841
rect 15311 26793 15320 26833
rect 15322 26793 15327 26833
rect 15331 26793 15337 26833
rect 15338 26793 15354 26833
rect 15322 26785 15329 26793
rect 15348 26785 15354 26793
rect 15324 26658 15326 26785
rect 15348 26658 15350 26785
rect 15358 26667 15364 26841
rect 15368 26833 15374 26841
rect 15380 26793 15386 26833
rect 15380 26667 15384 26793
rect 15316 26650 15326 26658
rect 15344 26650 15352 26658
rect 15308 26642 15316 26650
rect 15324 26639 15326 26650
rect 15336 26642 15344 26650
rect 15348 26639 15350 26650
rect 15396 26639 15398 26893
rect 15400 26667 15406 26841
rect 15420 26833 15422 26953
rect 15433 26841 15436 26851
rect 15444 26841 15446 26979
rect 15480 26956 15485 26966
rect 15492 26956 15495 26979
rect 15490 26953 15504 26956
rect 15490 26942 15495 26953
rect 15492 26917 15495 26942
rect 15521 26932 15528 26979
rect 15529 26955 15532 26965
rect 15540 26955 15542 26979
rect 15539 26939 15542 26955
rect 15580 26948 15589 26979
rect 15636 26971 15638 26979
rect 15635 26961 15640 26971
rect 15656 26961 15662 26979
rect 15636 26957 15640 26961
rect 15492 26893 15496 26917
rect 15425 26833 15433 26841
rect 15443 26833 15446 26841
rect 15407 26793 15416 26833
rect 15418 26793 15423 26833
rect 15427 26793 15433 26833
rect 15434 26793 15450 26833
rect 15418 26785 15425 26793
rect 15444 26785 15450 26793
rect 15420 26658 15422 26785
rect 15444 26658 15446 26785
rect 15454 26667 15460 26841
rect 15464 26833 15470 26841
rect 15492 26837 15494 26893
rect 15509 26847 15512 26893
rect 15509 26837 15519 26847
rect 15521 26837 15528 26916
rect 15482 26833 15501 26837
rect 15476 26793 15482 26833
rect 15492 26827 15501 26833
rect 15476 26667 15480 26793
rect 15492 26789 15502 26827
rect 15503 26789 15509 26833
rect 15412 26650 15422 26658
rect 15440 26650 15448 26658
rect 15404 26642 15412 26650
rect 15420 26639 15422 26650
rect 15432 26642 15440 26650
rect 15444 26639 15446 26650
rect 15492 26639 15494 26789
rect 15511 26785 15518 26833
rect 15520 26785 15529 26837
rect 15540 26833 15542 26939
rect 15566 26934 15568 26939
rect 15578 26934 15580 26939
rect 15580 26929 15588 26934
rect 15634 26931 15641 26957
rect 15590 26924 15598 26929
rect 15587 26883 15593 26909
rect 15612 26908 15614 26911
rect 15530 26789 15536 26833
rect 15538 26785 15545 26833
rect 15547 26789 15556 26843
rect 15568 26819 15573 26847
rect 15616 26839 15621 26841
rect 15586 26829 15590 26837
rect 15569 26789 15573 26819
rect 15574 26789 15585 26829
rect 15587 26789 15590 26829
rect 15521 26781 15528 26785
rect 15540 26658 15542 26785
rect 15569 26781 15572 26789
rect 15596 26667 15600 26789
rect 15616 26667 15622 26839
rect 15636 26829 15638 26931
rect 15660 26901 15662 26961
rect 15698 26915 15701 26925
rect 15708 26917 15710 26979
rect 15721 26977 15726 26979
rect 15730 26953 15737 26979
rect 15660 26885 15668 26901
rect 15708 26893 15712 26917
rect 15660 26861 15669 26885
rect 15649 26841 15652 26851
rect 15660 26841 15662 26861
rect 15641 26839 15648 26841
rect 15641 26829 15649 26839
rect 15659 26829 15662 26841
rect 15623 26793 15632 26829
rect 15634 26793 15639 26829
rect 15643 26793 15649 26829
rect 15650 26793 15666 26829
rect 15634 26785 15641 26793
rect 15660 26785 15666 26793
rect 15636 26658 15638 26785
rect 15660 26658 15662 26785
rect 15670 26667 15676 26839
rect 15680 26833 15686 26841
rect 15692 26793 15698 26833
rect 15692 26667 15696 26793
rect 15510 26650 15516 26658
rect 15538 26650 15544 26658
rect 15570 26650 15578 26658
rect 15598 26650 15612 26658
rect 15628 26650 15640 26658
rect 15656 26650 15668 26658
rect 15500 26642 15510 26650
rect 15528 26642 15538 26650
rect 15540 26639 15542 26650
rect 15578 26642 15586 26650
rect 15612 26642 15614 26650
rect 15626 26642 15628 26650
rect 15636 26639 15638 26650
rect 15640 26642 15642 26650
rect 15654 26642 15656 26650
rect 15660 26639 15662 26650
rect 15668 26642 15670 26650
rect 15708 26639 15710 26893
rect 15712 26667 15718 26841
rect 15732 26833 15734 26953
rect 15745 26841 15748 26851
rect 15756 26841 15758 26979
rect 15794 26915 15797 26925
rect 15804 26917 15806 26979
rect 15817 26977 15822 26979
rect 15826 26953 15833 26979
rect 15804 26893 15808 26917
rect 15737 26833 15745 26841
rect 15755 26833 15758 26841
rect 15719 26793 15728 26833
rect 15730 26793 15735 26833
rect 15739 26793 15745 26833
rect 15746 26793 15762 26833
rect 15730 26785 15737 26793
rect 15756 26785 15762 26793
rect 15732 26658 15734 26785
rect 15756 26658 15758 26785
rect 15766 26667 15772 26841
rect 15776 26833 15782 26841
rect 15788 26793 15794 26833
rect 15788 26667 15792 26793
rect 15724 26650 15734 26658
rect 15752 26650 15760 26658
rect 15716 26642 15724 26650
rect 15732 26639 15734 26650
rect 15744 26642 15752 26650
rect 15756 26639 15758 26650
rect 15804 26639 15806 26893
rect 15808 26667 15814 26841
rect 15828 26833 15830 26953
rect 15841 26841 15844 26851
rect 15852 26841 15854 26979
rect 15890 26915 15893 26925
rect 15900 26917 15902 26979
rect 15913 26977 15918 26979
rect 15922 26953 15929 26979
rect 15900 26893 15904 26917
rect 15833 26833 15841 26841
rect 15851 26833 15854 26841
rect 15815 26793 15824 26833
rect 15826 26793 15831 26833
rect 15835 26793 15841 26833
rect 15842 26793 15858 26833
rect 15826 26785 15833 26793
rect 15852 26785 15858 26793
rect 15828 26658 15830 26785
rect 15852 26658 15854 26785
rect 15862 26667 15868 26841
rect 15872 26833 15878 26841
rect 15884 26793 15890 26833
rect 15884 26667 15888 26793
rect 15820 26650 15830 26658
rect 15848 26650 15856 26658
rect 15812 26642 15820 26650
rect 15828 26639 15830 26650
rect 15840 26642 15848 26650
rect 15852 26639 15854 26650
rect 15900 26639 15902 26893
rect 15904 26667 15910 26841
rect 15924 26833 15926 26953
rect 15937 26841 15940 26851
rect 15948 26841 15950 26979
rect 15986 26915 15989 26925
rect 15996 26917 15998 26979
rect 16009 26977 16014 26979
rect 16018 26953 16025 26979
rect 15996 26893 16000 26917
rect 15929 26833 15937 26841
rect 15947 26833 15950 26841
rect 15911 26793 15920 26833
rect 15922 26793 15927 26833
rect 15931 26793 15937 26833
rect 15938 26793 15954 26833
rect 15922 26785 15929 26793
rect 15948 26785 15954 26793
rect 15924 26658 15926 26785
rect 15948 26658 15950 26785
rect 15958 26667 15964 26841
rect 15968 26833 15974 26841
rect 15980 26793 15986 26833
rect 15980 26667 15984 26793
rect 15916 26650 15926 26658
rect 15944 26650 15952 26658
rect 15908 26642 15916 26650
rect 15924 26639 15926 26650
rect 15936 26642 15944 26650
rect 15948 26639 15950 26650
rect 15996 26639 15998 26893
rect 16000 26667 16006 26841
rect 16020 26833 16022 26953
rect 16033 26841 16036 26851
rect 16044 26841 16046 26979
rect 16080 26956 16085 26966
rect 16092 26956 16095 26979
rect 16090 26953 16104 26956
rect 16090 26942 16095 26953
rect 16092 26917 16095 26942
rect 16121 26932 16128 26979
rect 16129 26955 16132 26965
rect 16140 26955 16142 26979
rect 16139 26939 16142 26955
rect 16180 26948 16189 26979
rect 16236 26971 16238 26979
rect 16235 26961 16240 26971
rect 16256 26961 16262 26979
rect 16236 26957 16240 26961
rect 16092 26893 16096 26917
rect 16025 26833 16033 26841
rect 16043 26833 16046 26841
rect 16007 26793 16016 26833
rect 16018 26793 16023 26833
rect 16027 26793 16033 26833
rect 16034 26793 16050 26833
rect 16018 26785 16025 26793
rect 16044 26785 16050 26793
rect 16020 26658 16022 26785
rect 16044 26658 16046 26785
rect 16054 26667 16060 26841
rect 16064 26833 16070 26841
rect 16092 26837 16094 26893
rect 16109 26847 16112 26893
rect 16109 26837 16119 26847
rect 16121 26837 16128 26916
rect 16082 26833 16101 26837
rect 16076 26793 16082 26833
rect 16092 26827 16101 26833
rect 16076 26667 16080 26793
rect 16092 26789 16102 26827
rect 16103 26789 16109 26833
rect 16012 26650 16022 26658
rect 16040 26650 16048 26658
rect 16004 26642 16012 26650
rect 16020 26639 16022 26650
rect 16032 26642 16040 26650
rect 16044 26639 16046 26650
rect 16092 26639 16094 26789
rect 16111 26785 16118 26833
rect 16120 26785 16129 26837
rect 16140 26833 16142 26939
rect 16166 26934 16168 26939
rect 16178 26934 16180 26939
rect 16180 26929 16188 26934
rect 16234 26931 16241 26957
rect 16190 26924 16198 26929
rect 16187 26883 16193 26909
rect 16212 26908 16214 26911
rect 16130 26789 16136 26833
rect 16138 26785 16145 26833
rect 16147 26789 16156 26843
rect 16168 26819 16173 26847
rect 16216 26839 16221 26841
rect 16186 26829 16190 26837
rect 16169 26789 16173 26819
rect 16174 26789 16185 26829
rect 16187 26789 16190 26829
rect 16121 26781 16128 26785
rect 16140 26658 16142 26785
rect 16169 26781 16172 26789
rect 16196 26667 16200 26789
rect 16216 26667 16222 26839
rect 16236 26829 16238 26931
rect 16260 26901 16262 26961
rect 16298 26915 16301 26925
rect 16308 26917 16310 26979
rect 16321 26977 16326 26979
rect 16330 26953 16337 26979
rect 16260 26885 16268 26901
rect 16308 26893 16312 26917
rect 16260 26861 16269 26885
rect 16249 26841 16252 26851
rect 16260 26841 16262 26861
rect 16241 26839 16248 26841
rect 16241 26829 16249 26839
rect 16259 26829 16262 26841
rect 16223 26793 16232 26829
rect 16234 26793 16239 26829
rect 16243 26793 16249 26829
rect 16250 26793 16266 26829
rect 16234 26785 16241 26793
rect 16260 26785 16266 26793
rect 16236 26658 16238 26785
rect 16260 26658 16262 26785
rect 16270 26667 16276 26839
rect 16280 26833 16286 26841
rect 16292 26793 16298 26833
rect 16292 26667 16296 26793
rect 16110 26650 16116 26658
rect 16138 26650 16144 26658
rect 16170 26650 16178 26658
rect 16198 26650 16212 26658
rect 16228 26650 16240 26658
rect 16256 26650 16268 26658
rect 16100 26642 16110 26650
rect 16128 26642 16138 26650
rect 16140 26639 16142 26650
rect 16178 26642 16186 26650
rect 16212 26642 16214 26650
rect 16226 26642 16228 26650
rect 16236 26639 16238 26650
rect 16240 26642 16242 26650
rect 16254 26642 16256 26650
rect 16260 26639 16262 26650
rect 16268 26642 16270 26650
rect 16308 26639 16310 26893
rect 16312 26667 16318 26841
rect 16332 26833 16334 26953
rect 16345 26841 16348 26851
rect 16356 26841 16358 26979
rect 16404 26917 16406 26979
rect 16407 26953 16423 26964
rect 16407 26917 16413 26953
rect 16404 26916 16413 26917
rect 16433 26916 16435 26964
rect 16404 26893 16408 26916
rect 16337 26833 16345 26841
rect 16355 26833 16358 26841
rect 16319 26793 16328 26833
rect 16330 26793 16335 26833
rect 16339 26793 16345 26833
rect 16346 26793 16362 26833
rect 16330 26785 16337 26793
rect 16356 26785 16362 26793
rect 16332 26658 16334 26785
rect 16356 26658 16358 26785
rect 16366 26667 16372 26841
rect 16376 26833 16382 26841
rect 16388 26793 16394 26833
rect 16388 26667 16392 26793
rect 16324 26650 16334 26658
rect 16352 26650 16360 26658
rect 16316 26642 16324 26650
rect 16332 26639 16334 26650
rect 16344 26642 16352 26650
rect 16356 26639 16358 26650
rect 16404 26639 16406 26893
rect 16452 26658 16454 26979
rect 16546 26977 16553 26979
rect 16546 26966 16555 26977
rect 16546 26961 16563 26966
rect 16483 26916 16495 26956
rect 16546 26900 16553 26961
rect 16568 26908 16571 26956
rect 16548 26851 16550 26900
rect 16547 26667 16554 26851
rect 16561 26841 16564 26851
rect 16572 26841 16574 26979
rect 16610 26915 16613 26925
rect 16620 26917 16622 26979
rect 16633 26977 16638 26979
rect 16642 26953 16649 26979
rect 16620 26893 16624 26917
rect 16571 26793 16574 26841
rect 16592 26833 16598 26841
rect 16548 26658 16550 26667
rect 16572 26658 16574 26793
rect 16604 26793 16610 26833
rect 16604 26667 16608 26793
rect 16418 26650 16428 26658
rect 16446 26650 16456 26658
rect 16478 26650 16486 26658
rect 16540 26650 16550 26658
rect 16568 26650 16578 26658
rect 16412 26642 16418 26650
rect 16440 26642 16446 26650
rect 16452 26639 16454 26650
rect 16486 26642 16494 26650
rect 16534 26642 16540 26650
rect 16548 26639 16550 26650
rect 16562 26642 16568 26650
rect 16572 26639 16574 26650
rect 16620 26639 16622 26893
rect 16624 26667 16630 26841
rect 16644 26833 16646 26953
rect 16657 26841 16660 26851
rect 16668 26841 16670 26979
rect 16716 26917 16719 26979
rect 16736 26972 16745 26979
rect 16740 26969 16744 26972
rect 16740 26953 16743 26969
rect 16703 26907 16708 26913
rect 16703 26903 16710 26907
rect 16716 26903 16720 26917
rect 16713 26893 16720 26903
rect 16713 26889 16718 26893
rect 16716 26843 16718 26889
rect 16733 26849 16737 26889
rect 16740 26849 16742 26953
rect 16649 26833 16657 26841
rect 16667 26833 16670 26841
rect 16631 26793 16640 26833
rect 16642 26793 16647 26833
rect 16651 26793 16657 26833
rect 16658 26793 16674 26833
rect 16642 26785 16649 26793
rect 16668 26785 16674 26793
rect 16644 26658 16646 26785
rect 16668 26658 16670 26785
rect 16678 26667 16684 26841
rect 16688 26833 16694 26841
rect 16700 26793 16706 26833
rect 16700 26667 16704 26793
rect 16716 26791 16726 26843
rect 16733 26839 16743 26849
rect 16745 26839 16752 26972
rect 16753 26953 16756 26963
rect 16764 26953 16766 26979
rect 16763 26937 16766 26953
rect 16740 26833 16742 26839
rect 16727 26791 16733 26833
rect 16636 26650 16646 26658
rect 16664 26650 16672 26658
rect 16628 26642 16636 26650
rect 16644 26639 16646 26650
rect 16656 26642 16664 26650
rect 16668 26639 16670 26650
rect 16716 26639 16718 26791
rect 16735 26785 16742 26833
rect 16744 26785 16753 26839
rect 16764 26833 16766 26937
rect 16779 26895 16781 26899
rect 16789 26881 16791 26895
rect 16754 26791 16760 26833
rect 16762 26785 16769 26833
rect 16771 26791 16780 26843
rect 16793 26791 16797 26849
rect 16810 26831 16814 26839
rect 16798 26791 16809 26831
rect 16811 26791 16814 26831
rect 16740 26658 16742 26785
rect 16745 26783 16752 26785
rect 16764 26658 16766 26785
rect 16793 26783 16796 26791
rect 16820 26667 16824 26791
rect 16730 26650 16742 26658
rect 16758 26650 16768 26658
rect 16790 26650 16798 26658
rect 16818 26650 16834 26658
rect 16724 26642 16730 26650
rect 16740 26639 16742 26650
rect 16752 26642 16758 26650
rect 16764 26639 16766 26650
rect 16798 26642 16806 26650
rect 16836 26639 16838 26979
rect 16862 26977 16864 26979
rect 16839 26959 16845 26964
rect 16839 26945 16854 26959
rect 16839 26929 16855 26945
rect 16839 26916 16845 26929
rect 16865 26916 16867 26964
rect 16884 26658 16886 26979
rect 16978 26977 16985 26979
rect 16978 26966 16987 26977
rect 16978 26961 16995 26966
rect 16915 26916 16927 26956
rect 16978 26900 16985 26961
rect 17000 26908 17003 26956
rect 16980 26851 16982 26900
rect 16979 26667 16986 26851
rect 16993 26841 16996 26851
rect 17004 26841 17006 26979
rect 17040 26956 17045 26966
rect 17052 26956 17055 26979
rect 17050 26953 17064 26956
rect 17050 26942 17055 26953
rect 17052 26917 17055 26942
rect 17081 26932 17088 26979
rect 17089 26955 17092 26965
rect 17100 26955 17102 26979
rect 17099 26939 17102 26955
rect 17140 26948 17149 26979
rect 17196 26971 17198 26979
rect 17195 26961 17200 26971
rect 17216 26961 17222 26979
rect 17196 26957 17200 26961
rect 17052 26893 17056 26917
rect 17003 26793 17006 26841
rect 17024 26833 17030 26841
rect 17052 26837 17054 26893
rect 17069 26847 17072 26893
rect 17069 26837 17079 26847
rect 17081 26837 17088 26916
rect 17042 26833 17061 26837
rect 16980 26658 16982 26667
rect 17004 26658 17006 26793
rect 17036 26793 17042 26833
rect 17052 26827 17061 26833
rect 17036 26667 17040 26793
rect 17052 26789 17062 26827
rect 17063 26789 17069 26833
rect 16850 26650 16862 26658
rect 16878 26650 16890 26658
rect 16910 26650 16918 26658
rect 16972 26650 16982 26658
rect 17000 26650 17010 26658
rect 16846 26642 16850 26650
rect 16874 26642 16878 26650
rect 16884 26639 16886 26650
rect 16918 26642 16926 26650
rect 16966 26642 16972 26650
rect 16980 26639 16982 26650
rect 16994 26642 17000 26650
rect 17004 26639 17006 26650
rect 17052 26639 17054 26789
rect 17071 26785 17078 26833
rect 17080 26785 17089 26837
rect 17100 26833 17102 26939
rect 17126 26934 17128 26939
rect 17138 26934 17140 26939
rect 17140 26929 17148 26934
rect 17194 26931 17201 26957
rect 17150 26924 17158 26929
rect 17147 26883 17153 26909
rect 17172 26908 17174 26911
rect 17090 26789 17096 26833
rect 17098 26785 17105 26833
rect 17107 26789 17116 26843
rect 17128 26819 17133 26847
rect 17176 26839 17181 26841
rect 17146 26829 17150 26837
rect 17129 26789 17133 26819
rect 17134 26789 17145 26829
rect 17147 26789 17150 26829
rect 17081 26781 17088 26785
rect 17100 26658 17102 26785
rect 17129 26781 17132 26789
rect 17156 26667 17160 26789
rect 17176 26667 17182 26839
rect 17196 26829 17198 26931
rect 17220 26901 17222 26961
rect 17258 26915 17261 26925
rect 17268 26917 17270 26979
rect 17281 26977 17286 26979
rect 17290 26953 17297 26979
rect 17220 26885 17228 26901
rect 17268 26893 17272 26917
rect 17220 26861 17229 26885
rect 17209 26841 17212 26851
rect 17220 26841 17222 26861
rect 17201 26839 17208 26841
rect 17201 26829 17209 26839
rect 17219 26829 17222 26841
rect 17183 26793 17192 26829
rect 17194 26793 17199 26829
rect 17203 26793 17209 26829
rect 17210 26793 17226 26829
rect 17194 26785 17201 26793
rect 17220 26785 17226 26793
rect 17196 26658 17198 26785
rect 17220 26658 17222 26785
rect 17230 26667 17236 26839
rect 17240 26833 17246 26841
rect 17252 26793 17258 26833
rect 17252 26667 17256 26793
rect 17070 26650 17076 26658
rect 17098 26650 17104 26658
rect 17130 26650 17138 26658
rect 17158 26650 17172 26658
rect 17188 26650 17200 26658
rect 17216 26650 17228 26658
rect 17060 26642 17070 26650
rect 17088 26642 17098 26650
rect 17100 26639 17102 26650
rect 17138 26642 17146 26650
rect 17172 26642 17174 26650
rect 17186 26642 17188 26650
rect 17196 26639 17198 26650
rect 17200 26642 17202 26650
rect 17214 26642 17216 26650
rect 17220 26639 17222 26650
rect 17228 26642 17230 26650
rect 17268 26639 17270 26893
rect 17272 26667 17278 26841
rect 17292 26833 17294 26953
rect 17305 26841 17308 26851
rect 17316 26841 17318 26979
rect 17362 26893 17381 26902
rect 17474 26882 17481 26979
rect 17524 26976 17527 26979
rect 17600 26968 17603 26979
rect 17641 26970 17644 26979
rect 17659 26978 17745 26979
rect 17694 26960 17697 26961
rect 17504 26952 17510 26960
rect 17517 26952 17531 26960
rect 17591 26952 17600 26953
rect 17660 26952 17662 26960
rect 17669 26952 17703 26960
rect 17524 26950 17527 26952
rect 17600 26950 17603 26952
rect 17510 26902 17517 26950
rect 17520 26902 17521 26942
rect 17505 26894 17514 26902
rect 17524 26894 17531 26942
rect 17542 26902 17549 26950
rect 17593 26947 17607 26950
rect 17600 26942 17607 26947
rect 17581 26902 17584 26942
rect 17536 26894 17581 26902
rect 17586 26894 17593 26942
rect 17601 26894 17607 26942
rect 17658 26902 17660 26942
rect 17662 26902 17669 26950
rect 17689 26947 17710 26950
rect 17703 26942 17710 26947
rect 17756 26942 17760 26978
rect 17677 26902 17678 26942
rect 17627 26894 17634 26902
rect 17680 26894 17687 26942
rect 17691 26902 17695 26942
rect 17703 26902 17707 26942
rect 17734 26902 17735 26942
rect 17710 26894 17717 26902
rect 17743 26894 17750 26942
rect 17524 26882 17527 26894
rect 17600 26892 17607 26894
rect 17600 26882 17603 26892
rect 17464 26874 17536 26882
rect 17581 26874 17658 26882
rect 17474 26872 17481 26874
rect 17484 26856 17488 26862
rect 17297 26833 17305 26841
rect 17315 26833 17318 26841
rect 17279 26793 17288 26833
rect 17290 26793 17295 26833
rect 17299 26793 17305 26833
rect 17306 26793 17322 26833
rect 17290 26785 17297 26793
rect 17316 26785 17322 26793
rect 17292 26658 17294 26785
rect 17316 26658 17318 26785
rect 17326 26667 17332 26841
rect 17336 26833 17342 26841
rect 17348 26793 17354 26833
rect 17348 26667 17352 26793
rect 17372 26667 17374 26843
rect 17400 26824 17405 26833
rect 17375 26785 17388 26824
rect 17398 26785 17400 26824
rect 17402 26785 17405 26824
rect 17408 26785 17418 26824
rect 17474 26816 17481 26856
rect 17524 26841 17527 26874
rect 17528 26864 17531 26874
rect 17538 26854 17541 26864
rect 17538 26848 17554 26854
rect 17582 26848 17594 26854
rect 17496 26824 17500 26834
rect 17510 26826 17532 26834
rect 17510 26825 17526 26826
rect 17600 26824 17603 26874
rect 17626 26854 17748 26859
rect 17652 26839 17670 26846
rect 17607 26826 17627 26834
rect 17756 26826 17760 26894
rect 17506 26820 17524 26824
rect 17393 26777 17398 26785
rect 17466 26768 17473 26816
rect 17506 26776 17512 26820
rect 17542 26776 17549 26824
rect 17600 26816 17608 26824
rect 17662 26816 17669 26824
rect 17582 26776 17584 26816
rect 17484 26768 17500 26775
rect 17506 26768 17510 26776
rect 17586 26768 17593 26816
rect 17601 26768 17608 26816
rect 17644 26777 17652 26816
rect 17644 26776 17660 26777
rect 17474 26705 17481 26768
rect 17600 26765 17608 26768
rect 17627 26765 17634 26776
rect 17652 26768 17660 26776
rect 17680 26768 17687 26816
rect 17689 26776 17693 26816
rect 17703 26776 17705 26824
rect 17710 26768 17717 26816
rect 17722 26778 17728 26816
rect 17756 26778 17763 26826
rect 17765 26778 17769 26816
rect 17743 26768 17750 26778
rect 17826 26771 17830 26818
rect 17899 26815 17902 26841
rect 17910 26815 17916 26979
rect 17940 26824 17947 26979
rect 18081 26917 18087 26979
rect 18100 26969 18103 26979
rect 18108 26969 18112 26979
rect 18108 26953 18111 26969
rect 18071 26907 18076 26913
rect 18071 26903 18078 26907
rect 18081 26893 18088 26917
rect 18081 26889 18086 26893
rect 18084 26841 18086 26889
rect 18100 26891 18103 26953
rect 18100 26889 18105 26891
rect 18100 26851 18103 26889
rect 18108 26851 18110 26953
rect 18097 26841 18110 26851
rect 17844 26783 17845 26813
rect 17891 26805 17893 26815
rect 17910 26805 17917 26815
rect 17930 26805 17937 26824
rect 17953 26823 17965 26824
rect 17952 26807 17965 26823
rect 17901 26789 17903 26805
rect 17920 26789 17937 26805
rect 17826 26770 17843 26771
rect 17712 26767 17715 26768
rect 17756 26767 17760 26768
rect 17488 26747 17524 26755
rect 17600 26753 17603 26765
rect 17910 26763 17916 26789
rect 17922 26776 17937 26789
rect 17957 26776 17964 26807
rect 17992 26793 17993 26841
rect 18017 26826 18023 26841
rect 18056 26833 18062 26841
rect 18084 26833 18093 26841
rect 18101 26833 18110 26841
rect 18113 26841 18117 26979
rect 18127 26841 18130 26979
rect 18017 26816 18024 26826
rect 17998 26793 18008 26816
rect 18010 26793 18014 26816
rect 18016 26793 18017 26816
rect 18019 26793 18024 26816
rect 18025 26793 18035 26816
rect 18010 26785 18016 26793
rect 18037 26785 18041 26816
rect 17576 26747 17624 26753
rect 17682 26747 17693 26755
rect 17523 26737 17524 26747
rect 17548 26745 17549 26747
rect 17542 26737 17549 26745
rect 17600 26743 17603 26747
rect 17474 26697 17490 26705
rect 17464 26685 17472 26695
rect 17474 26689 17483 26697
rect 17498 26687 17500 26715
rect 17523 26689 17531 26737
rect 17548 26697 17549 26737
rect 17569 26689 17576 26737
rect 17586 26727 17602 26737
rect 17662 26735 17669 26745
rect 17712 26735 17718 26755
rect 17726 26737 17735 26745
rect 17738 26737 17745 26755
rect 17790 26747 17807 26755
rect 17817 26747 17830 26755
rect 17828 26746 17830 26747
rect 17662 26719 17678 26735
rect 17640 26693 17646 26699
rect 17738 26697 17747 26737
rect 17800 26697 17811 26737
rect 17829 26697 17830 26746
rect 17883 26737 17889 26755
rect 17895 26747 17903 26759
rect 17940 26755 17947 26776
rect 17906 26751 17930 26755
rect 17937 26751 17948 26755
rect 17906 26747 17919 26751
rect 17895 26745 17905 26747
rect 17910 26745 17916 26747
rect 17940 26745 17947 26751
rect 17958 26745 17965 26747
rect 17899 26742 17910 26745
rect 17917 26742 17924 26745
rect 17899 26737 17908 26742
rect 17929 26737 17938 26745
rect 17957 26737 17965 26745
rect 17971 26737 17975 26751
rect 17876 26697 17879 26737
rect 17881 26697 17888 26737
rect 17892 26697 17896 26737
rect 17899 26697 17906 26737
rect 17911 26697 17918 26737
rect 17922 26697 17927 26737
rect 17930 26697 17937 26737
rect 17939 26697 17948 26737
rect 17949 26697 17955 26737
rect 17957 26697 17964 26737
rect 17636 26689 17640 26693
rect 17702 26685 17708 26695
rect 17738 26689 17745 26697
rect 17876 26689 17896 26697
rect 17910 26689 17917 26697
rect 17939 26689 17947 26697
rect 17968 26689 17975 26737
rect 17992 26689 17994 26747
rect 17474 26677 17482 26685
rect 17712 26677 17718 26685
rect 17942 26677 17945 26689
rect 17474 26669 17590 26677
rect 17712 26669 17719 26677
rect 17735 26669 17753 26677
rect 17769 26669 17784 26677
rect 17942 26669 17949 26677
rect 17965 26669 17992 26677
rect 18008 26669 18011 26677
rect 18046 26667 18051 26826
rect 18068 26793 18074 26833
rect 18082 26793 18093 26833
rect 18095 26793 18098 26833
rect 18100 26793 18111 26833
rect 18113 26793 18120 26841
rect 18132 26833 18134 26979
rect 18176 26978 18182 26979
rect 18169 26841 18172 26851
rect 18180 26841 18182 26978
rect 18148 26833 18152 26841
rect 18176 26833 18182 26841
rect 18202 26833 18206 26841
rect 18122 26793 18125 26833
rect 18068 26667 18072 26793
rect 17284 26650 17294 26658
rect 17312 26650 17320 26658
rect 17382 26650 17388 26658
rect 17410 26650 17416 26658
rect 17442 26650 17450 26658
rect 17470 26650 17478 26658
rect 17498 26650 17506 26658
rect 17526 26650 17534 26658
rect 17537 26656 17550 26658
rect 17554 26650 17562 26658
rect 17582 26650 17590 26658
rect 17595 26656 17606 26658
rect 17610 26650 17618 26658
rect 17638 26650 17646 26658
rect 17666 26650 17674 26658
rect 17694 26650 17702 26658
rect 17722 26650 17730 26658
rect 17750 26656 17768 26658
rect 17750 26650 17758 26656
rect 17806 26650 17812 26661
rect 17834 26650 17840 26661
rect 17876 26653 17884 26661
rect 17888 26653 17896 26661
rect 17904 26653 17912 26661
rect 17916 26653 17924 26661
rect 17932 26653 17940 26661
rect 17944 26653 17952 26661
rect 17960 26653 17968 26661
rect 17972 26653 17988 26658
rect 18004 26653 18016 26658
rect 18032 26653 18044 26658
rect 17888 26652 17904 26653
rect 17916 26652 17932 26653
rect 17944 26652 17960 26653
rect 17972 26652 17980 26653
rect 17276 26642 17284 26650
rect 17292 26639 17294 26650
rect 17304 26642 17312 26650
rect 17316 26639 17318 26650
rect 17372 26642 17382 26650
rect 17400 26642 17410 26650
rect 17450 26642 17458 26650
rect 17478 26642 17486 26650
rect 17506 26642 17514 26650
rect 17534 26642 17542 26650
rect 17562 26642 17570 26650
rect 17590 26642 17598 26650
rect 17618 26642 17626 26650
rect 17646 26642 17654 26650
rect 17674 26642 17682 26650
rect 17702 26642 17710 26650
rect 17730 26642 17738 26650
rect 17758 26642 17766 26650
rect 17812 26645 17822 26650
rect 17840 26645 17850 26650
rect 17896 26645 17904 26652
rect 17924 26645 17932 26652
rect 17952 26645 17960 26652
rect 18000 26642 18004 26653
rect 18028 26642 18032 26653
rect 18064 26650 18080 26658
rect 17448 26639 17484 26642
rect 17834 26639 17868 26641
rect 18084 26639 18086 26793
rect 18100 26785 18107 26793
rect 18108 26658 18110 26793
rect 18127 26785 18134 26833
rect 18136 26793 18138 26833
rect 18132 26658 18134 26785
rect 18158 26667 18162 26833
rect 18163 26793 18174 26833
rect 18176 26793 18183 26833
rect 18185 26793 18188 26833
rect 18190 26793 18201 26833
rect 18203 26793 18206 26833
rect 18096 26650 18110 26658
rect 18124 26650 18136 26658
rect 18156 26650 18164 26658
rect 18092 26642 18096 26650
rect 18108 26639 18110 26650
rect 18120 26642 18124 26650
rect 18132 26639 18134 26650
rect 18164 26642 18172 26650
rect 18180 26639 18182 26793
rect 18183 26785 18188 26793
rect 18212 26667 18216 26793
rect 18252 26658 18254 26979
rect 18256 26970 18257 26979
rect 18348 26969 18352 26979
rect 18257 26919 18264 26967
rect 18348 26956 18358 26969
rect 18346 26942 18350 26956
rect 18283 26667 18292 26843
rect 18348 26658 18350 26942
rect 18359 26942 18360 26956
rect 18367 26942 18374 26959
rect 18385 26955 18388 26965
rect 18396 26955 18398 26979
rect 18359 26932 18374 26942
rect 18395 26939 18398 26955
rect 18436 26948 18445 26979
rect 18492 26971 18494 26979
rect 18491 26961 18496 26971
rect 18512 26961 18518 26979
rect 18492 26957 18496 26961
rect 18359 26916 18375 26932
rect 18359 26911 18374 26916
rect 18359 26847 18368 26911
rect 18359 26837 18375 26847
rect 18376 26667 18385 26837
rect 18396 26658 18398 26939
rect 18422 26934 18424 26939
rect 18434 26934 18436 26939
rect 18436 26929 18444 26934
rect 18490 26931 18497 26957
rect 18446 26924 18454 26929
rect 18443 26883 18449 26909
rect 18468 26908 18470 26911
rect 18424 26819 18429 26847
rect 18472 26839 18477 26841
rect 18442 26829 18446 26837
rect 18425 26789 18429 26819
rect 18430 26789 18441 26829
rect 18443 26789 18446 26829
rect 18425 26781 18428 26789
rect 18452 26667 18456 26789
rect 18472 26667 18478 26839
rect 18492 26829 18494 26931
rect 18516 26901 18518 26961
rect 18554 26915 18557 26925
rect 18564 26917 18566 26979
rect 18577 26977 18582 26979
rect 18586 26953 18593 26979
rect 18516 26885 18524 26901
rect 18564 26893 18568 26917
rect 18516 26861 18525 26885
rect 18505 26841 18508 26851
rect 18516 26841 18518 26861
rect 18497 26839 18504 26841
rect 18497 26829 18505 26839
rect 18515 26829 18518 26841
rect 18479 26793 18488 26829
rect 18490 26793 18495 26829
rect 18499 26793 18505 26829
rect 18506 26793 18522 26829
rect 18490 26785 18497 26793
rect 18516 26785 18522 26793
rect 18492 26658 18494 26785
rect 18516 26658 18518 26785
rect 18526 26667 18532 26839
rect 18536 26833 18542 26841
rect 18548 26793 18554 26833
rect 18548 26667 18552 26793
rect 18184 26650 18192 26658
rect 18246 26650 18256 26658
rect 18274 26650 18284 26658
rect 18306 26650 18314 26658
rect 18334 26650 18350 26658
rect 18366 26650 18378 26658
rect 18394 26650 18406 26658
rect 18426 26650 18434 26658
rect 18454 26650 18468 26658
rect 18484 26650 18496 26658
rect 18512 26650 18524 26658
rect 18192 26642 18200 26650
rect 18240 26642 18246 26650
rect 18252 26639 18254 26650
rect 18268 26642 18274 26650
rect 18314 26642 18322 26650
rect 18348 26639 18350 26650
rect 18362 26642 18366 26650
rect 18390 26642 18394 26650
rect 18396 26639 18398 26650
rect 18434 26642 18442 26650
rect 18468 26642 18470 26650
rect 18482 26642 18484 26650
rect 18492 26639 18494 26650
rect 18496 26642 18498 26650
rect 18510 26642 18512 26650
rect 18516 26639 18518 26650
rect 18524 26642 18526 26650
rect 18564 26639 18566 26893
rect 18568 26667 18574 26841
rect 18588 26833 18590 26953
rect 18601 26841 18604 26851
rect 18612 26841 18614 26979
rect 18650 26915 18653 26925
rect 18660 26917 18662 26979
rect 18673 26977 18678 26979
rect 18682 26953 18689 26979
rect 18660 26893 18664 26917
rect 18593 26833 18601 26841
rect 18611 26833 18614 26841
rect 18575 26793 18584 26833
rect 18586 26793 18591 26833
rect 18595 26793 18601 26833
rect 18602 26793 18618 26833
rect 18586 26785 18593 26793
rect 18612 26785 18618 26793
rect 18588 26658 18590 26785
rect 18612 26658 18614 26785
rect 18622 26667 18628 26841
rect 18632 26833 18638 26841
rect 18644 26793 18650 26833
rect 18644 26667 18648 26793
rect 18580 26650 18590 26658
rect 18608 26650 18616 26658
rect 18572 26642 18580 26650
rect 18588 26639 18590 26650
rect 18600 26642 18608 26650
rect 18612 26639 18614 26650
rect 18660 26639 18662 26893
rect 18664 26667 18670 26841
rect 18684 26833 18686 26953
rect 18697 26841 18700 26851
rect 18708 26841 18710 26979
rect 18746 26915 18749 26925
rect 18756 26917 18758 26979
rect 18769 26977 18774 26979
rect 18778 26953 18785 26979
rect 18756 26893 18760 26917
rect 18689 26833 18697 26841
rect 18707 26833 18710 26841
rect 18671 26793 18680 26833
rect 18682 26793 18687 26833
rect 18691 26793 18697 26833
rect 18698 26793 18714 26833
rect 18682 26785 18689 26793
rect 18708 26785 18714 26793
rect 18684 26658 18686 26785
rect 18708 26658 18710 26785
rect 18718 26667 18724 26841
rect 18728 26833 18734 26841
rect 18740 26793 18746 26833
rect 18740 26667 18744 26793
rect 18676 26650 18686 26658
rect 18704 26650 18712 26658
rect 18668 26642 18676 26650
rect 18684 26639 18686 26650
rect 18696 26642 18704 26650
rect 18708 26639 18710 26650
rect 18756 26639 18758 26893
rect 18760 26667 18766 26841
rect 18780 26833 18782 26953
rect 18793 26841 18796 26851
rect 18804 26841 18806 26979
rect 18849 26917 18855 26979
rect 18868 26969 18871 26979
rect 18876 26969 18880 26979
rect 18876 26953 18879 26969
rect 18839 26907 18844 26913
rect 18839 26903 18846 26907
rect 18849 26893 18856 26917
rect 18849 26889 18854 26893
rect 18852 26841 18854 26889
rect 18868 26891 18871 26953
rect 18868 26889 18873 26891
rect 18868 26851 18871 26889
rect 18876 26851 18878 26953
rect 18865 26841 18878 26851
rect 18785 26833 18793 26841
rect 18803 26833 18806 26841
rect 18767 26793 18776 26833
rect 18778 26793 18783 26833
rect 18787 26793 18793 26833
rect 18794 26793 18810 26833
rect 18778 26785 18785 26793
rect 18804 26785 18810 26793
rect 18780 26658 18782 26785
rect 18804 26658 18806 26785
rect 18814 26667 18820 26841
rect 18824 26833 18830 26841
rect 18852 26833 18861 26841
rect 18869 26833 18878 26841
rect 18881 26841 18885 26979
rect 18895 26841 18898 26979
rect 18836 26793 18842 26833
rect 18850 26793 18861 26833
rect 18863 26793 18866 26833
rect 18868 26793 18879 26833
rect 18881 26793 18888 26841
rect 18900 26833 18902 26979
rect 18944 26978 18950 26979
rect 18937 26841 18940 26851
rect 18948 26841 18950 26978
rect 18996 26903 18998 26979
rect 19009 26977 19015 26979
rect 19018 26970 19025 26979
rect 19020 26903 19022 26970
rect 18996 26901 19027 26903
rect 18916 26833 18920 26841
rect 18944 26833 18950 26841
rect 18970 26833 18974 26841
rect 18890 26793 18893 26833
rect 18836 26667 18840 26793
rect 18772 26650 18782 26658
rect 18800 26650 18808 26658
rect 18832 26650 18848 26658
rect 18764 26642 18772 26650
rect 18780 26639 18782 26650
rect 18792 26642 18800 26650
rect 18804 26639 18806 26650
rect 18852 26639 18854 26793
rect 18868 26785 18875 26793
rect 18876 26658 18878 26793
rect 18895 26785 18902 26833
rect 18904 26793 18906 26833
rect 18900 26658 18902 26785
rect 18926 26667 18930 26833
rect 18931 26793 18942 26833
rect 18944 26793 18951 26833
rect 18953 26793 18956 26833
rect 18958 26793 18969 26833
rect 18971 26793 18974 26833
rect 18864 26650 18878 26658
rect 18892 26650 18904 26658
rect 18924 26650 18932 26658
rect 18860 26642 18864 26650
rect 18876 26639 18878 26650
rect 18888 26642 18892 26650
rect 18900 26639 18902 26650
rect 18932 26642 18940 26650
rect 18948 26639 18950 26793
rect 18951 26785 18956 26793
rect 18980 26667 18984 26793
rect 18996 26658 18998 26901
rect 19000 26667 19006 26841
rect 19020 26833 19022 26901
rect 19033 26841 19036 26851
rect 19044 26841 19046 26979
rect 19082 26915 19085 26925
rect 19092 26917 19094 26979
rect 19105 26977 19110 26979
rect 19114 26953 19121 26979
rect 19092 26893 19096 26917
rect 19025 26833 19033 26841
rect 19043 26833 19046 26841
rect 19007 26793 19016 26833
rect 19018 26793 19023 26833
rect 19027 26793 19033 26833
rect 19034 26793 19050 26833
rect 19018 26785 19025 26793
rect 19044 26785 19050 26793
rect 19020 26658 19022 26785
rect 19044 26658 19046 26785
rect 19054 26667 19060 26841
rect 19064 26833 19070 26841
rect 19076 26793 19082 26833
rect 19076 26667 19080 26793
rect 18952 26650 18960 26658
rect 18980 26650 18998 26658
rect 19012 26650 19024 26658
rect 19040 26650 19052 26658
rect 18960 26642 18968 26650
rect 18996 26639 18998 26650
rect 19008 26642 19012 26650
rect 19020 26639 19022 26650
rect 19036 26642 19040 26650
rect 19044 26639 19046 26650
rect 19092 26639 19094 26893
rect 19096 26667 19102 26841
rect 19116 26833 19118 26953
rect 19129 26841 19132 26851
rect 19140 26841 19142 26979
rect 19188 26917 19190 26979
rect 19191 26953 19207 26964
rect 19191 26917 19197 26953
rect 19188 26916 19197 26917
rect 19217 26916 19219 26964
rect 19188 26893 19192 26916
rect 19121 26833 19129 26841
rect 19139 26833 19142 26841
rect 19103 26793 19112 26833
rect 19114 26793 19119 26833
rect 19123 26793 19129 26833
rect 19130 26793 19146 26833
rect 19114 26785 19121 26793
rect 19140 26785 19146 26793
rect 19116 26658 19118 26785
rect 19140 26658 19142 26785
rect 19150 26667 19156 26841
rect 19160 26833 19166 26841
rect 19172 26793 19178 26833
rect 19172 26667 19176 26793
rect 19108 26650 19118 26658
rect 19136 26650 19144 26658
rect 19100 26642 19108 26650
rect 19116 26639 19118 26650
rect 19128 26642 19136 26650
rect 19140 26639 19142 26650
rect 19188 26639 19190 26893
rect 19236 26658 19238 26979
rect 19267 26916 19279 26956
rect 19332 26658 19334 26979
rect 19425 26969 19432 26979
rect 19336 26919 19352 26956
rect 19354 26911 19355 26956
rect 19363 26667 19365 26966
rect 19425 26959 19435 26969
rect 19444 26959 19447 26979
rect 19415 26903 19420 26913
rect 19428 26903 19430 26959
rect 19439 26911 19451 26959
rect 19439 26903 19447 26911
rect 19425 26889 19430 26903
rect 19202 26650 19212 26658
rect 19230 26650 19240 26658
rect 19262 26650 19270 26658
rect 19326 26650 19334 26658
rect 19354 26650 19362 26658
rect 19386 26650 19394 26658
rect 19414 26650 19424 26658
rect 19428 26650 19430 26889
rect 19476 26658 19478 26979
rect 19520 26978 19526 26979
rect 19513 26841 19516 26851
rect 19524 26841 19526 26978
rect 19572 26903 19574 26979
rect 19585 26977 19591 26979
rect 19594 26970 19601 26979
rect 19596 26903 19598 26970
rect 19572 26901 19603 26903
rect 19492 26833 19496 26841
rect 19520 26833 19526 26841
rect 19546 26833 19550 26841
rect 19502 26667 19506 26833
rect 19507 26793 19518 26833
rect 19520 26793 19527 26833
rect 19529 26793 19532 26833
rect 19534 26793 19545 26833
rect 19547 26793 19550 26833
rect 19442 26650 19452 26658
rect 19470 26650 19480 26658
rect 19500 26650 19508 26658
rect 19196 26642 19202 26650
rect 19224 26642 19230 26650
rect 19236 26639 19238 26650
rect 19270 26642 19278 26650
rect 19318 26642 19326 26650
rect 19332 26639 19334 26650
rect 19346 26642 19354 26650
rect 19394 26642 19402 26650
rect 19424 26642 19430 26650
rect 19452 26642 19458 26650
rect 19428 26639 19430 26642
rect 19476 26639 19478 26650
rect 19480 26642 19486 26650
rect 19508 26642 19516 26650
rect 19524 26639 19526 26793
rect 19527 26785 19532 26793
rect 19556 26667 19560 26793
rect 19572 26658 19574 26901
rect 19576 26667 19582 26841
rect 19596 26833 19598 26901
rect 19609 26841 19612 26851
rect 19620 26841 19622 26979
rect 19665 26917 19671 26979
rect 19684 26969 19687 26979
rect 19692 26969 19696 26979
rect 19692 26953 19695 26969
rect 19655 26907 19660 26913
rect 19655 26903 19662 26907
rect 19665 26893 19672 26917
rect 19665 26889 19670 26893
rect 19668 26841 19670 26889
rect 19684 26891 19687 26953
rect 19684 26889 19689 26891
rect 19684 26851 19687 26889
rect 19692 26851 19694 26953
rect 19681 26841 19694 26851
rect 19601 26833 19609 26841
rect 19619 26833 19622 26841
rect 19583 26793 19592 26833
rect 19594 26793 19599 26833
rect 19603 26793 19609 26833
rect 19610 26793 19626 26833
rect 19594 26785 19601 26793
rect 19620 26785 19626 26793
rect 19596 26658 19598 26785
rect 19620 26658 19622 26785
rect 19630 26667 19636 26841
rect 19640 26833 19646 26841
rect 19668 26833 19677 26841
rect 19685 26833 19694 26841
rect 19697 26841 19701 26979
rect 19711 26841 19714 26979
rect 19652 26793 19658 26833
rect 19666 26793 19677 26833
rect 19679 26793 19682 26833
rect 19684 26793 19695 26833
rect 19697 26793 19704 26841
rect 19716 26833 19718 26979
rect 19760 26978 19766 26979
rect 19753 26841 19756 26851
rect 19764 26841 19766 26978
rect 19799 26903 19804 26913
rect 19812 26903 19814 26979
rect 19832 26972 19841 26979
rect 19809 26889 19814 26903
rect 19812 26843 19814 26889
rect 19732 26833 19736 26841
rect 19760 26833 19766 26841
rect 19786 26833 19790 26841
rect 19706 26793 19709 26833
rect 19652 26667 19656 26793
rect 19528 26650 19536 26658
rect 19556 26650 19574 26658
rect 19588 26650 19600 26658
rect 19616 26650 19628 26658
rect 19648 26650 19664 26658
rect 19536 26642 19544 26650
rect 19572 26639 19574 26650
rect 19584 26642 19588 26650
rect 19596 26639 19598 26650
rect 19612 26642 19616 26650
rect 19620 26639 19622 26650
rect 19668 26639 19670 26793
rect 19684 26785 19691 26793
rect 19692 26658 19694 26793
rect 19711 26785 19718 26833
rect 19720 26793 19722 26833
rect 19716 26658 19718 26785
rect 19742 26667 19746 26833
rect 19747 26793 19758 26833
rect 19760 26793 19767 26833
rect 19769 26793 19772 26833
rect 19774 26793 19785 26833
rect 19787 26793 19790 26833
rect 19680 26650 19694 26658
rect 19708 26650 19720 26658
rect 19740 26650 19748 26658
rect 19676 26642 19680 26650
rect 19692 26639 19694 26650
rect 19704 26642 19708 26650
rect 19716 26639 19718 26650
rect 19748 26642 19756 26650
rect 19764 26639 19766 26793
rect 19767 26785 19772 26793
rect 19796 26667 19800 26793
rect 19812 26791 19822 26843
rect 19830 26839 19833 26849
rect 19836 26833 19838 26972
rect 19841 26839 19848 26972
rect 19849 26953 19852 26963
rect 19860 26953 19862 26979
rect 19859 26937 19862 26953
rect 19823 26791 19829 26833
rect 19768 26650 19776 26658
rect 19796 26650 19810 26658
rect 19812 26650 19814 26791
rect 19831 26785 19838 26833
rect 19840 26785 19849 26839
rect 19860 26833 19862 26937
rect 19875 26895 19877 26899
rect 19885 26881 19887 26895
rect 19850 26791 19856 26833
rect 19858 26785 19865 26833
rect 19867 26791 19876 26843
rect 19889 26791 19893 26849
rect 19906 26831 19910 26839
rect 19894 26791 19905 26831
rect 19907 26791 19910 26831
rect 19836 26658 19838 26785
rect 19841 26783 19848 26785
rect 19860 26658 19862 26785
rect 19889 26783 19892 26791
rect 19916 26667 19920 26791
rect 19826 26650 19838 26658
rect 19854 26650 19866 26658
rect 19886 26650 19894 26658
rect 19776 26642 19784 26650
rect 19810 26642 19814 26650
rect 19824 26642 19826 26650
rect 19836 26642 19840 26650
rect 19852 26642 19854 26650
rect 19812 26639 19814 26642
rect 19836 26639 19838 26642
rect 19860 26639 19862 26650
rect 19866 26642 19868 26650
rect 19894 26642 19902 26650
rect 19932 26639 19934 26979
rect 19956 26977 19970 26979
rect 19956 26969 19958 26977
rect 19955 26961 19960 26969
rect 19956 26955 19960 26961
rect 19954 26929 19961 26955
rect 19936 26667 19942 26841
rect 19956 26831 19958 26929
rect 19969 26841 19972 26851
rect 19980 26841 19982 26979
rect 20028 26917 20031 26979
rect 20048 26972 20057 26979
rect 20052 26969 20056 26972
rect 20052 26953 20055 26969
rect 20015 26907 20020 26913
rect 20015 26903 20022 26907
rect 20028 26903 20032 26917
rect 20025 26893 20032 26903
rect 20025 26889 20030 26893
rect 20028 26843 20030 26889
rect 20045 26849 20049 26889
rect 20052 26849 20054 26953
rect 19961 26831 19969 26841
rect 19979 26831 19982 26841
rect 19943 26793 19952 26831
rect 19954 26793 19959 26831
rect 19963 26793 19969 26831
rect 19970 26793 19986 26831
rect 19954 26785 19961 26793
rect 19980 26785 19986 26793
rect 19956 26658 19958 26785
rect 19980 26658 19982 26785
rect 19990 26667 19996 26841
rect 20000 26833 20006 26841
rect 20012 26793 20018 26833
rect 20012 26667 20016 26793
rect 20028 26791 20038 26843
rect 20045 26839 20055 26849
rect 20057 26839 20064 26972
rect 20065 26953 20068 26963
rect 20076 26953 20078 26979
rect 20075 26937 20078 26953
rect 20052 26833 20054 26839
rect 20039 26791 20045 26833
rect 19948 26650 19958 26658
rect 19976 26650 19986 26658
rect 19942 26642 19948 26650
rect 19956 26639 19958 26650
rect 19970 26642 19976 26650
rect 19980 26639 19982 26650
rect 20028 26639 20030 26791
rect 20047 26785 20054 26833
rect 20056 26785 20065 26839
rect 20076 26833 20078 26937
rect 20091 26895 20093 26899
rect 20101 26881 20103 26895
rect 20066 26791 20072 26833
rect 20074 26785 20081 26833
rect 20083 26791 20092 26843
rect 20105 26791 20109 26849
rect 20122 26831 20126 26839
rect 20110 26791 20121 26831
rect 20123 26791 20126 26831
rect 20052 26658 20054 26785
rect 20057 26783 20064 26785
rect 20076 26658 20078 26785
rect 20105 26783 20108 26791
rect 20132 26667 20136 26791
rect 20042 26650 20054 26658
rect 20070 26650 20080 26658
rect 20102 26650 20110 26658
rect 20036 26642 20042 26650
rect 20052 26639 20054 26650
rect 20064 26642 20070 26650
rect 20076 26639 20078 26650
rect 20110 26642 20118 26650
rect 20148 26639 20150 26979
rect 20172 26977 20186 26979
rect 20172 26969 20174 26977
rect 20171 26961 20176 26969
rect 20172 26955 20176 26961
rect 20170 26929 20177 26955
rect 20152 26667 20158 26841
rect 20172 26831 20174 26929
rect 20185 26841 20188 26851
rect 20196 26841 20198 26979
rect 20234 26915 20237 26925
rect 20244 26917 20246 26979
rect 20257 26977 20262 26979
rect 20266 26953 20273 26979
rect 20244 26893 20248 26917
rect 20177 26831 20185 26841
rect 20195 26831 20198 26841
rect 20159 26793 20168 26831
rect 20170 26793 20175 26831
rect 20179 26793 20185 26831
rect 20186 26793 20202 26831
rect 20170 26785 20177 26793
rect 20196 26785 20202 26793
rect 20172 26658 20174 26785
rect 20196 26658 20198 26785
rect 20206 26667 20212 26841
rect 20216 26833 20222 26841
rect 20228 26793 20234 26833
rect 20228 26667 20232 26793
rect 20164 26650 20174 26658
rect 20192 26650 20202 26658
rect 20158 26642 20164 26650
rect 20172 26639 20174 26650
rect 20186 26642 20192 26650
rect 20196 26639 20198 26650
rect 20244 26639 20246 26893
rect 20248 26667 20254 26841
rect 20268 26833 20270 26953
rect 20281 26841 20284 26851
rect 20292 26841 20294 26979
rect 20340 26917 20342 26979
rect 20343 26953 20359 26964
rect 20343 26917 20349 26953
rect 20340 26916 20349 26917
rect 20369 26916 20371 26964
rect 20340 26893 20344 26916
rect 20273 26833 20281 26841
rect 20291 26833 20294 26841
rect 20255 26793 20264 26833
rect 20266 26793 20271 26833
rect 20275 26793 20281 26833
rect 20282 26793 20298 26833
rect 20266 26785 20273 26793
rect 20292 26785 20298 26793
rect 20268 26658 20270 26785
rect 20292 26658 20294 26785
rect 20302 26667 20308 26841
rect 20312 26833 20318 26841
rect 20324 26793 20330 26833
rect 20324 26667 20328 26793
rect 20260 26650 20270 26658
rect 20288 26650 20296 26658
rect 20252 26642 20260 26650
rect 20268 26639 20270 26650
rect 20280 26642 20288 26650
rect 20292 26639 20294 26650
rect 20340 26639 20342 26893
rect 20388 26658 20390 26979
rect 20482 26977 20489 26979
rect 20482 26966 20491 26977
rect 20482 26961 20499 26966
rect 20419 26916 20431 26956
rect 20482 26900 20489 26961
rect 20504 26908 20507 26956
rect 20484 26851 20486 26900
rect 20483 26667 20490 26851
rect 20497 26841 20500 26851
rect 20508 26841 20510 26979
rect 20556 26917 20559 26979
rect 20576 26972 20585 26979
rect 20580 26969 20584 26972
rect 20580 26953 20583 26969
rect 20543 26907 20548 26913
rect 20543 26903 20550 26907
rect 20556 26903 20560 26917
rect 20553 26893 20560 26903
rect 20553 26889 20558 26893
rect 20556 26843 20558 26889
rect 20573 26849 20577 26889
rect 20580 26849 20582 26953
rect 20507 26793 20510 26841
rect 20528 26833 20534 26841
rect 20484 26658 20486 26667
rect 20508 26658 20510 26793
rect 20540 26793 20546 26833
rect 20540 26667 20544 26793
rect 20556 26791 20566 26843
rect 20573 26839 20583 26849
rect 20585 26839 20592 26972
rect 20593 26953 20596 26963
rect 20604 26953 20606 26979
rect 20603 26937 20606 26953
rect 20580 26833 20582 26839
rect 20567 26791 20573 26833
rect 20354 26650 20364 26658
rect 20382 26650 20392 26658
rect 20414 26650 20422 26658
rect 20476 26650 20486 26658
rect 20504 26650 20514 26658
rect 20348 26642 20354 26650
rect 20376 26642 20382 26650
rect 20388 26639 20390 26650
rect 20422 26642 20430 26650
rect 20470 26642 20476 26650
rect 20484 26639 20486 26650
rect 20498 26642 20504 26650
rect 20508 26639 20510 26650
rect 20556 26639 20558 26791
rect 20575 26785 20582 26833
rect 20584 26785 20593 26839
rect 20604 26833 20606 26937
rect 20700 26969 20702 26979
rect 20913 26969 20920 26979
rect 20700 26955 20704 26969
rect 20824 26967 20833 26969
rect 20705 26955 20712 26967
rect 20700 26945 20712 26955
rect 20619 26895 20621 26899
rect 20629 26881 20631 26895
rect 20594 26791 20600 26833
rect 20602 26785 20609 26833
rect 20611 26791 20620 26843
rect 20633 26791 20637 26849
rect 20650 26831 20654 26839
rect 20638 26791 20649 26831
rect 20651 26791 20654 26831
rect 20580 26658 20582 26785
rect 20585 26783 20592 26785
rect 20604 26658 20606 26785
rect 20633 26783 20636 26791
rect 20660 26667 20664 26791
rect 20700 26658 20702 26945
rect 20704 26929 20712 26945
rect 20705 26919 20712 26929
rect 20824 26919 20835 26967
rect 20913 26959 20923 26969
rect 20932 26959 20935 26979
rect 20903 26903 20908 26913
rect 20916 26903 20918 26959
rect 20927 26911 20939 26959
rect 20927 26903 20935 26911
rect 20913 26889 20918 26903
rect 20731 26667 20740 26841
rect 20570 26650 20582 26658
rect 20598 26650 20608 26658
rect 20630 26650 20638 26658
rect 20694 26650 20702 26658
rect 20722 26650 20730 26658
rect 20754 26650 20762 26658
rect 20782 26650 20798 26658
rect 20814 26650 20826 26658
rect 20842 26650 20854 26658
rect 20874 26650 20882 26658
rect 20902 26650 20912 26658
rect 20916 26650 20918 26889
rect 20964 26658 20966 26979
rect 21008 26978 21014 26979
rect 21001 26841 21004 26851
rect 21012 26841 21014 26978
rect 21060 26903 21062 26979
rect 21073 26977 21079 26979
rect 21082 26970 21089 26979
rect 21084 26903 21086 26970
rect 21060 26901 21091 26903
rect 20980 26833 20984 26841
rect 21008 26833 21014 26841
rect 21034 26833 21038 26841
rect 20990 26667 20994 26833
rect 20995 26793 21006 26833
rect 21008 26793 21015 26833
rect 21017 26793 21020 26833
rect 21022 26793 21033 26833
rect 21035 26793 21038 26833
rect 20930 26650 20940 26658
rect 20958 26650 20968 26658
rect 20988 26650 20996 26658
rect 20564 26642 20570 26650
rect 20580 26639 20582 26650
rect 20592 26642 20598 26650
rect 20604 26639 20606 26650
rect 20638 26642 20646 26650
rect 20686 26642 20694 26650
rect 20700 26639 20702 26650
rect 20714 26642 20722 26650
rect 20762 26642 20770 26650
rect 20810 26642 20814 26650
rect 20838 26642 20842 26650
rect 20882 26642 20890 26650
rect 20912 26642 20918 26650
rect 20940 26642 20946 26650
rect 20916 26639 20918 26642
rect 20964 26639 20966 26650
rect 20968 26642 20974 26650
rect 20996 26642 21004 26650
rect 21012 26639 21014 26793
rect 21015 26785 21020 26793
rect 21044 26667 21048 26793
rect 21060 26658 21062 26901
rect 21064 26667 21070 26841
rect 21084 26833 21086 26901
rect 21097 26841 21100 26851
rect 21108 26841 21110 26979
rect 21156 26917 21158 26979
rect 21159 26953 21175 26964
rect 21159 26917 21165 26953
rect 21156 26916 21165 26917
rect 21185 26916 21187 26964
rect 21156 26893 21160 26916
rect 21089 26833 21097 26841
rect 21107 26833 21110 26841
rect 21071 26793 21080 26833
rect 21082 26793 21087 26833
rect 21091 26793 21097 26833
rect 21098 26793 21114 26833
rect 21082 26785 21089 26793
rect 21108 26785 21114 26793
rect 21084 26658 21086 26785
rect 21108 26658 21110 26785
rect 21118 26667 21124 26841
rect 21128 26833 21134 26841
rect 21140 26793 21146 26833
rect 21140 26667 21144 26793
rect 21016 26650 21024 26658
rect 21044 26650 21062 26658
rect 21076 26650 21088 26658
rect 21104 26650 21116 26658
rect 21024 26642 21032 26650
rect 21060 26639 21062 26650
rect 21072 26642 21076 26650
rect 21084 26639 21086 26650
rect 21100 26642 21104 26650
rect 21108 26639 21110 26650
rect 21156 26639 21158 26893
rect 21204 26658 21206 26979
rect 21235 26916 21247 26956
rect 21297 26908 21299 26956
rect 21300 26851 21302 26979
rect 21319 26908 21323 26956
rect 21289 26841 21292 26851
rect 21299 26667 21302 26851
rect 21318 26841 21323 26851
rect 21300 26658 21302 26667
rect 21324 26658 21326 26979
rect 21368 26978 21374 26979
rect 21361 26841 21364 26851
rect 21372 26841 21374 26978
rect 21420 26903 21422 26979
rect 21433 26977 21439 26979
rect 21442 26970 21449 26979
rect 21444 26903 21446 26970
rect 21420 26901 21451 26903
rect 21328 26667 21333 26841
rect 21340 26833 21344 26841
rect 21368 26833 21374 26841
rect 21394 26833 21398 26841
rect 21350 26667 21354 26833
rect 21355 26793 21366 26833
rect 21368 26793 21375 26833
rect 21377 26793 21380 26833
rect 21382 26793 21393 26833
rect 21395 26793 21398 26833
rect 21170 26650 21180 26658
rect 21198 26650 21208 26658
rect 21230 26650 21238 26658
rect 21258 26650 21272 26658
rect 21288 26650 21302 26658
rect 21316 26650 21328 26658
rect 21348 26650 21356 26658
rect 21164 26642 21170 26650
rect 21192 26642 21198 26650
rect 21204 26639 21206 26650
rect 21238 26642 21246 26650
rect 21272 26642 21274 26650
rect 21286 26642 21288 26650
rect 21300 26639 21302 26650
rect 21314 26642 21316 26650
rect 21324 26639 21326 26650
rect 21328 26642 21330 26650
rect 21356 26642 21364 26650
rect 21372 26639 21374 26793
rect 21375 26785 21380 26793
rect 21404 26667 21408 26793
rect 21420 26658 21422 26901
rect 21424 26667 21430 26841
rect 21444 26833 21446 26901
rect 21457 26841 21460 26851
rect 21468 26841 21470 26979
rect 21513 26917 21519 26979
rect 21532 26969 21535 26979
rect 21540 26969 21544 26979
rect 21540 26953 21543 26969
rect 21503 26907 21508 26913
rect 21503 26903 21510 26907
rect 21513 26893 21520 26917
rect 21513 26889 21518 26893
rect 21516 26841 21518 26889
rect 21532 26891 21535 26953
rect 21532 26889 21537 26891
rect 21532 26851 21535 26889
rect 21540 26851 21542 26953
rect 21529 26841 21542 26851
rect 21449 26833 21457 26841
rect 21467 26833 21470 26841
rect 21431 26793 21440 26833
rect 21442 26793 21447 26833
rect 21451 26793 21457 26833
rect 21458 26793 21474 26833
rect 21442 26785 21449 26793
rect 21468 26785 21474 26793
rect 21444 26658 21446 26785
rect 21468 26658 21470 26785
rect 21478 26667 21484 26841
rect 21488 26833 21494 26841
rect 21516 26833 21525 26841
rect 21533 26833 21542 26841
rect 21545 26841 21549 26979
rect 21559 26841 21562 26979
rect 21500 26793 21506 26833
rect 21514 26793 21525 26833
rect 21527 26793 21530 26833
rect 21532 26793 21543 26833
rect 21545 26793 21552 26841
rect 21564 26833 21566 26979
rect 21608 26978 21614 26979
rect 21601 26841 21604 26851
rect 21612 26841 21614 26978
rect 21647 26903 21652 26913
rect 21660 26903 21662 26979
rect 21680 26972 21689 26979
rect 21657 26889 21662 26903
rect 21660 26843 21662 26889
rect 21580 26833 21584 26841
rect 21608 26833 21614 26841
rect 21634 26833 21638 26841
rect 21554 26793 21557 26833
rect 21500 26667 21504 26793
rect 21376 26650 21384 26658
rect 21404 26650 21422 26658
rect 21436 26650 21448 26658
rect 21464 26650 21476 26658
rect 21496 26650 21512 26658
rect 21384 26642 21392 26650
rect 21420 26639 21422 26650
rect 21432 26642 21436 26650
rect 21444 26639 21446 26650
rect 21460 26642 21464 26650
rect 21468 26639 21470 26650
rect 21516 26639 21518 26793
rect 21532 26785 21539 26793
rect 21540 26658 21542 26793
rect 21559 26785 21566 26833
rect 21568 26793 21570 26833
rect 21564 26658 21566 26785
rect 21590 26667 21594 26833
rect 21595 26793 21606 26833
rect 21608 26793 21615 26833
rect 21617 26793 21620 26833
rect 21622 26793 21633 26833
rect 21635 26793 21638 26833
rect 21528 26650 21542 26658
rect 21556 26650 21568 26658
rect 21588 26650 21596 26658
rect 21524 26642 21528 26650
rect 21540 26639 21542 26650
rect 21552 26642 21556 26650
rect 21564 26639 21566 26650
rect 21596 26642 21604 26650
rect 21612 26639 21614 26793
rect 21615 26785 21620 26793
rect 21644 26667 21648 26793
rect 21660 26791 21670 26843
rect 21678 26839 21681 26849
rect 21684 26833 21686 26972
rect 21689 26839 21696 26972
rect 21697 26953 21700 26963
rect 21708 26953 21710 26979
rect 21707 26937 21710 26953
rect 21671 26791 21677 26833
rect 21616 26650 21624 26658
rect 21644 26650 21658 26658
rect 21660 26650 21662 26791
rect 21679 26785 21686 26833
rect 21688 26785 21697 26839
rect 21708 26833 21710 26937
rect 21767 26903 21772 26913
rect 21780 26903 21782 26979
rect 21803 26977 21816 26979
rect 21803 26972 21806 26977
rect 21723 26895 21725 26899
rect 21733 26881 21735 26895
rect 21777 26889 21782 26903
rect 21698 26791 21704 26833
rect 21706 26785 21713 26833
rect 21715 26791 21724 26843
rect 21737 26791 21741 26849
rect 21780 26841 21782 26889
rect 21804 26969 21806 26972
rect 21804 26945 21808 26969
rect 21754 26831 21758 26839
rect 21742 26791 21753 26831
rect 21755 26791 21758 26831
rect 21780 26791 21790 26841
rect 21798 26839 21801 26849
rect 21804 26831 21806 26945
rect 21809 26839 21816 26972
rect 21817 26953 21820 26963
rect 21828 26953 21830 26979
rect 21827 26937 21830 26953
rect 21791 26791 21797 26831
rect 21684 26658 21686 26785
rect 21689 26783 21696 26785
rect 21708 26658 21710 26785
rect 21737 26783 21740 26791
rect 21764 26667 21768 26791
rect 21674 26650 21686 26658
rect 21702 26650 21714 26658
rect 21734 26650 21742 26658
rect 21762 26650 21778 26658
rect 21624 26642 21632 26650
rect 21658 26642 21662 26650
rect 21672 26642 21674 26650
rect 21684 26642 21688 26650
rect 21700 26642 21702 26650
rect 21660 26639 21662 26642
rect 21684 26639 21686 26642
rect 21708 26639 21710 26650
rect 21714 26642 21716 26650
rect 21742 26642 21750 26650
rect 21780 26639 21782 26791
rect 21799 26783 21806 26831
rect 21808 26783 21817 26839
rect 21828 26831 21830 26937
rect 21887 26903 21892 26913
rect 21900 26903 21902 26979
rect 21923 26977 21936 26979
rect 21923 26972 21926 26977
rect 21843 26895 21845 26899
rect 21853 26881 21855 26895
rect 21897 26889 21902 26903
rect 21818 26791 21824 26831
rect 21826 26783 21833 26831
rect 21835 26791 21844 26841
rect 21857 26791 21861 26849
rect 21900 26841 21902 26889
rect 21924 26969 21926 26972
rect 21924 26945 21928 26969
rect 21874 26831 21878 26839
rect 21862 26791 21873 26831
rect 21875 26791 21878 26831
rect 21900 26791 21910 26841
rect 21918 26839 21921 26849
rect 21924 26831 21926 26945
rect 21929 26839 21936 26972
rect 21937 26953 21940 26963
rect 21948 26953 21950 26979
rect 22017 26964 22022 26979
rect 21947 26937 21950 26953
rect 21911 26791 21917 26831
rect 21857 26783 21860 26791
rect 21804 26658 21806 26783
rect 21828 26658 21830 26783
rect 21884 26667 21888 26791
rect 21794 26650 21806 26658
rect 21822 26650 21834 26658
rect 21854 26650 21862 26658
rect 21882 26650 21898 26658
rect 21790 26642 21794 26650
rect 21804 26639 21806 26650
rect 21818 26642 21822 26650
rect 21828 26639 21830 26650
rect 21862 26642 21870 26650
rect 21900 26639 21902 26791
rect 21919 26783 21926 26831
rect 21928 26783 21937 26839
rect 21948 26831 21950 26937
rect 22007 26903 22012 26913
rect 22020 26903 22022 26964
rect 22036 26945 22039 26979
rect 22044 26969 22046 26979
rect 22044 26945 22048 26969
rect 21963 26895 21965 26899
rect 21973 26881 21975 26895
rect 22017 26889 22022 26903
rect 21938 26791 21944 26831
rect 21946 26783 21953 26831
rect 21955 26791 21964 26841
rect 21977 26791 21981 26849
rect 22020 26841 22022 26889
rect 22036 26851 22039 26929
rect 22033 26841 22039 26851
rect 22044 26891 22046 26945
rect 22049 26891 22053 26979
rect 22044 26841 22053 26891
rect 22063 26841 22066 26979
rect 21994 26831 21998 26839
rect 22020 26831 22029 26841
rect 22043 26831 22056 26841
rect 22068 26831 22070 26979
rect 22112 26978 22118 26979
rect 22105 26841 22108 26851
rect 22116 26841 22118 26978
rect 22151 26903 22156 26913
rect 22164 26903 22166 26979
rect 22184 26972 22193 26979
rect 22161 26889 22166 26903
rect 22164 26843 22166 26889
rect 22084 26833 22088 26841
rect 22112 26833 22118 26841
rect 22138 26833 22142 26841
rect 21982 26791 21993 26831
rect 21995 26791 21998 26831
rect 22018 26793 22029 26831
rect 22031 26793 22034 26831
rect 22036 26793 22047 26831
rect 22049 26793 22056 26831
rect 22058 26793 22061 26831
rect 21977 26783 21980 26791
rect 21924 26658 21926 26783
rect 21948 26658 21950 26783
rect 22004 26667 22008 26791
rect 21914 26650 21926 26658
rect 21942 26650 21954 26658
rect 21974 26650 21982 26658
rect 22002 26650 22016 26658
rect 21910 26642 21914 26650
rect 21924 26639 21926 26650
rect 21938 26642 21942 26650
rect 21948 26639 21950 26650
rect 21982 26642 21990 26650
rect 22016 26642 22018 26650
rect 22020 26639 22022 26793
rect 22036 26785 22043 26793
rect 22044 26658 22046 26793
rect 22063 26785 22070 26831
rect 22072 26793 22074 26831
rect 22068 26658 22070 26785
rect 22094 26667 22098 26833
rect 22099 26793 22110 26833
rect 22112 26793 22119 26833
rect 22121 26793 22124 26833
rect 22126 26793 22137 26833
rect 22139 26793 22142 26833
rect 22032 26650 22046 26658
rect 22060 26650 22072 26658
rect 22092 26650 22100 26658
rect 22030 26642 22032 26650
rect 22044 26639 22046 26650
rect 22058 26642 22060 26650
rect 22068 26639 22070 26650
rect 22072 26642 22074 26650
rect 22100 26642 22108 26650
rect 22116 26639 22118 26793
rect 22119 26785 22124 26793
rect 22148 26667 22152 26793
rect 22164 26791 22174 26843
rect 22182 26839 22185 26849
rect 22188 26833 22190 26972
rect 22193 26839 22200 26972
rect 22201 26953 22204 26963
rect 22212 26953 22214 26979
rect 22321 26977 22324 26979
rect 22211 26937 22214 26953
rect 22175 26791 22181 26833
rect 22120 26650 22128 26658
rect 22148 26650 22162 26658
rect 22164 26650 22166 26791
rect 22183 26785 22190 26833
rect 22192 26785 22201 26839
rect 22212 26833 22214 26937
rect 22227 26895 22229 26899
rect 22237 26881 22239 26895
rect 22394 26882 22401 26979
rect 22444 26976 22447 26979
rect 22520 26968 22523 26979
rect 22561 26970 22564 26979
rect 22579 26978 22665 26979
rect 22614 26960 22617 26961
rect 22424 26952 22430 26960
rect 22437 26952 22451 26960
rect 22511 26952 22520 26953
rect 22580 26952 22582 26960
rect 22589 26952 22623 26960
rect 22444 26950 22447 26952
rect 22520 26950 22523 26952
rect 22430 26902 22437 26950
rect 22440 26902 22441 26942
rect 22425 26894 22434 26902
rect 22444 26894 22451 26942
rect 22462 26902 22469 26950
rect 22513 26947 22527 26950
rect 22520 26942 22527 26947
rect 22501 26902 22504 26942
rect 22456 26894 22501 26902
rect 22506 26894 22513 26942
rect 22521 26894 22527 26942
rect 22578 26902 22580 26942
rect 22582 26902 22589 26950
rect 22609 26947 22630 26950
rect 22623 26942 22630 26947
rect 22676 26942 22680 26978
rect 22597 26902 22598 26942
rect 22547 26894 22554 26902
rect 22600 26894 22607 26942
rect 22611 26902 22615 26942
rect 22623 26902 22627 26942
rect 22654 26902 22655 26942
rect 22630 26894 22637 26902
rect 22663 26894 22670 26942
rect 22444 26882 22447 26894
rect 22520 26892 22527 26894
rect 22520 26882 22523 26892
rect 22384 26874 22456 26882
rect 22501 26874 22578 26882
rect 22394 26872 22401 26874
rect 22404 26856 22408 26862
rect 22202 26791 22208 26833
rect 22210 26785 22217 26833
rect 22219 26791 22228 26843
rect 22241 26791 22245 26849
rect 22258 26831 22262 26839
rect 22246 26791 22257 26831
rect 22259 26791 22262 26831
rect 22188 26658 22190 26785
rect 22193 26783 22200 26785
rect 22212 26658 22214 26785
rect 22241 26783 22244 26791
rect 22268 26667 22272 26791
rect 22292 26667 22294 26841
rect 22320 26824 22325 26831
rect 22295 26783 22308 26824
rect 22318 26783 22320 26824
rect 22322 26783 22325 26824
rect 22328 26783 22338 26824
rect 22394 26816 22401 26856
rect 22444 26841 22447 26874
rect 22448 26864 22451 26874
rect 22458 26854 22461 26864
rect 22458 26848 22474 26854
rect 22502 26848 22514 26854
rect 22416 26824 22420 26834
rect 22430 26826 22452 26834
rect 22430 26825 22446 26826
rect 22520 26824 22523 26874
rect 22546 26854 22668 26859
rect 22572 26839 22590 26846
rect 22527 26826 22547 26834
rect 22676 26826 22680 26894
rect 22426 26820 22444 26824
rect 22313 26776 22318 26783
rect 22386 26768 22393 26816
rect 22426 26776 22432 26820
rect 22462 26776 22469 26824
rect 22520 26816 22528 26824
rect 22582 26816 22589 26824
rect 22502 26776 22504 26816
rect 22404 26768 22420 26775
rect 22426 26768 22430 26776
rect 22506 26768 22513 26816
rect 22521 26768 22528 26816
rect 22564 26777 22572 26816
rect 22564 26776 22580 26777
rect 22394 26705 22401 26768
rect 22520 26765 22528 26768
rect 22547 26765 22554 26776
rect 22572 26768 22580 26776
rect 22600 26768 22607 26816
rect 22609 26776 22613 26816
rect 22623 26776 22625 26824
rect 22630 26768 22637 26816
rect 22642 26778 22648 26816
rect 22676 26778 22683 26826
rect 22685 26778 22689 26816
rect 22663 26768 22670 26778
rect 22746 26771 22750 26818
rect 22819 26815 22822 26841
rect 22830 26815 22836 26979
rect 22860 26824 22867 26979
rect 22936 26841 22941 26979
rect 22951 26841 22953 26979
rect 23000 26978 23006 26979
rect 22993 26841 22996 26851
rect 23004 26841 23006 26978
rect 23039 26903 23044 26913
rect 23052 26903 23054 26979
rect 23049 26889 23054 26903
rect 23052 26841 23054 26889
rect 23068 26851 23071 26970
rect 23065 26841 23071 26851
rect 23076 26891 23078 26979
rect 23081 26891 23085 26979
rect 23076 26841 23085 26891
rect 23095 26841 23098 26979
rect 22764 26783 22765 26813
rect 22811 26805 22813 26815
rect 22830 26805 22837 26815
rect 22850 26805 22857 26824
rect 22873 26823 22885 26824
rect 22872 26807 22885 26823
rect 22821 26789 22823 26805
rect 22840 26789 22857 26805
rect 22746 26770 22763 26771
rect 22632 26767 22635 26768
rect 22676 26767 22680 26768
rect 22408 26747 22444 26755
rect 22520 26753 22523 26765
rect 22830 26763 22836 26789
rect 22842 26776 22857 26789
rect 22877 26776 22884 26807
rect 22906 26793 22913 26841
rect 22918 26793 22922 26816
rect 22924 26785 22931 26816
rect 22933 26793 22934 26816
rect 22936 26793 22943 26841
rect 22972 26833 22976 26841
rect 23000 26833 23006 26841
rect 23026 26833 23030 26841
rect 23052 26833 23061 26841
rect 23075 26833 23088 26841
rect 23100 26833 23102 26979
rect 23144 26978 23150 26979
rect 23137 26841 23140 26851
rect 23148 26841 23150 26978
rect 23196 26903 23198 26979
rect 23209 26977 23215 26979
rect 23218 26970 23225 26979
rect 23220 26903 23222 26970
rect 23196 26901 23227 26903
rect 23116 26833 23120 26841
rect 23144 26833 23150 26841
rect 23170 26833 23174 26841
rect 22945 26793 22949 26816
rect 22951 26785 22958 26816
rect 22960 26793 22961 26816
rect 22496 26747 22544 26753
rect 22602 26747 22613 26755
rect 22443 26737 22444 26747
rect 22468 26745 22469 26747
rect 22462 26737 22469 26745
rect 22520 26743 22523 26747
rect 22394 26697 22410 26705
rect 22384 26685 22392 26695
rect 22394 26689 22403 26697
rect 22418 26687 22420 26715
rect 22443 26689 22451 26737
rect 22468 26697 22469 26737
rect 22489 26689 22496 26737
rect 22506 26727 22522 26737
rect 22582 26735 22589 26745
rect 22632 26735 22638 26755
rect 22646 26737 22655 26745
rect 22658 26737 22665 26755
rect 22710 26747 22727 26755
rect 22737 26747 22750 26755
rect 22748 26746 22750 26747
rect 22582 26719 22598 26735
rect 22560 26693 22566 26699
rect 22658 26697 22667 26737
rect 22720 26697 22731 26737
rect 22749 26697 22750 26746
rect 22803 26737 22809 26755
rect 22815 26747 22823 26759
rect 22860 26755 22867 26776
rect 22826 26751 22850 26755
rect 22857 26751 22868 26755
rect 22826 26747 22839 26751
rect 22815 26745 22825 26747
rect 22830 26745 22836 26747
rect 22860 26745 22867 26751
rect 22878 26745 22885 26747
rect 22819 26742 22830 26745
rect 22837 26742 22844 26745
rect 22819 26737 22828 26742
rect 22849 26737 22858 26745
rect 22877 26737 22885 26745
rect 22891 26737 22895 26751
rect 22796 26697 22799 26737
rect 22801 26697 22808 26737
rect 22812 26697 22816 26737
rect 22819 26697 22826 26737
rect 22831 26697 22838 26737
rect 22842 26697 22847 26737
rect 22850 26697 22857 26737
rect 22859 26697 22868 26737
rect 22869 26697 22875 26737
rect 22877 26697 22884 26737
rect 22556 26689 22560 26693
rect 22622 26685 22628 26695
rect 22658 26689 22665 26697
rect 22796 26689 22816 26697
rect 22830 26689 22837 26697
rect 22859 26689 22867 26697
rect 22888 26689 22895 26737
rect 22906 26747 22911 26771
rect 22906 26689 22914 26747
rect 22394 26677 22402 26685
rect 22632 26677 22638 26685
rect 22862 26677 22865 26689
rect 22394 26669 22510 26677
rect 22632 26669 22639 26677
rect 22655 26669 22673 26677
rect 22689 26669 22704 26677
rect 22862 26669 22869 26677
rect 22885 26669 22906 26677
rect 22922 26669 22931 26677
rect 22982 26667 22986 26833
rect 22987 26793 22998 26833
rect 23000 26793 23007 26833
rect 23009 26793 23012 26833
rect 23014 26793 23025 26833
rect 23027 26793 23030 26833
rect 23050 26793 23061 26833
rect 23063 26793 23066 26833
rect 23068 26793 23079 26833
rect 23081 26793 23088 26833
rect 23090 26793 23093 26833
rect 22178 26650 22190 26658
rect 22206 26650 22218 26658
rect 22238 26650 22246 26658
rect 22302 26650 22310 26658
rect 22330 26650 22338 26658
rect 22362 26650 22370 26658
rect 22390 26650 22398 26658
rect 22418 26650 22426 26658
rect 22446 26650 22454 26658
rect 22457 26656 22470 26658
rect 22474 26650 22482 26658
rect 22502 26650 22510 26658
rect 22515 26656 22526 26658
rect 22530 26650 22538 26658
rect 22558 26650 22566 26658
rect 22586 26650 22594 26658
rect 22614 26650 22622 26658
rect 22642 26650 22650 26658
rect 22670 26656 22688 26658
rect 22670 26650 22678 26656
rect 22726 26650 22732 26661
rect 22754 26650 22760 26661
rect 22796 26653 22804 26661
rect 22808 26653 22816 26661
rect 22824 26653 22832 26661
rect 22836 26653 22844 26661
rect 22852 26653 22860 26661
rect 22864 26653 22872 26661
rect 22880 26653 22888 26661
rect 22892 26653 22904 26658
rect 22920 26653 22932 26658
rect 22948 26653 22960 26658
rect 22808 26652 22824 26653
rect 22836 26652 22852 26653
rect 22864 26652 22880 26653
rect 22892 26652 22900 26653
rect 22128 26642 22136 26650
rect 22162 26642 22166 26650
rect 22176 26642 22178 26650
rect 22188 26642 22192 26650
rect 22204 26642 22206 26650
rect 22164 26639 22166 26642
rect 22188 26639 22190 26642
rect 22212 26639 22214 26650
rect 22218 26642 22220 26650
rect 22246 26642 22254 26650
rect 22294 26642 22302 26650
rect 22322 26642 22330 26650
rect 22370 26642 22378 26650
rect 22398 26642 22406 26650
rect 22426 26642 22434 26650
rect 22454 26642 22462 26650
rect 22482 26642 22490 26650
rect 22510 26642 22518 26650
rect 22538 26642 22546 26650
rect 22566 26642 22574 26650
rect 22594 26642 22602 26650
rect 22622 26642 22630 26650
rect 22650 26642 22658 26650
rect 22678 26642 22686 26650
rect 22732 26645 22742 26650
rect 22760 26645 22770 26650
rect 22816 26645 22824 26652
rect 22844 26645 22852 26652
rect 22872 26645 22880 26652
rect 22904 26642 22908 26653
rect 22932 26642 22936 26653
rect 22960 26642 22964 26653
rect 22980 26650 22988 26658
rect 22988 26642 22996 26650
rect 22368 26639 22404 26642
rect 22754 26639 22788 26641
rect 23004 26639 23006 26793
rect 23007 26785 23012 26793
rect 23036 26667 23040 26793
rect 23008 26650 23016 26658
rect 23036 26650 23048 26658
rect 23052 26650 23054 26793
rect 23068 26785 23075 26793
rect 23076 26658 23078 26793
rect 23095 26785 23102 26833
rect 23104 26793 23106 26833
rect 23100 26658 23102 26785
rect 23126 26667 23130 26833
rect 23131 26793 23142 26833
rect 23144 26793 23151 26833
rect 23153 26793 23156 26833
rect 23158 26793 23169 26833
rect 23171 26793 23174 26833
rect 23064 26650 23078 26658
rect 23092 26650 23104 26658
rect 23124 26650 23132 26658
rect 23016 26642 23024 26650
rect 23048 26642 23054 26650
rect 23052 26639 23054 26642
rect 23076 26642 23080 26650
rect 23076 26639 23078 26642
rect 23100 26639 23102 26650
rect 23104 26642 23108 26650
rect 23132 26642 23140 26650
rect 23148 26639 23150 26793
rect 23151 26785 23156 26793
rect 23180 26667 23184 26793
rect 23196 26658 23198 26901
rect 23200 26667 23206 26841
rect 23220 26833 23222 26901
rect 23233 26841 23236 26851
rect 23244 26841 23246 26979
rect 23282 26915 23285 26925
rect 23292 26917 23294 26979
rect 23305 26977 23310 26979
rect 23314 26953 23321 26979
rect 23292 26893 23296 26917
rect 23225 26833 23233 26841
rect 23243 26833 23246 26841
rect 23207 26793 23216 26833
rect 23218 26793 23223 26833
rect 23227 26793 23233 26833
rect 23234 26793 23250 26833
rect 23218 26785 23225 26793
rect 23244 26785 23250 26793
rect 23220 26658 23222 26785
rect 23244 26658 23246 26785
rect 23254 26667 23260 26841
rect 23264 26833 23270 26841
rect 23276 26793 23282 26833
rect 23276 26667 23280 26793
rect 23152 26650 23160 26658
rect 23180 26650 23198 26658
rect 23212 26650 23224 26658
rect 23240 26650 23252 26658
rect 23160 26642 23168 26650
rect 23196 26639 23198 26650
rect 23208 26642 23212 26650
rect 23220 26639 23222 26650
rect 23236 26642 23240 26650
rect 23244 26639 23246 26650
rect 23292 26639 23294 26893
rect 23296 26667 23302 26841
rect 23316 26833 23318 26953
rect 23329 26841 23332 26851
rect 23340 26841 23342 26979
rect 23385 26917 23391 26979
rect 23404 26969 23407 26979
rect 23412 26969 23416 26979
rect 23412 26953 23415 26969
rect 23375 26907 23380 26913
rect 23375 26903 23382 26907
rect 23385 26893 23392 26917
rect 23385 26889 23390 26893
rect 23388 26841 23390 26889
rect 23404 26891 23407 26953
rect 23404 26889 23409 26891
rect 23404 26851 23407 26889
rect 23412 26851 23414 26953
rect 23401 26841 23414 26851
rect 23321 26833 23329 26841
rect 23339 26833 23342 26841
rect 23303 26793 23312 26833
rect 23314 26793 23319 26833
rect 23323 26793 23329 26833
rect 23330 26793 23346 26833
rect 23314 26785 23321 26793
rect 23340 26785 23346 26793
rect 23316 26658 23318 26785
rect 23340 26658 23342 26785
rect 23350 26667 23356 26841
rect 23360 26833 23366 26841
rect 23388 26833 23397 26841
rect 23405 26833 23414 26841
rect 23417 26841 23421 26979
rect 23431 26841 23434 26979
rect 23372 26793 23378 26833
rect 23386 26793 23397 26833
rect 23399 26793 23402 26833
rect 23404 26793 23415 26833
rect 23417 26793 23424 26841
rect 23436 26833 23438 26979
rect 23480 26978 23486 26979
rect 23473 26841 23476 26851
rect 23484 26841 23486 26978
rect 23532 26903 23534 26979
rect 23545 26977 23551 26979
rect 23554 26970 23561 26979
rect 23556 26903 23558 26970
rect 23532 26901 23563 26903
rect 23452 26833 23456 26841
rect 23480 26833 23486 26841
rect 23506 26833 23510 26841
rect 23426 26793 23429 26833
rect 23372 26667 23376 26793
rect 23308 26650 23318 26658
rect 23336 26650 23344 26658
rect 23368 26650 23384 26658
rect 23300 26642 23308 26650
rect 23316 26639 23318 26650
rect 23328 26642 23336 26650
rect 23340 26639 23342 26650
rect 23388 26639 23390 26793
rect 23404 26785 23411 26793
rect 23412 26658 23414 26793
rect 23431 26785 23438 26833
rect 23440 26793 23442 26833
rect 23436 26658 23438 26785
rect 23462 26667 23466 26833
rect 23467 26793 23478 26833
rect 23480 26793 23487 26833
rect 23489 26793 23492 26833
rect 23494 26793 23505 26833
rect 23507 26793 23510 26833
rect 23400 26650 23414 26658
rect 23428 26650 23440 26658
rect 23460 26650 23468 26658
rect 23396 26642 23400 26650
rect 23412 26639 23414 26650
rect 23424 26642 23428 26650
rect 23436 26639 23438 26650
rect 23468 26642 23476 26650
rect 23484 26639 23486 26793
rect 23487 26785 23492 26793
rect 23516 26667 23520 26793
rect 23532 26658 23534 26901
rect 23536 26667 23542 26841
rect 23556 26833 23558 26901
rect 23569 26841 23572 26851
rect 23580 26841 23582 26979
rect 23618 26915 23621 26925
rect 23628 26917 23630 26979
rect 23641 26977 23646 26979
rect 23650 26953 23657 26979
rect 23628 26893 23632 26917
rect 23561 26833 23569 26841
rect 23579 26833 23582 26841
rect 23543 26793 23552 26833
rect 23554 26793 23559 26833
rect 23563 26793 23569 26833
rect 23570 26793 23586 26833
rect 23554 26785 23561 26793
rect 23580 26785 23586 26793
rect 23556 26658 23558 26785
rect 23580 26658 23582 26785
rect 23590 26667 23596 26841
rect 23600 26833 23606 26841
rect 23612 26793 23618 26833
rect 23612 26667 23616 26793
rect 23488 26650 23496 26658
rect 23516 26650 23534 26658
rect 23548 26650 23560 26658
rect 23576 26650 23588 26658
rect 23496 26642 23504 26650
rect 23532 26639 23534 26650
rect 23544 26642 23548 26650
rect 23556 26639 23558 26650
rect 23572 26642 23576 26650
rect 23580 26639 23582 26650
rect 23628 26639 23630 26893
rect 23632 26667 23638 26841
rect 23652 26833 23654 26953
rect 23665 26841 23668 26851
rect 23676 26841 23678 26979
rect 23721 26917 23727 26979
rect 23740 26969 23743 26979
rect 23748 26969 23752 26979
rect 23748 26953 23751 26969
rect 23711 26907 23716 26913
rect 23711 26903 23718 26907
rect 23721 26893 23728 26917
rect 23721 26889 23726 26893
rect 23724 26841 23726 26889
rect 23740 26891 23743 26953
rect 23740 26889 23745 26891
rect 23740 26851 23743 26889
rect 23748 26851 23750 26953
rect 23737 26841 23750 26851
rect 23657 26833 23665 26841
rect 23675 26833 23678 26841
rect 23639 26793 23648 26833
rect 23650 26793 23655 26833
rect 23659 26793 23665 26833
rect 23666 26793 23682 26833
rect 23650 26785 23657 26793
rect 23676 26785 23682 26793
rect 23652 26658 23654 26785
rect 23676 26658 23678 26785
rect 23686 26667 23692 26841
rect 23696 26833 23702 26841
rect 23724 26833 23733 26841
rect 23741 26833 23750 26841
rect 23753 26841 23757 26979
rect 23767 26841 23770 26979
rect 23708 26793 23714 26833
rect 23722 26793 23733 26833
rect 23735 26793 23738 26833
rect 23740 26793 23751 26833
rect 23753 26793 23760 26841
rect 23772 26833 23774 26979
rect 23816 26978 23822 26979
rect 23809 26841 23812 26851
rect 23820 26841 23822 26978
rect 23855 26903 23860 26913
rect 23868 26903 23870 26979
rect 23888 26972 23897 26979
rect 23865 26889 23870 26903
rect 23868 26843 23870 26889
rect 23788 26833 23792 26841
rect 23816 26833 23822 26841
rect 23842 26833 23846 26841
rect 23762 26793 23765 26833
rect 23708 26667 23712 26793
rect 23644 26650 23654 26658
rect 23672 26650 23680 26658
rect 23704 26650 23720 26658
rect 23636 26642 23644 26650
rect 23652 26639 23654 26650
rect 23664 26642 23672 26650
rect 23676 26639 23678 26650
rect 23724 26639 23726 26793
rect 23740 26785 23747 26793
rect 23748 26658 23750 26793
rect 23767 26785 23774 26833
rect 23776 26793 23778 26833
rect 23772 26658 23774 26785
rect 23798 26667 23802 26833
rect 23803 26793 23814 26833
rect 23816 26793 23823 26833
rect 23825 26793 23828 26833
rect 23830 26793 23841 26833
rect 23843 26793 23846 26833
rect 23736 26650 23750 26658
rect 23764 26650 23776 26658
rect 23796 26650 23804 26658
rect 23732 26642 23736 26650
rect 23748 26639 23750 26650
rect 23760 26642 23764 26650
rect 23772 26639 23774 26650
rect 23804 26642 23812 26650
rect 23820 26639 23822 26793
rect 23823 26785 23828 26793
rect 23852 26667 23856 26793
rect 23868 26791 23878 26843
rect 23886 26839 23889 26849
rect 23892 26833 23894 26972
rect 23897 26839 23904 26972
rect 23905 26953 23908 26963
rect 23916 26953 23918 26979
rect 23915 26937 23918 26953
rect 23879 26791 23885 26833
rect 23824 26650 23832 26658
rect 23852 26650 23866 26658
rect 23868 26650 23870 26791
rect 23887 26785 23894 26833
rect 23896 26785 23905 26839
rect 23916 26833 23918 26937
rect 23931 26895 23933 26899
rect 23941 26881 23943 26895
rect 23906 26791 23912 26833
rect 23914 26785 23921 26833
rect 23923 26791 23932 26843
rect 23945 26791 23949 26849
rect 23962 26831 23966 26839
rect 23950 26791 23961 26831
rect 23963 26791 23966 26831
rect 23892 26658 23894 26785
rect 23897 26783 23904 26785
rect 23916 26658 23918 26785
rect 23945 26783 23948 26791
rect 23972 26667 23976 26791
rect 23882 26650 23894 26658
rect 23910 26650 23922 26658
rect 23942 26650 23950 26658
rect 23832 26642 23840 26650
rect 23866 26642 23870 26650
rect 23880 26642 23882 26650
rect 23892 26642 23896 26650
rect 23908 26642 23910 26650
rect 23868 26639 23870 26642
rect 23892 26639 23894 26642
rect 23916 26639 23918 26650
rect 23922 26642 23924 26650
rect 23950 26642 23958 26650
rect 23988 26639 23990 26979
rect 24012 26977 24026 26979
rect 24012 26969 24014 26977
rect 24011 26961 24016 26969
rect 24012 26955 24016 26961
rect 24010 26929 24017 26955
rect 23992 26667 23998 26841
rect 24012 26831 24014 26929
rect 24025 26841 24028 26851
rect 24036 26841 24038 26979
rect 24084 26917 24086 26979
rect 24087 26953 24103 26964
rect 24087 26917 24093 26953
rect 24084 26916 24093 26917
rect 24113 26916 24115 26964
rect 24084 26893 24088 26916
rect 24017 26831 24025 26841
rect 24035 26831 24038 26841
rect 23999 26793 24008 26831
rect 24010 26793 24015 26831
rect 24019 26793 24025 26831
rect 24026 26793 24042 26831
rect 24010 26785 24017 26793
rect 24036 26785 24042 26793
rect 24012 26658 24014 26785
rect 24036 26658 24038 26785
rect 24046 26667 24052 26841
rect 24056 26833 24062 26841
rect 24068 26793 24074 26833
rect 24068 26667 24072 26793
rect 24004 26650 24014 26658
rect 24032 26650 24042 26658
rect 23998 26642 24004 26650
rect 24012 26639 24014 26650
rect 24026 26642 24032 26650
rect 24036 26639 24038 26650
rect 24084 26639 24086 26893
rect 24132 26658 24134 26979
rect 24163 26916 24175 26956
rect 24225 26908 24227 26956
rect 24228 26851 24230 26979
rect 24247 26908 24251 26956
rect 24217 26841 24220 26851
rect 24227 26667 24230 26851
rect 24246 26841 24251 26851
rect 24228 26658 24230 26667
rect 24252 26658 24254 26979
rect 24296 26978 24302 26979
rect 24289 26841 24292 26851
rect 24300 26841 24302 26978
rect 24335 26903 24340 26913
rect 24348 26903 24350 26979
rect 24368 26972 24377 26979
rect 24345 26889 24350 26903
rect 24348 26843 24350 26889
rect 24256 26667 24261 26841
rect 24268 26833 24272 26841
rect 24296 26833 24302 26841
rect 24322 26833 24326 26841
rect 24278 26667 24282 26833
rect 24283 26793 24294 26833
rect 24296 26793 24303 26833
rect 24305 26793 24308 26833
rect 24310 26793 24321 26833
rect 24323 26793 24326 26833
rect 24098 26650 24108 26658
rect 24126 26650 24136 26658
rect 24158 26650 24166 26658
rect 24186 26650 24200 26658
rect 24216 26650 24230 26658
rect 24244 26650 24256 26658
rect 24276 26650 24284 26658
rect 24092 26642 24098 26650
rect 24120 26642 24126 26650
rect 24132 26639 24134 26650
rect 24166 26642 24174 26650
rect 24200 26642 24202 26650
rect 24214 26642 24216 26650
rect 24228 26639 24230 26650
rect 24242 26642 24244 26650
rect 24252 26639 24254 26650
rect 24256 26642 24258 26650
rect 24284 26642 24292 26650
rect 24300 26639 24302 26793
rect 24303 26785 24308 26793
rect 24332 26667 24336 26793
rect 24348 26791 24358 26843
rect 24366 26839 24369 26849
rect 24372 26833 24374 26972
rect 24377 26839 24384 26972
rect 24385 26953 24388 26963
rect 24396 26953 24398 26979
rect 24395 26937 24398 26953
rect 24359 26791 24365 26833
rect 24304 26650 24312 26658
rect 24332 26650 24346 26658
rect 24348 26650 24350 26791
rect 24367 26785 24374 26833
rect 24376 26785 24385 26839
rect 24396 26833 24398 26937
rect 24411 26895 24413 26899
rect 24421 26881 24423 26895
rect 24386 26791 24392 26833
rect 24394 26785 24401 26833
rect 24403 26791 24412 26843
rect 24425 26791 24429 26849
rect 24442 26831 24446 26839
rect 24430 26791 24441 26831
rect 24443 26791 24446 26831
rect 24372 26658 24374 26785
rect 24377 26783 24384 26785
rect 24396 26658 24398 26785
rect 24425 26783 24428 26791
rect 24452 26667 24456 26791
rect 24362 26650 24374 26658
rect 24390 26650 24402 26658
rect 24422 26650 24430 26658
rect 24312 26642 24320 26650
rect 24346 26642 24350 26650
rect 24360 26642 24362 26650
rect 24372 26642 24376 26650
rect 24388 26642 24390 26650
rect 24348 26639 24350 26642
rect 24372 26639 24374 26642
rect 24396 26639 24398 26650
rect 24402 26642 24404 26650
rect 24430 26642 24438 26650
rect 24468 26639 24470 26979
rect 24492 26977 24506 26979
rect 24492 26969 24494 26977
rect 24491 26961 24496 26969
rect 24492 26955 24496 26961
rect 24490 26929 24497 26955
rect 24472 26667 24478 26841
rect 24492 26831 24494 26929
rect 24505 26841 24508 26851
rect 24516 26841 24518 26979
rect 24561 26917 24567 26979
rect 24580 26969 24583 26979
rect 24588 26969 24592 26979
rect 24588 26953 24591 26969
rect 24551 26907 24556 26913
rect 24551 26903 24558 26907
rect 24561 26893 24568 26917
rect 24561 26889 24566 26893
rect 24564 26841 24566 26889
rect 24580 26891 24583 26953
rect 24580 26889 24585 26891
rect 24580 26851 24583 26889
rect 24588 26851 24590 26953
rect 24577 26841 24590 26851
rect 24497 26831 24505 26841
rect 24515 26831 24518 26841
rect 24479 26793 24488 26831
rect 24490 26793 24495 26831
rect 24499 26793 24505 26831
rect 24506 26793 24522 26831
rect 24490 26785 24497 26793
rect 24516 26785 24522 26793
rect 24492 26658 24494 26785
rect 24516 26658 24518 26785
rect 24526 26667 24532 26841
rect 24536 26833 24542 26841
rect 24564 26833 24573 26841
rect 24581 26833 24590 26841
rect 24593 26841 24597 26979
rect 24607 26841 24610 26979
rect 24548 26793 24554 26833
rect 24562 26793 24573 26833
rect 24575 26793 24578 26833
rect 24580 26793 24591 26833
rect 24593 26793 24600 26841
rect 24612 26833 24614 26979
rect 24656 26978 24662 26979
rect 24649 26841 24652 26851
rect 24660 26841 24662 26978
rect 24695 26903 24700 26913
rect 24708 26903 24710 26979
rect 24728 26972 24737 26979
rect 24705 26889 24710 26903
rect 24708 26843 24710 26889
rect 24628 26833 24632 26841
rect 24656 26833 24662 26841
rect 24682 26833 24686 26841
rect 24602 26793 24605 26833
rect 24548 26667 24552 26793
rect 24484 26650 24494 26658
rect 24512 26650 24522 26658
rect 24544 26650 24560 26658
rect 24478 26642 24484 26650
rect 24492 26639 24494 26650
rect 24506 26642 24512 26650
rect 24516 26639 24518 26650
rect 24564 26639 24566 26793
rect 24580 26785 24587 26793
rect 24588 26658 24590 26793
rect 24607 26785 24614 26833
rect 24616 26793 24618 26833
rect 24612 26658 24614 26785
rect 24638 26667 24642 26833
rect 24643 26793 24654 26833
rect 24656 26793 24663 26833
rect 24665 26793 24668 26833
rect 24670 26793 24681 26833
rect 24683 26793 24686 26833
rect 24576 26650 24590 26658
rect 24604 26650 24616 26658
rect 24636 26650 24644 26658
rect 24572 26642 24576 26650
rect 24588 26639 24590 26650
rect 24600 26642 24604 26650
rect 24612 26639 24614 26650
rect 24644 26642 24652 26650
rect 24660 26639 24662 26793
rect 24663 26785 24668 26793
rect 24692 26667 24696 26793
rect 24708 26791 24718 26843
rect 24726 26839 24729 26849
rect 24732 26833 24734 26972
rect 24737 26839 24744 26972
rect 24745 26953 24748 26963
rect 24756 26953 24758 26979
rect 24755 26937 24758 26953
rect 24719 26791 24725 26833
rect 24664 26650 24672 26658
rect 24692 26650 24706 26658
rect 24708 26650 24710 26791
rect 24727 26785 24734 26833
rect 24736 26785 24745 26839
rect 24756 26833 24758 26937
rect 24815 26903 24820 26913
rect 24828 26903 24830 26979
rect 24851 26977 24864 26979
rect 24851 26972 24854 26977
rect 24771 26895 24773 26899
rect 24781 26881 24783 26895
rect 24825 26889 24830 26903
rect 24746 26791 24752 26833
rect 24754 26785 24761 26833
rect 24763 26791 24772 26843
rect 24785 26791 24789 26849
rect 24828 26841 24830 26889
rect 24852 26969 24854 26972
rect 24852 26945 24856 26969
rect 24802 26831 24806 26839
rect 24790 26791 24801 26831
rect 24803 26791 24806 26831
rect 24828 26791 24838 26841
rect 24846 26839 24849 26849
rect 24852 26831 24854 26945
rect 24857 26839 24864 26972
rect 24865 26953 24868 26963
rect 24876 26953 24878 26979
rect 24945 26964 24950 26979
rect 24875 26937 24878 26953
rect 24839 26791 24845 26831
rect 24732 26658 24734 26785
rect 24737 26783 24744 26785
rect 24756 26658 24758 26785
rect 24785 26783 24788 26791
rect 24812 26667 24816 26791
rect 24722 26650 24734 26658
rect 24750 26650 24762 26658
rect 24782 26650 24790 26658
rect 24810 26650 24826 26658
rect 24672 26642 24680 26650
rect 24706 26642 24710 26650
rect 24720 26642 24722 26650
rect 24732 26642 24736 26650
rect 24748 26642 24750 26650
rect 24708 26639 24710 26642
rect 24732 26639 24734 26642
rect 24756 26639 24758 26650
rect 24762 26642 24764 26650
rect 24790 26642 24798 26650
rect 24828 26639 24830 26791
rect 24847 26783 24854 26831
rect 24856 26783 24865 26839
rect 24876 26831 24878 26937
rect 24935 26903 24940 26913
rect 24948 26903 24950 26964
rect 24964 26945 24967 26979
rect 24972 26969 24974 26979
rect 24972 26945 24976 26969
rect 24891 26895 24893 26899
rect 24901 26881 24903 26895
rect 24945 26889 24950 26903
rect 24866 26791 24872 26831
rect 24874 26783 24881 26831
rect 24883 26791 24892 26841
rect 24905 26791 24909 26849
rect 24948 26841 24950 26889
rect 24964 26851 24967 26929
rect 24961 26841 24967 26851
rect 24972 26891 24974 26945
rect 24977 26891 24981 26979
rect 24972 26841 24981 26891
rect 24991 26841 24994 26979
rect 24922 26831 24926 26839
rect 24948 26831 24957 26841
rect 24971 26831 24984 26841
rect 24996 26831 24998 26979
rect 25040 26978 25046 26979
rect 25033 26841 25036 26851
rect 25044 26841 25046 26978
rect 25012 26833 25016 26841
rect 25040 26833 25046 26841
rect 25066 26833 25070 26841
rect 24910 26791 24921 26831
rect 24923 26791 24926 26831
rect 24946 26793 24957 26831
rect 24959 26793 24962 26831
rect 24964 26793 24975 26831
rect 24977 26793 24984 26831
rect 24986 26793 24989 26831
rect 24905 26783 24908 26791
rect 24852 26658 24854 26783
rect 24876 26658 24878 26783
rect 24932 26667 24936 26791
rect 24842 26650 24854 26658
rect 24870 26650 24882 26658
rect 24902 26650 24910 26658
rect 24930 26650 24944 26658
rect 24838 26642 24842 26650
rect 24852 26639 24854 26650
rect 24866 26642 24870 26650
rect 24876 26639 24878 26650
rect 24910 26642 24918 26650
rect 24944 26642 24946 26650
rect 24948 26639 24950 26793
rect 24964 26785 24971 26793
rect 24972 26658 24974 26793
rect 24991 26785 24998 26831
rect 25000 26793 25002 26831
rect 24996 26658 24998 26785
rect 25022 26667 25026 26833
rect 25027 26793 25038 26833
rect 25040 26793 25047 26833
rect 25049 26793 25052 26833
rect 25054 26793 25065 26833
rect 25067 26793 25070 26833
rect 24960 26650 24974 26658
rect 24988 26650 25000 26658
rect 25020 26650 25028 26658
rect 24958 26642 24960 26650
rect 24972 26639 24974 26650
rect 24986 26642 24988 26650
rect 24996 26639 24998 26650
rect 25000 26642 25002 26650
rect 25028 26642 25036 26650
rect 25044 26639 25046 26793
rect 25047 26785 25052 26793
rect 25076 26667 25080 26793
rect 25048 26650 25056 26658
rect 25076 26650 25090 26658
rect 25092 26650 25094 26979
rect 25110 26970 25111 26974
rect 25095 26916 25101 26964
rect 25121 26916 25123 26964
rect 25140 26658 25142 26979
rect 25171 26916 25183 26956
rect 25226 26916 25233 26964
rect 25235 26916 25241 26956
rect 25243 26908 25250 26956
rect 25260 26658 25262 26979
rect 25355 26972 25358 26979
rect 25356 26956 25358 26972
rect 25380 26966 25382 26979
rect 25291 26916 25303 26956
rect 25353 26908 25358 26956
rect 25369 26953 25372 26963
rect 25378 26953 25379 26956
rect 25380 26953 25389 26966
rect 25378 26937 25382 26953
rect 25378 26908 25379 26937
rect 25356 26849 25358 26908
rect 25355 26791 25359 26849
rect 25356 26658 25358 26791
rect 25380 26658 25382 26937
rect 25395 26895 25397 26899
rect 25387 26791 25389 26889
rect 25405 26881 25407 26895
rect 25409 26791 25413 26849
rect 25426 26831 25430 26839
rect 25414 26791 25425 26831
rect 25427 26791 25430 26831
rect 25409 26783 25412 26791
rect 25436 26667 25440 26791
rect 25106 26650 25118 26658
rect 25134 26650 25146 26658
rect 25166 26650 25174 26658
rect 25194 26650 25210 26658
rect 25226 26650 25238 26658
rect 25254 26650 25266 26658
rect 25286 26650 25294 26658
rect 25314 26650 25330 26658
rect 25346 26650 25358 26658
rect 25374 26650 25386 26658
rect 25406 26650 25414 26658
rect 25056 26642 25064 26650
rect 25090 26642 25094 26650
rect 25104 26642 25106 26650
rect 25118 26642 25120 26650
rect 25132 26642 25134 26650
rect 25092 26639 25094 26642
rect 25140 26639 25142 26650
rect 25146 26642 25148 26650
rect 25174 26642 25182 26650
rect 25222 26642 25226 26650
rect 25250 26642 25254 26650
rect 25260 26639 25262 26650
rect 25294 26642 25302 26650
rect 25342 26642 25346 26650
rect 25356 26639 25358 26650
rect 25370 26642 25374 26650
rect 25380 26639 25382 26650
rect 25414 26642 25422 26650
rect 25452 26639 25454 26979
rect 25476 26977 25490 26979
rect 25476 26969 25478 26977
rect 25475 26961 25480 26969
rect 25476 26955 25480 26961
rect 25474 26929 25481 26955
rect 25456 26667 25462 26841
rect 25476 26831 25478 26929
rect 25489 26841 25492 26851
rect 25500 26841 25502 26979
rect 25545 26917 25551 26979
rect 25564 26969 25567 26979
rect 25572 26969 25576 26979
rect 25572 26953 25575 26969
rect 25535 26907 25540 26913
rect 25535 26903 25542 26907
rect 25545 26893 25552 26917
rect 25545 26889 25550 26893
rect 25548 26841 25550 26889
rect 25564 26891 25567 26953
rect 25564 26889 25569 26891
rect 25564 26851 25567 26889
rect 25572 26851 25574 26953
rect 25561 26841 25574 26851
rect 25481 26831 25489 26841
rect 25499 26831 25502 26841
rect 25463 26793 25472 26831
rect 25474 26793 25479 26831
rect 25483 26793 25489 26831
rect 25490 26793 25506 26831
rect 25474 26785 25481 26793
rect 25500 26785 25506 26793
rect 25476 26658 25478 26785
rect 25500 26658 25502 26785
rect 25510 26667 25516 26841
rect 25520 26833 25526 26841
rect 25548 26833 25557 26841
rect 25565 26833 25574 26841
rect 25577 26841 25581 26979
rect 25591 26841 25594 26979
rect 25532 26793 25538 26833
rect 25546 26793 25557 26833
rect 25559 26793 25562 26833
rect 25564 26793 25575 26833
rect 25577 26793 25584 26841
rect 25596 26833 25598 26979
rect 25640 26978 25646 26979
rect 25633 26841 25636 26851
rect 25644 26841 25646 26978
rect 25802 26882 25809 26979
rect 25852 26976 25855 26979
rect 25928 26968 25931 26979
rect 25969 26970 25972 26979
rect 25987 26978 26073 26979
rect 26022 26960 26025 26961
rect 25832 26952 25838 26960
rect 25845 26952 25859 26960
rect 25919 26952 25928 26953
rect 25988 26952 25990 26960
rect 25997 26952 26031 26960
rect 25852 26950 25855 26952
rect 25928 26950 25931 26952
rect 25838 26902 25845 26950
rect 25848 26902 25849 26942
rect 25833 26894 25842 26902
rect 25852 26894 25859 26942
rect 25870 26902 25877 26950
rect 25921 26947 25935 26950
rect 25928 26942 25935 26947
rect 25909 26902 25912 26942
rect 25864 26894 25909 26902
rect 25914 26894 25921 26942
rect 25929 26894 25935 26942
rect 25986 26902 25988 26942
rect 25990 26902 25997 26950
rect 26017 26947 26038 26950
rect 26031 26942 26038 26947
rect 26084 26942 26088 26978
rect 26005 26902 26006 26942
rect 25955 26894 25962 26902
rect 26008 26894 26015 26942
rect 26019 26902 26023 26942
rect 26031 26902 26035 26942
rect 26062 26902 26063 26942
rect 26038 26894 26045 26902
rect 26071 26894 26078 26942
rect 25852 26882 25855 26894
rect 25928 26892 25935 26894
rect 25928 26882 25931 26892
rect 25792 26874 25864 26882
rect 25909 26874 25986 26882
rect 25802 26872 25809 26874
rect 25812 26856 25816 26862
rect 25612 26833 25616 26841
rect 25640 26833 25646 26841
rect 25666 26833 25670 26841
rect 25586 26793 25589 26833
rect 25532 26667 25536 26793
rect 25468 26650 25478 26658
rect 25496 26650 25506 26658
rect 25528 26650 25544 26658
rect 25462 26642 25468 26650
rect 25476 26639 25478 26650
rect 25490 26642 25496 26650
rect 25500 26639 25502 26650
rect 25548 26639 25550 26793
rect 25564 26785 25571 26793
rect 25572 26658 25574 26793
rect 25591 26785 25598 26833
rect 25600 26793 25602 26833
rect 25596 26658 25598 26785
rect 25622 26667 25626 26833
rect 25627 26793 25638 26833
rect 25640 26793 25647 26833
rect 25649 26793 25652 26833
rect 25654 26793 25665 26833
rect 25667 26793 25670 26833
rect 25560 26650 25574 26658
rect 25588 26650 25600 26658
rect 25620 26650 25628 26658
rect 25556 26642 25560 26650
rect 25572 26639 25574 26650
rect 25584 26642 25588 26650
rect 25596 26639 25598 26650
rect 25628 26642 25636 26650
rect 25644 26639 25646 26793
rect 25647 26785 25652 26793
rect 25676 26667 25680 26793
rect 25700 26667 25702 26843
rect 25728 26824 25733 26833
rect 25703 26785 25716 26824
rect 25726 26785 25728 26824
rect 25730 26785 25733 26824
rect 25736 26785 25746 26824
rect 25802 26816 25809 26856
rect 25852 26841 25855 26874
rect 25856 26864 25859 26874
rect 25866 26854 25869 26864
rect 25866 26848 25882 26854
rect 25910 26848 25922 26854
rect 25824 26824 25828 26834
rect 25838 26826 25860 26834
rect 25838 26825 25854 26826
rect 25928 26824 25931 26874
rect 25954 26854 26076 26859
rect 25980 26839 25998 26846
rect 25935 26826 25955 26834
rect 26084 26826 26088 26894
rect 25834 26820 25852 26824
rect 25721 26777 25726 26785
rect 25794 26768 25801 26816
rect 25834 26776 25840 26820
rect 25870 26776 25877 26824
rect 25928 26816 25936 26824
rect 25990 26816 25997 26824
rect 25910 26776 25912 26816
rect 25812 26768 25828 26775
rect 25834 26768 25838 26776
rect 25914 26768 25921 26816
rect 25929 26768 25936 26816
rect 25972 26777 25980 26816
rect 25972 26776 25988 26777
rect 25802 26705 25809 26768
rect 25928 26765 25936 26768
rect 25955 26765 25962 26776
rect 25980 26768 25988 26776
rect 26008 26768 26015 26816
rect 26017 26776 26021 26816
rect 26031 26776 26033 26824
rect 26038 26768 26045 26816
rect 26050 26778 26056 26816
rect 26084 26778 26091 26826
rect 26093 26778 26097 26816
rect 26071 26768 26078 26778
rect 26154 26771 26158 26818
rect 26227 26815 26230 26841
rect 26238 26815 26244 26979
rect 26268 26824 26275 26979
rect 26426 26882 26433 26979
rect 26476 26976 26479 26979
rect 26552 26968 26555 26979
rect 26593 26970 26596 26979
rect 26611 26978 26697 26979
rect 26646 26960 26649 26961
rect 26456 26952 26462 26960
rect 26469 26952 26483 26960
rect 26543 26952 26552 26953
rect 26612 26952 26614 26960
rect 26621 26952 26655 26960
rect 26476 26950 26479 26952
rect 26552 26950 26555 26952
rect 26462 26902 26469 26950
rect 26472 26902 26473 26942
rect 26457 26894 26466 26902
rect 26476 26894 26483 26942
rect 26494 26902 26501 26950
rect 26545 26947 26559 26950
rect 26552 26942 26559 26947
rect 26533 26902 26536 26942
rect 26488 26894 26533 26902
rect 26538 26894 26545 26942
rect 26553 26894 26559 26942
rect 26610 26902 26612 26942
rect 26614 26902 26621 26950
rect 26641 26947 26662 26950
rect 26655 26942 26662 26947
rect 26708 26942 26712 26978
rect 26629 26902 26630 26942
rect 26579 26894 26586 26902
rect 26632 26894 26639 26942
rect 26643 26902 26647 26942
rect 26655 26902 26659 26942
rect 26686 26902 26687 26942
rect 26662 26894 26669 26902
rect 26695 26894 26702 26942
rect 26476 26882 26479 26894
rect 26552 26892 26559 26894
rect 26552 26882 26555 26892
rect 26416 26874 26488 26882
rect 26533 26874 26610 26882
rect 26426 26872 26433 26874
rect 26436 26856 26440 26862
rect 26172 26783 26173 26813
rect 26219 26805 26221 26815
rect 26238 26805 26245 26815
rect 26258 26805 26265 26824
rect 26281 26823 26293 26824
rect 26280 26807 26293 26823
rect 26324 26816 26326 26824
rect 26344 26816 26350 26824
rect 26426 26816 26433 26856
rect 26476 26841 26479 26874
rect 26480 26864 26483 26874
rect 26490 26854 26493 26864
rect 26490 26848 26506 26854
rect 26534 26848 26546 26854
rect 26448 26824 26452 26834
rect 26462 26826 26484 26834
rect 26462 26825 26478 26826
rect 26552 26824 26555 26874
rect 26578 26854 26700 26859
rect 26604 26839 26622 26846
rect 26559 26826 26579 26834
rect 26708 26826 26712 26894
rect 26458 26820 26476 26824
rect 26229 26789 26231 26805
rect 26248 26789 26265 26805
rect 26154 26770 26171 26771
rect 26040 26767 26043 26768
rect 26084 26767 26088 26768
rect 25816 26747 25852 26755
rect 25928 26753 25931 26765
rect 26238 26763 26244 26789
rect 26250 26776 26265 26789
rect 26285 26776 26292 26807
rect 26324 26776 26340 26816
rect 26350 26776 26351 26816
rect 26353 26776 26357 26816
rect 26360 26776 26369 26816
rect 25904 26747 25952 26753
rect 26010 26747 26021 26755
rect 25851 26737 25852 26747
rect 25876 26745 25877 26747
rect 25870 26737 25877 26745
rect 25928 26743 25931 26747
rect 25802 26697 25818 26705
rect 25792 26685 25800 26695
rect 25802 26689 25811 26697
rect 25826 26687 25828 26715
rect 25851 26689 25859 26737
rect 25876 26697 25877 26737
rect 25897 26689 25904 26737
rect 25914 26727 25930 26737
rect 25990 26735 25997 26745
rect 26040 26735 26046 26755
rect 26054 26737 26063 26745
rect 26066 26737 26073 26755
rect 26118 26747 26135 26755
rect 26145 26747 26158 26755
rect 26156 26746 26158 26747
rect 25990 26719 26006 26735
rect 25968 26693 25974 26699
rect 26066 26697 26075 26737
rect 26128 26697 26139 26737
rect 26157 26697 26158 26746
rect 26211 26737 26217 26755
rect 26223 26747 26231 26759
rect 26268 26755 26275 26776
rect 26340 26768 26342 26775
rect 26351 26768 26357 26776
rect 26418 26768 26425 26816
rect 26458 26776 26464 26820
rect 26494 26776 26501 26824
rect 26552 26816 26560 26824
rect 26614 26816 26621 26824
rect 26534 26776 26536 26816
rect 26436 26768 26452 26775
rect 26458 26768 26462 26776
rect 26538 26768 26545 26816
rect 26553 26768 26560 26816
rect 26596 26777 26604 26816
rect 26596 26776 26612 26777
rect 26234 26751 26258 26755
rect 26265 26751 26276 26755
rect 26234 26747 26247 26751
rect 26223 26745 26233 26747
rect 26238 26745 26244 26747
rect 26268 26745 26275 26751
rect 26286 26745 26293 26747
rect 26227 26742 26238 26745
rect 26245 26742 26252 26745
rect 26227 26737 26236 26742
rect 26257 26737 26266 26745
rect 26285 26737 26293 26745
rect 26299 26737 26303 26751
rect 26204 26697 26207 26737
rect 26209 26697 26216 26737
rect 26220 26697 26224 26737
rect 26227 26697 26234 26737
rect 26239 26697 26246 26737
rect 26250 26697 26255 26737
rect 26258 26697 26265 26737
rect 26267 26697 26276 26737
rect 26277 26697 26283 26737
rect 26285 26697 26292 26737
rect 25964 26689 25968 26693
rect 26030 26685 26036 26695
rect 26066 26689 26073 26697
rect 26204 26689 26224 26697
rect 26238 26689 26245 26697
rect 26267 26689 26275 26697
rect 26296 26689 26303 26737
rect 26351 26713 26357 26737
rect 26350 26697 26366 26713
rect 26426 26705 26433 26768
rect 26552 26765 26560 26768
rect 26579 26765 26586 26776
rect 26604 26768 26612 26776
rect 26632 26768 26639 26816
rect 26641 26776 26645 26816
rect 26655 26776 26657 26824
rect 26662 26768 26669 26816
rect 26674 26778 26680 26816
rect 26708 26778 26715 26826
rect 26717 26778 26721 26816
rect 26695 26768 26702 26778
rect 26778 26771 26782 26818
rect 26851 26815 26854 26841
rect 26862 26815 26868 26979
rect 26892 26824 26899 26979
rect 26968 26919 26975 26967
rect 27060 26921 27062 26979
rect 27063 26969 27064 26979
rect 27063 26921 27070 26969
rect 27083 26961 27097 26969
rect 27060 26915 27070 26921
rect 26796 26783 26797 26813
rect 26843 26805 26845 26815
rect 26862 26805 26869 26815
rect 26882 26805 26889 26824
rect 26905 26823 26917 26824
rect 26904 26807 26917 26823
rect 26853 26789 26855 26805
rect 26872 26789 26889 26805
rect 26778 26770 26795 26771
rect 26664 26767 26667 26768
rect 26708 26767 26712 26768
rect 26440 26747 26476 26755
rect 26552 26753 26555 26765
rect 26862 26763 26868 26789
rect 26874 26776 26889 26789
rect 26909 26776 26916 26807
rect 26528 26747 26576 26753
rect 26634 26747 26645 26755
rect 26475 26737 26476 26747
rect 26500 26745 26501 26747
rect 26494 26737 26501 26745
rect 26552 26743 26555 26747
rect 26426 26697 26442 26705
rect 26350 26689 26352 26697
rect 26353 26689 26366 26693
rect 25802 26677 25810 26685
rect 26040 26677 26046 26685
rect 26270 26677 26273 26689
rect 26416 26685 26424 26695
rect 26426 26689 26435 26697
rect 26450 26687 26452 26715
rect 26475 26689 26483 26737
rect 26500 26697 26501 26737
rect 26521 26689 26528 26737
rect 26538 26727 26554 26737
rect 26614 26735 26621 26745
rect 26664 26735 26670 26755
rect 26678 26737 26687 26745
rect 26690 26737 26697 26755
rect 26742 26747 26759 26755
rect 26769 26747 26782 26755
rect 26780 26746 26782 26747
rect 26614 26719 26630 26735
rect 26592 26693 26598 26699
rect 26690 26697 26699 26737
rect 26752 26697 26763 26737
rect 26781 26697 26782 26746
rect 26835 26737 26841 26755
rect 26847 26747 26855 26759
rect 26892 26755 26899 26776
rect 26858 26751 26882 26755
rect 26889 26751 26900 26755
rect 26858 26747 26871 26751
rect 26847 26745 26857 26747
rect 26862 26745 26868 26747
rect 26892 26745 26899 26751
rect 26910 26745 26917 26747
rect 26851 26742 26862 26745
rect 26869 26742 26876 26745
rect 26851 26737 26860 26742
rect 26881 26737 26890 26745
rect 26909 26737 26917 26745
rect 26923 26737 26927 26751
rect 26828 26697 26831 26737
rect 26833 26697 26840 26737
rect 26844 26697 26848 26737
rect 26851 26697 26858 26737
rect 26863 26697 26870 26737
rect 26874 26697 26879 26737
rect 26882 26697 26889 26737
rect 26891 26697 26900 26737
rect 26901 26697 26907 26737
rect 26909 26697 26916 26737
rect 26588 26689 26592 26693
rect 26654 26685 26660 26695
rect 26690 26689 26697 26697
rect 26828 26689 26848 26697
rect 26862 26689 26869 26697
rect 26891 26689 26899 26697
rect 26920 26689 26927 26737
rect 26426 26677 26434 26685
rect 26664 26677 26670 26685
rect 26894 26677 26897 26689
rect 25802 26669 25918 26677
rect 26040 26669 26047 26677
rect 26063 26669 26081 26677
rect 26097 26669 26112 26677
rect 26270 26669 26277 26677
rect 26293 26669 26324 26677
rect 26426 26669 26542 26677
rect 26664 26669 26671 26677
rect 26687 26669 26705 26677
rect 26721 26669 26736 26677
rect 26894 26669 26901 26677
rect 26917 26669 26963 26677
rect 26995 26667 27003 26826
rect 25648 26650 25656 26658
rect 25710 26650 25720 26658
rect 25738 26650 25748 26658
rect 25770 26650 25778 26658
rect 25798 26650 25806 26658
rect 25826 26650 25834 26658
rect 25854 26650 25862 26658
rect 25865 26656 25878 26658
rect 25882 26650 25890 26658
rect 25910 26650 25918 26658
rect 25923 26656 25934 26658
rect 25938 26650 25946 26658
rect 25966 26650 25974 26658
rect 25994 26650 26002 26658
rect 26022 26650 26030 26658
rect 26050 26650 26058 26658
rect 26078 26656 26096 26658
rect 26078 26650 26086 26656
rect 26134 26650 26140 26661
rect 26162 26650 26168 26661
rect 26204 26653 26212 26661
rect 26216 26653 26224 26661
rect 26232 26653 26240 26661
rect 26244 26653 26252 26661
rect 26260 26653 26268 26661
rect 26272 26653 26280 26661
rect 26288 26653 26296 26661
rect 26318 26653 26328 26658
rect 26334 26653 26344 26658
rect 26346 26653 26356 26658
rect 26362 26653 26372 26658
rect 26216 26652 26232 26653
rect 26244 26652 26260 26653
rect 26272 26652 26288 26653
rect 26300 26652 26308 26653
rect 26318 26652 26334 26653
rect 26346 26652 26362 26653
rect 26374 26652 26384 26658
rect 25656 26642 25664 26650
rect 25704 26642 25710 26650
rect 25732 26642 25738 26650
rect 25778 26642 25786 26650
rect 25806 26642 25814 26650
rect 25834 26642 25842 26650
rect 25862 26642 25870 26650
rect 25890 26642 25898 26650
rect 25918 26642 25926 26650
rect 25946 26642 25954 26650
rect 25974 26642 25982 26650
rect 26002 26642 26010 26650
rect 26030 26642 26038 26650
rect 26058 26642 26066 26650
rect 26086 26642 26094 26650
rect 26140 26645 26150 26650
rect 26168 26645 26178 26650
rect 26224 26645 26232 26652
rect 26252 26645 26260 26652
rect 26280 26645 26288 26652
rect 26328 26642 26334 26652
rect 26356 26642 26362 26652
rect 26394 26650 26402 26658
rect 26422 26650 26430 26658
rect 26450 26650 26458 26658
rect 26478 26650 26486 26658
rect 26489 26656 26502 26658
rect 26506 26650 26514 26658
rect 26534 26650 26542 26658
rect 26547 26656 26558 26658
rect 26562 26650 26570 26658
rect 26590 26650 26598 26658
rect 26618 26650 26626 26658
rect 26646 26650 26654 26658
rect 26674 26650 26682 26658
rect 26702 26656 26720 26658
rect 26702 26650 26710 26656
rect 26758 26650 26764 26661
rect 26786 26650 26792 26661
rect 26828 26653 26836 26661
rect 26840 26653 26848 26661
rect 26856 26653 26864 26661
rect 26868 26653 26876 26661
rect 26884 26653 26892 26661
rect 26896 26653 26904 26661
rect 26912 26653 26920 26661
rect 27060 26658 27062 26915
rect 27071 26911 27074 26915
rect 27082 26911 27087 26959
rect 27081 26841 27087 26851
rect 27097 26841 27100 26851
rect 27108 26841 27110 26979
rect 27180 26969 27185 26979
rect 27180 26953 27183 26969
rect 27184 26967 27185 26969
rect 27184 26953 27192 26967
rect 27091 26793 27097 26841
rect 27107 26793 27110 26841
rect 27128 26833 27134 26841
rect 27108 26658 27110 26793
rect 27140 26793 27146 26833
rect 27140 26667 27144 26793
rect 27180 26658 27182 26953
rect 27185 26919 27192 26953
rect 27276 26921 27278 26979
rect 27279 26969 27280 26979
rect 27279 26921 27286 26969
rect 27299 26961 27313 26969
rect 27276 26915 27286 26921
rect 27211 26667 27220 26843
rect 27276 26658 27278 26915
rect 27287 26911 27290 26915
rect 27298 26911 27303 26959
rect 27297 26841 27303 26851
rect 27313 26841 27316 26851
rect 27324 26841 27326 26979
rect 27369 26917 27375 26979
rect 27388 26969 27391 26979
rect 27396 26969 27400 26979
rect 27396 26953 27399 26969
rect 27359 26907 27364 26913
rect 27359 26903 27366 26907
rect 27369 26893 27376 26917
rect 27369 26889 27374 26893
rect 27372 26841 27374 26889
rect 27388 26891 27391 26953
rect 27388 26889 27393 26891
rect 27388 26851 27391 26889
rect 27396 26851 27398 26953
rect 27385 26841 27398 26851
rect 27307 26793 27313 26841
rect 27323 26793 27326 26841
rect 27344 26833 27350 26841
rect 27372 26833 27381 26841
rect 27389 26833 27398 26841
rect 27401 26841 27405 26979
rect 27415 26841 27418 26979
rect 27324 26658 27326 26793
rect 27356 26793 27362 26833
rect 27370 26793 27381 26833
rect 27383 26793 27386 26833
rect 27388 26793 27399 26833
rect 27401 26793 27408 26841
rect 27420 26833 27422 26979
rect 27464 26978 27470 26979
rect 27457 26841 27460 26851
rect 27468 26841 27470 26978
rect 27516 26903 27518 26979
rect 27529 26977 27535 26979
rect 27538 26970 27545 26979
rect 27540 26903 27542 26970
rect 27516 26901 27547 26903
rect 27436 26833 27440 26841
rect 27464 26833 27470 26841
rect 27490 26833 27494 26841
rect 27410 26793 27413 26833
rect 27356 26667 27360 26793
rect 26942 26653 26952 26658
rect 26958 26653 26968 26658
rect 26970 26653 26980 26658
rect 26986 26653 26996 26658
rect 26840 26652 26856 26653
rect 26868 26652 26884 26653
rect 26896 26652 26912 26653
rect 26924 26652 26932 26653
rect 26942 26652 26958 26653
rect 26970 26652 26986 26653
rect 26998 26652 27008 26658
rect 26402 26642 26410 26650
rect 26430 26642 26438 26650
rect 26458 26642 26466 26650
rect 26486 26642 26494 26650
rect 26514 26642 26522 26650
rect 26542 26642 26550 26650
rect 26570 26642 26578 26650
rect 26598 26642 26606 26650
rect 26626 26642 26634 26650
rect 26654 26642 26662 26650
rect 26682 26642 26690 26650
rect 26710 26642 26718 26650
rect 26764 26645 26774 26650
rect 26792 26645 26802 26650
rect 26848 26645 26856 26652
rect 26876 26645 26884 26652
rect 26904 26645 26912 26652
rect 26952 26642 26958 26652
rect 26980 26642 26986 26652
rect 27018 26650 27026 26658
rect 27046 26650 27062 26658
rect 27076 26650 27088 26658
rect 27104 26650 27116 26658
rect 27174 26650 27182 26658
rect 27202 26650 27208 26658
rect 27234 26650 27242 26658
rect 27262 26650 27278 26658
rect 27292 26650 27304 26658
rect 27320 26650 27332 26658
rect 27352 26650 27368 26658
rect 27026 26642 27034 26650
rect 25776 26639 25812 26642
rect 26162 26639 26196 26641
rect 26400 26639 26436 26642
rect 26786 26639 26820 26641
rect 27060 26639 27062 26650
rect 27074 26642 27076 26650
rect 27088 26642 27090 26650
rect 27102 26642 27104 26650
rect 27108 26639 27110 26650
rect 27116 26642 27118 26650
rect 27164 26642 27174 26650
rect 27180 26639 27182 26650
rect 27192 26642 27202 26650
rect 27242 26642 27250 26650
rect 27276 26639 27278 26650
rect 27290 26642 27292 26650
rect 27304 26642 27306 26650
rect 27318 26642 27320 26650
rect 27324 26639 27326 26650
rect 27332 26642 27334 26650
rect 27372 26639 27374 26793
rect 27388 26785 27395 26793
rect 27396 26658 27398 26793
rect 27415 26785 27422 26833
rect 27424 26793 27426 26833
rect 27420 26658 27422 26785
rect 27446 26667 27450 26833
rect 27451 26793 27462 26833
rect 27464 26793 27471 26833
rect 27473 26793 27476 26833
rect 27478 26793 27489 26833
rect 27491 26793 27494 26833
rect 27384 26650 27398 26658
rect 27412 26650 27424 26658
rect 27444 26650 27452 26658
rect 27380 26642 27384 26650
rect 27396 26639 27398 26650
rect 27408 26642 27412 26650
rect 27420 26639 27422 26650
rect 27452 26642 27460 26650
rect 27468 26639 27470 26793
rect 27471 26785 27476 26793
rect 27500 26667 27504 26793
rect 27516 26658 27518 26901
rect 27520 26667 27526 26841
rect 27540 26833 27542 26901
rect 27553 26841 27556 26851
rect 27564 26841 27566 26979
rect 27610 26893 27629 26902
rect 27722 26882 27729 26979
rect 27772 26976 27775 26979
rect 27848 26968 27851 26979
rect 27889 26970 27892 26979
rect 27907 26978 27993 26979
rect 28049 26978 28054 26979
rect 27942 26960 27945 26961
rect 27752 26952 27758 26960
rect 27765 26952 27779 26960
rect 27839 26952 27848 26953
rect 27908 26952 27910 26960
rect 27917 26952 27951 26960
rect 27772 26950 27775 26952
rect 27848 26950 27851 26952
rect 27758 26902 27765 26950
rect 27768 26902 27769 26942
rect 27753 26894 27762 26902
rect 27772 26894 27779 26942
rect 27790 26902 27797 26950
rect 27841 26947 27855 26950
rect 27848 26942 27855 26947
rect 27829 26902 27832 26942
rect 27784 26894 27829 26902
rect 27834 26894 27841 26942
rect 27849 26894 27855 26942
rect 27906 26902 27908 26942
rect 27910 26902 27917 26950
rect 27937 26947 27958 26950
rect 27951 26942 27958 26947
rect 28004 26942 28008 26978
rect 27925 26902 27926 26942
rect 27875 26894 27882 26902
rect 27928 26894 27935 26942
rect 27939 26902 27943 26942
rect 27951 26902 27955 26942
rect 27982 26902 27983 26942
rect 27958 26894 27965 26902
rect 27991 26894 27998 26942
rect 28037 26894 28059 26895
rect 27772 26882 27775 26894
rect 27848 26892 27855 26894
rect 27848 26882 27851 26892
rect 27712 26874 27784 26882
rect 27829 26874 27906 26882
rect 27722 26872 27729 26874
rect 27732 26856 27736 26862
rect 27545 26833 27553 26841
rect 27563 26833 27566 26841
rect 27527 26793 27536 26833
rect 27538 26793 27543 26833
rect 27547 26793 27553 26833
rect 27554 26793 27570 26833
rect 27538 26785 27545 26793
rect 27564 26785 27570 26793
rect 27540 26658 27542 26785
rect 27564 26658 27566 26785
rect 27574 26667 27580 26841
rect 27584 26833 27590 26841
rect 27596 26793 27602 26833
rect 27596 26667 27600 26793
rect 27620 26667 27622 26843
rect 27648 26824 27653 26833
rect 27623 26785 27636 26824
rect 27646 26785 27648 26824
rect 27650 26785 27653 26824
rect 27656 26785 27666 26824
rect 27722 26816 27729 26856
rect 27772 26841 27775 26874
rect 27776 26864 27779 26874
rect 27786 26854 27789 26864
rect 27786 26848 27802 26854
rect 27830 26848 27842 26854
rect 27744 26824 27748 26834
rect 27758 26826 27780 26834
rect 27758 26825 27774 26826
rect 27848 26824 27851 26874
rect 27874 26854 27996 26859
rect 27900 26839 27918 26846
rect 27855 26826 27875 26834
rect 28004 26826 28008 26894
rect 28143 26887 28150 26913
rect 28125 26835 28131 26875
rect 28125 26827 28141 26835
rect 27754 26820 27772 26824
rect 27641 26777 27646 26785
rect 27714 26768 27721 26816
rect 27754 26776 27760 26820
rect 27790 26776 27797 26824
rect 27848 26816 27856 26824
rect 27910 26816 27917 26824
rect 27830 26776 27832 26816
rect 27732 26768 27748 26775
rect 27754 26768 27758 26776
rect 27834 26768 27841 26816
rect 27849 26768 27856 26816
rect 27892 26777 27900 26816
rect 27892 26776 27908 26777
rect 27722 26705 27729 26768
rect 27848 26765 27856 26768
rect 27875 26765 27882 26776
rect 27900 26768 27908 26776
rect 27928 26768 27935 26816
rect 27937 26776 27941 26816
rect 27951 26776 27953 26824
rect 27958 26768 27965 26816
rect 27970 26778 27976 26816
rect 28004 26778 28011 26826
rect 28013 26778 28017 26816
rect 28053 26789 28069 26805
rect 27991 26768 27998 26778
rect 28092 26777 28093 26818
rect 28151 26815 28158 26979
rect 28181 26883 28188 26979
rect 28163 26835 28168 26875
rect 28173 26835 28180 26883
rect 28200 26875 28206 26883
rect 28225 26879 28226 26905
rect 28247 26885 28290 26893
rect 28237 26875 28239 26883
rect 28255 26875 28257 26877
rect 28262 26875 28265 26883
rect 28200 26865 28207 26875
rect 28200 26835 28206 26865
rect 28211 26849 28217 26865
rect 28237 26835 28253 26875
rect 28255 26835 28262 26875
rect 28264 26835 28282 26875
rect 28301 26857 28302 26979
rect 28442 26882 28449 26979
rect 28492 26976 28495 26979
rect 28568 26968 28571 26979
rect 28609 26970 28612 26979
rect 28627 26978 28713 26979
rect 28769 26978 28774 26979
rect 28662 26960 28665 26961
rect 28472 26952 28478 26960
rect 28485 26952 28499 26960
rect 28559 26952 28568 26953
rect 28628 26952 28630 26960
rect 28637 26952 28671 26960
rect 28492 26950 28495 26952
rect 28568 26950 28571 26952
rect 28478 26902 28485 26950
rect 28488 26902 28489 26942
rect 28473 26894 28482 26902
rect 28492 26894 28499 26942
rect 28510 26902 28517 26950
rect 28561 26947 28575 26950
rect 28568 26942 28575 26947
rect 28549 26902 28552 26942
rect 28504 26894 28549 26902
rect 28554 26894 28561 26942
rect 28569 26894 28575 26942
rect 28626 26902 28628 26942
rect 28630 26902 28637 26950
rect 28657 26947 28678 26950
rect 28671 26942 28678 26947
rect 28724 26942 28728 26978
rect 28645 26902 28646 26942
rect 28595 26894 28602 26902
rect 28648 26894 28655 26942
rect 28659 26902 28663 26942
rect 28671 26902 28675 26942
rect 28702 26902 28703 26942
rect 28678 26894 28685 26902
rect 28711 26894 28718 26942
rect 28757 26894 28779 26895
rect 28492 26882 28495 26894
rect 28568 26892 28575 26894
rect 28568 26882 28571 26892
rect 28432 26874 28504 26882
rect 28549 26874 28626 26882
rect 28442 26872 28449 26874
rect 28452 26856 28456 26862
rect 28181 26815 28188 26835
rect 28251 26827 28257 26835
rect 28266 26827 28270 26835
rect 28280 26827 28282 26835
rect 28151 26807 28188 26815
rect 28151 26795 28158 26807
rect 28145 26787 28158 26795
rect 28151 26781 28158 26787
rect 28067 26770 28093 26777
rect 28181 26775 28188 26807
rect 28207 26787 28242 26795
rect 27960 26767 27963 26768
rect 28004 26767 28008 26768
rect 28145 26765 28146 26767
rect 27736 26747 27772 26755
rect 27848 26753 27851 26765
rect 28145 26757 28149 26765
rect 28158 26757 28159 26775
rect 28180 26767 28200 26775
rect 28172 26765 28176 26767
rect 28181 26765 28188 26767
rect 28301 26765 28302 26841
rect 28313 26827 28315 26835
rect 28328 26827 28356 26836
rect 28340 26776 28343 26824
rect 28361 26776 28366 26824
rect 28442 26816 28449 26856
rect 28492 26841 28495 26874
rect 28496 26864 28499 26874
rect 28506 26854 28509 26864
rect 28506 26848 28522 26854
rect 28550 26848 28562 26854
rect 28464 26824 28468 26834
rect 28478 26826 28500 26834
rect 28478 26825 28494 26826
rect 28568 26824 28571 26874
rect 28594 26854 28716 26859
rect 28620 26839 28638 26846
rect 28575 26826 28595 26834
rect 28724 26826 28728 26894
rect 28863 26887 28870 26913
rect 28845 26835 28851 26875
rect 28845 26827 28861 26835
rect 28474 26820 28492 26824
rect 28308 26767 28321 26775
rect 28434 26768 28441 26816
rect 28474 26776 28480 26820
rect 28510 26776 28517 26824
rect 28568 26816 28576 26824
rect 28630 26816 28637 26824
rect 28550 26776 28552 26816
rect 28452 26768 28468 26775
rect 28474 26768 28478 26776
rect 28554 26768 28561 26816
rect 28569 26768 28576 26816
rect 28612 26777 28620 26816
rect 28612 26776 28628 26777
rect 28303 26765 28305 26767
rect 28172 26757 28180 26765
rect 28199 26757 28207 26765
rect 28225 26757 28227 26759
rect 28232 26757 28234 26765
rect 28255 26757 28257 26759
rect 28262 26757 28265 26765
rect 28301 26757 28311 26765
rect 27824 26747 27872 26753
rect 27930 26747 27941 26755
rect 27771 26737 27772 26747
rect 27796 26745 27797 26747
rect 27790 26737 27797 26745
rect 27848 26743 27851 26747
rect 27722 26697 27738 26705
rect 27712 26685 27720 26695
rect 27722 26689 27731 26697
rect 27746 26687 27748 26715
rect 27771 26689 27779 26737
rect 27796 26697 27797 26737
rect 27817 26689 27824 26737
rect 27834 26727 27850 26737
rect 27910 26735 27917 26745
rect 27960 26735 27966 26755
rect 27974 26737 27983 26745
rect 27986 26737 27993 26755
rect 27910 26719 27926 26735
rect 27888 26693 27894 26699
rect 27986 26697 27995 26737
rect 28155 26717 28159 26757
rect 28163 26717 28171 26757
rect 28173 26717 28179 26757
rect 28155 26709 28171 26717
rect 28181 26709 28188 26757
rect 28190 26717 28198 26757
rect 28200 26717 28206 26757
rect 28225 26717 28232 26757
rect 28239 26717 28253 26757
rect 28255 26717 28262 26757
rect 28264 26717 28280 26757
rect 28301 26717 28308 26757
rect 28209 26709 28210 26717
rect 28225 26709 28227 26717
rect 28255 26709 28257 26717
rect 28285 26709 28292 26717
rect 27884 26689 27888 26693
rect 27950 26685 27956 26695
rect 27986 26689 27993 26697
rect 28212 26689 28217 26697
rect 27722 26677 27730 26685
rect 27960 26677 27966 26685
rect 27722 26669 27838 26677
rect 27960 26669 27967 26677
rect 27983 26669 28001 26677
rect 28017 26669 28032 26677
rect 28185 26669 28237 26677
rect 28253 26669 28294 26677
rect 28313 26667 28321 26757
rect 28368 26713 28373 26757
rect 28366 26709 28382 26713
rect 28442 26705 28449 26768
rect 28568 26765 28576 26768
rect 28595 26765 28602 26776
rect 28620 26768 28628 26776
rect 28648 26768 28655 26816
rect 28657 26776 28661 26816
rect 28671 26776 28673 26824
rect 28678 26768 28685 26816
rect 28690 26778 28696 26816
rect 28724 26778 28731 26826
rect 28733 26778 28737 26816
rect 28773 26789 28789 26805
rect 28711 26768 28718 26778
rect 28812 26777 28813 26818
rect 28871 26815 28878 26979
rect 28901 26883 28908 26979
rect 28883 26835 28888 26875
rect 28893 26835 28900 26883
rect 28920 26875 28926 26883
rect 28945 26879 28946 26905
rect 28967 26885 29010 26893
rect 28957 26875 28959 26883
rect 28975 26875 28977 26877
rect 28982 26875 28985 26883
rect 28920 26865 28927 26875
rect 28920 26835 28926 26865
rect 28931 26849 28937 26865
rect 28957 26835 28973 26875
rect 28975 26835 28982 26875
rect 28984 26835 29002 26875
rect 29021 26857 29022 26979
rect 29162 26882 29169 26979
rect 29212 26976 29215 26979
rect 29288 26968 29291 26979
rect 29329 26970 29332 26979
rect 29347 26978 29433 26979
rect 29489 26978 29494 26979
rect 29382 26960 29385 26961
rect 29192 26952 29198 26960
rect 29205 26952 29219 26960
rect 29279 26952 29288 26953
rect 29348 26952 29350 26960
rect 29357 26952 29391 26960
rect 29212 26950 29215 26952
rect 29288 26950 29291 26952
rect 29198 26902 29205 26950
rect 29208 26902 29209 26942
rect 29193 26894 29202 26902
rect 29212 26894 29219 26942
rect 29230 26902 29237 26950
rect 29281 26947 29295 26950
rect 29288 26942 29295 26947
rect 29269 26902 29272 26942
rect 29224 26894 29269 26902
rect 29274 26894 29281 26942
rect 29289 26894 29295 26942
rect 29346 26902 29348 26942
rect 29350 26902 29357 26950
rect 29377 26947 29398 26950
rect 29391 26942 29398 26947
rect 29444 26942 29448 26978
rect 29365 26902 29366 26942
rect 29315 26894 29322 26902
rect 29368 26894 29375 26942
rect 29379 26902 29383 26942
rect 29391 26902 29395 26942
rect 29422 26902 29423 26942
rect 29398 26894 29405 26902
rect 29431 26894 29438 26942
rect 29477 26894 29499 26895
rect 29212 26882 29215 26894
rect 29288 26892 29295 26894
rect 29288 26882 29291 26892
rect 29152 26874 29224 26882
rect 29269 26874 29346 26882
rect 29162 26872 29169 26874
rect 29172 26856 29176 26862
rect 28901 26815 28908 26835
rect 28971 26827 28977 26835
rect 28986 26827 28990 26835
rect 29000 26827 29002 26835
rect 28871 26807 28908 26815
rect 28871 26795 28878 26807
rect 28865 26787 28878 26795
rect 28871 26781 28878 26787
rect 28787 26770 28813 26777
rect 28901 26775 28908 26807
rect 28927 26787 28962 26795
rect 28680 26767 28683 26768
rect 28724 26767 28728 26768
rect 28865 26765 28866 26767
rect 28456 26747 28492 26755
rect 28568 26753 28571 26765
rect 28865 26757 28869 26765
rect 28878 26757 28879 26775
rect 28900 26767 28920 26775
rect 28892 26765 28896 26767
rect 28901 26765 28908 26767
rect 29021 26765 29022 26841
rect 29033 26827 29035 26835
rect 29048 26827 29076 26836
rect 29060 26776 29063 26824
rect 29081 26776 29086 26824
rect 29162 26816 29169 26856
rect 29212 26841 29215 26874
rect 29216 26864 29219 26874
rect 29226 26854 29229 26864
rect 29226 26848 29242 26854
rect 29270 26848 29282 26854
rect 29184 26824 29188 26834
rect 29198 26826 29220 26834
rect 29198 26825 29214 26826
rect 29288 26824 29291 26874
rect 29314 26854 29436 26859
rect 29340 26839 29358 26846
rect 29295 26826 29315 26834
rect 29444 26826 29448 26894
rect 29583 26887 29590 26913
rect 29565 26835 29571 26875
rect 29565 26827 29581 26835
rect 29194 26820 29212 26824
rect 29028 26767 29041 26775
rect 29154 26768 29161 26816
rect 29194 26776 29200 26820
rect 29230 26776 29237 26824
rect 29288 26816 29296 26824
rect 29350 26816 29357 26824
rect 29270 26776 29272 26816
rect 29172 26768 29188 26775
rect 29194 26768 29198 26776
rect 29274 26768 29281 26816
rect 29289 26768 29296 26816
rect 29332 26777 29340 26816
rect 29332 26776 29348 26777
rect 29023 26765 29025 26767
rect 28892 26757 28900 26765
rect 28919 26757 28927 26765
rect 28945 26757 28947 26759
rect 28952 26757 28954 26765
rect 28975 26757 28977 26759
rect 28982 26757 28985 26765
rect 29021 26757 29031 26765
rect 28544 26747 28592 26753
rect 28650 26747 28661 26755
rect 28491 26737 28492 26747
rect 28516 26745 28517 26747
rect 28510 26737 28517 26745
rect 28568 26743 28571 26747
rect 28442 26697 28458 26705
rect 28432 26685 28440 26695
rect 28442 26689 28451 26697
rect 28466 26687 28468 26715
rect 28491 26689 28499 26737
rect 28516 26697 28517 26737
rect 28537 26689 28544 26737
rect 28554 26727 28570 26737
rect 28630 26735 28637 26745
rect 28680 26735 28686 26755
rect 28694 26737 28703 26745
rect 28706 26737 28713 26755
rect 28630 26719 28646 26735
rect 28608 26693 28614 26699
rect 28706 26697 28715 26737
rect 28875 26717 28879 26757
rect 28883 26717 28891 26757
rect 28893 26717 28899 26757
rect 28875 26709 28891 26717
rect 28901 26709 28908 26757
rect 28910 26717 28918 26757
rect 28920 26717 28926 26757
rect 28945 26717 28952 26757
rect 28959 26717 28973 26757
rect 28975 26717 28982 26757
rect 28984 26717 29000 26757
rect 29021 26717 29028 26757
rect 28929 26709 28930 26717
rect 28945 26709 28947 26717
rect 28975 26709 28977 26717
rect 29005 26709 29012 26717
rect 28604 26689 28608 26693
rect 28670 26685 28676 26695
rect 28706 26689 28713 26697
rect 28932 26689 28937 26697
rect 28442 26677 28450 26685
rect 28680 26677 28686 26685
rect 28442 26669 28558 26677
rect 28680 26669 28687 26677
rect 28703 26669 28721 26677
rect 28737 26669 28752 26677
rect 28905 26669 28957 26677
rect 28973 26669 29014 26677
rect 29033 26667 29041 26757
rect 29088 26713 29093 26757
rect 29086 26709 29102 26713
rect 29162 26705 29169 26768
rect 29288 26765 29296 26768
rect 29315 26765 29322 26776
rect 29340 26768 29348 26776
rect 29368 26768 29375 26816
rect 29377 26776 29381 26816
rect 29391 26776 29393 26824
rect 29398 26768 29405 26816
rect 29410 26778 29416 26816
rect 29444 26778 29451 26826
rect 29453 26778 29457 26816
rect 29493 26789 29509 26805
rect 29431 26768 29438 26778
rect 29532 26777 29533 26818
rect 29591 26815 29598 26979
rect 29621 26883 29628 26979
rect 29603 26835 29608 26875
rect 29613 26835 29620 26883
rect 29640 26875 29646 26883
rect 29665 26879 29666 26905
rect 29687 26885 29730 26893
rect 29677 26875 29679 26883
rect 29695 26875 29697 26877
rect 29702 26875 29705 26883
rect 29640 26865 29647 26875
rect 29640 26835 29646 26865
rect 29651 26849 29657 26865
rect 29677 26835 29693 26875
rect 29695 26835 29702 26875
rect 29704 26835 29722 26875
rect 29741 26857 29742 26979
rect 29882 26882 29889 26979
rect 29932 26976 29935 26979
rect 30008 26968 30011 26979
rect 30049 26970 30052 26979
rect 30067 26978 30153 26979
rect 30209 26978 30214 26979
rect 30102 26960 30105 26961
rect 29912 26952 29918 26960
rect 29925 26952 29939 26960
rect 29999 26952 30008 26953
rect 30068 26952 30070 26960
rect 30077 26952 30111 26960
rect 29932 26950 29935 26952
rect 30008 26950 30011 26952
rect 29918 26902 29925 26950
rect 29928 26902 29929 26942
rect 29913 26894 29922 26902
rect 29932 26894 29939 26942
rect 29950 26902 29957 26950
rect 30001 26947 30015 26950
rect 30008 26942 30015 26947
rect 29989 26902 29992 26942
rect 29944 26894 29989 26902
rect 29994 26894 30001 26942
rect 30009 26894 30015 26942
rect 30066 26902 30068 26942
rect 30070 26902 30077 26950
rect 30097 26947 30118 26950
rect 30111 26942 30118 26947
rect 30164 26942 30168 26978
rect 30085 26902 30086 26942
rect 30035 26894 30042 26902
rect 30088 26894 30095 26942
rect 30099 26902 30103 26942
rect 30111 26902 30115 26942
rect 30142 26902 30143 26942
rect 30118 26894 30125 26902
rect 30151 26894 30158 26942
rect 30197 26894 30219 26895
rect 29932 26882 29935 26894
rect 30008 26892 30015 26894
rect 30008 26882 30011 26892
rect 29872 26874 29944 26882
rect 29989 26874 30066 26882
rect 29882 26872 29889 26874
rect 29892 26856 29896 26862
rect 29621 26815 29628 26835
rect 29691 26827 29697 26835
rect 29706 26827 29710 26835
rect 29720 26827 29722 26835
rect 29591 26807 29628 26815
rect 29591 26795 29598 26807
rect 29585 26787 29598 26795
rect 29591 26781 29598 26787
rect 29507 26770 29533 26777
rect 29621 26775 29628 26807
rect 29647 26787 29682 26795
rect 29400 26767 29403 26768
rect 29444 26767 29448 26768
rect 29585 26765 29586 26767
rect 29176 26747 29212 26755
rect 29288 26753 29291 26765
rect 29585 26757 29589 26765
rect 29598 26757 29599 26775
rect 29620 26767 29640 26775
rect 29612 26765 29616 26767
rect 29621 26765 29628 26767
rect 29741 26765 29742 26841
rect 29753 26827 29755 26835
rect 29768 26827 29796 26836
rect 29780 26776 29783 26824
rect 29801 26776 29806 26824
rect 29882 26816 29889 26856
rect 29932 26841 29935 26874
rect 29936 26864 29939 26874
rect 29946 26854 29949 26864
rect 29946 26848 29962 26854
rect 29990 26848 30002 26854
rect 29904 26824 29908 26834
rect 29918 26826 29940 26834
rect 29918 26825 29934 26826
rect 30008 26824 30011 26874
rect 30034 26854 30156 26859
rect 30060 26839 30078 26846
rect 30015 26826 30035 26834
rect 30164 26826 30168 26894
rect 30303 26887 30310 26913
rect 30285 26835 30291 26875
rect 30285 26827 30301 26835
rect 29914 26820 29932 26824
rect 29748 26767 29761 26775
rect 29874 26768 29881 26816
rect 29914 26776 29920 26820
rect 29950 26776 29957 26824
rect 30008 26816 30016 26824
rect 30070 26816 30077 26824
rect 29990 26776 29992 26816
rect 29892 26768 29908 26775
rect 29914 26768 29918 26776
rect 29994 26768 30001 26816
rect 30009 26768 30016 26816
rect 30052 26777 30060 26816
rect 30052 26776 30068 26777
rect 29743 26765 29745 26767
rect 29612 26757 29620 26765
rect 29639 26757 29647 26765
rect 29665 26757 29667 26759
rect 29672 26757 29674 26765
rect 29695 26757 29697 26759
rect 29702 26757 29705 26765
rect 29741 26757 29751 26765
rect 29264 26747 29312 26753
rect 29370 26747 29381 26755
rect 29211 26737 29212 26747
rect 29236 26745 29237 26747
rect 29230 26737 29237 26745
rect 29288 26743 29291 26747
rect 29162 26697 29178 26705
rect 29152 26685 29160 26695
rect 29162 26689 29171 26697
rect 29186 26687 29188 26715
rect 29211 26689 29219 26737
rect 29236 26697 29237 26737
rect 29257 26689 29264 26737
rect 29274 26727 29290 26737
rect 29350 26735 29357 26745
rect 29400 26735 29406 26755
rect 29414 26737 29423 26745
rect 29426 26737 29433 26755
rect 29350 26719 29366 26735
rect 29328 26693 29334 26699
rect 29426 26697 29435 26737
rect 29595 26717 29599 26757
rect 29603 26717 29611 26757
rect 29613 26717 29619 26757
rect 29595 26709 29611 26717
rect 29621 26709 29628 26757
rect 29630 26717 29638 26757
rect 29640 26717 29646 26757
rect 29665 26717 29672 26757
rect 29679 26717 29693 26757
rect 29695 26717 29702 26757
rect 29704 26717 29720 26757
rect 29741 26717 29748 26757
rect 29649 26709 29650 26717
rect 29665 26709 29667 26717
rect 29695 26709 29697 26717
rect 29725 26709 29732 26717
rect 29324 26689 29328 26693
rect 29390 26685 29396 26695
rect 29426 26689 29433 26697
rect 29652 26689 29657 26697
rect 29162 26677 29170 26685
rect 29400 26677 29406 26685
rect 29162 26669 29278 26677
rect 29400 26669 29407 26677
rect 29423 26669 29441 26677
rect 29457 26669 29472 26677
rect 29625 26669 29677 26677
rect 29693 26669 29734 26677
rect 29753 26667 29761 26757
rect 29808 26713 29813 26757
rect 29806 26709 29822 26713
rect 29882 26705 29889 26768
rect 30008 26765 30016 26768
rect 30035 26765 30042 26776
rect 30060 26768 30068 26776
rect 30088 26768 30095 26816
rect 30097 26776 30101 26816
rect 30111 26776 30113 26824
rect 30118 26768 30125 26816
rect 30130 26778 30136 26816
rect 30164 26778 30171 26826
rect 30173 26778 30177 26816
rect 30213 26789 30229 26805
rect 30151 26768 30158 26778
rect 30252 26777 30253 26818
rect 30311 26815 30318 26979
rect 30341 26883 30348 26979
rect 30323 26835 30328 26875
rect 30333 26835 30340 26883
rect 30360 26875 30366 26883
rect 30385 26879 30386 26905
rect 30407 26885 30450 26893
rect 30397 26875 30399 26883
rect 30415 26875 30417 26877
rect 30422 26875 30425 26883
rect 30360 26865 30367 26875
rect 30360 26835 30366 26865
rect 30371 26849 30377 26865
rect 30397 26835 30413 26875
rect 30415 26835 30422 26875
rect 30424 26835 30442 26875
rect 30461 26857 30462 26979
rect 30479 26903 30484 26913
rect 30492 26903 30494 26979
rect 30489 26889 30494 26903
rect 30492 26885 30494 26889
rect 30492 26843 30499 26885
rect 30511 26849 30516 26875
rect 30341 26815 30348 26835
rect 30411 26827 30417 26835
rect 30426 26827 30430 26835
rect 30440 26827 30442 26835
rect 30311 26807 30348 26815
rect 30311 26795 30318 26807
rect 30305 26787 30318 26795
rect 30311 26781 30318 26787
rect 30227 26770 30253 26777
rect 30341 26775 30348 26807
rect 30367 26787 30402 26795
rect 30120 26767 30123 26768
rect 30164 26767 30168 26768
rect 30305 26765 30306 26767
rect 29896 26747 29932 26755
rect 30008 26753 30011 26765
rect 30305 26757 30309 26765
rect 30318 26757 30319 26775
rect 30340 26767 30360 26775
rect 30332 26765 30336 26767
rect 30341 26765 30348 26767
rect 30461 26765 30462 26841
rect 30492 26839 30500 26843
rect 30510 26839 30516 26849
rect 30521 26839 30528 26972
rect 30529 26953 30532 26963
rect 30540 26953 30542 26979
rect 30609 26964 30614 26979
rect 30539 26937 30542 26953
rect 30473 26827 30475 26835
rect 30492 26827 30499 26839
rect 30500 26827 30509 26839
rect 30511 26827 30516 26839
rect 30492 26791 30498 26827
rect 30520 26817 30528 26839
rect 30468 26767 30481 26775
rect 30463 26765 30465 26767
rect 30332 26757 30340 26765
rect 30359 26757 30367 26765
rect 30385 26757 30387 26759
rect 30392 26757 30394 26765
rect 30415 26757 30417 26759
rect 30422 26757 30425 26765
rect 30461 26757 30471 26765
rect 29984 26747 30032 26753
rect 30090 26747 30101 26755
rect 29931 26737 29932 26747
rect 29956 26745 29957 26747
rect 29950 26737 29957 26745
rect 30008 26743 30011 26747
rect 29882 26697 29898 26705
rect 29872 26685 29880 26695
rect 29882 26689 29891 26697
rect 29906 26687 29908 26715
rect 29931 26689 29939 26737
rect 29956 26697 29957 26737
rect 29977 26689 29984 26737
rect 29994 26727 30010 26737
rect 30070 26735 30077 26745
rect 30120 26735 30126 26755
rect 30134 26737 30143 26745
rect 30146 26737 30153 26755
rect 30070 26719 30086 26735
rect 30048 26693 30054 26699
rect 30146 26697 30155 26737
rect 30315 26717 30319 26757
rect 30323 26717 30331 26757
rect 30333 26717 30339 26757
rect 30315 26709 30331 26717
rect 30341 26709 30348 26757
rect 30350 26717 30358 26757
rect 30360 26717 30366 26757
rect 30385 26717 30392 26757
rect 30399 26717 30413 26757
rect 30415 26717 30422 26757
rect 30424 26717 30440 26757
rect 30461 26717 30468 26757
rect 30369 26709 30370 26717
rect 30385 26709 30387 26717
rect 30415 26709 30417 26717
rect 30445 26709 30452 26717
rect 30044 26689 30048 26693
rect 30110 26685 30116 26695
rect 30146 26689 30153 26697
rect 30372 26689 30377 26697
rect 29882 26677 29890 26685
rect 30120 26677 30126 26685
rect 29882 26669 29998 26677
rect 30120 26669 30127 26677
rect 30143 26669 30161 26677
rect 30177 26669 30192 26677
rect 30345 26669 30397 26677
rect 30413 26669 30454 26677
rect 30473 26667 30481 26757
rect 27472 26650 27480 26658
rect 27500 26650 27518 26658
rect 27532 26650 27544 26658
rect 27560 26650 27572 26658
rect 27630 26650 27636 26658
rect 27658 26650 27664 26658
rect 27690 26650 27698 26658
rect 27718 26650 27726 26658
rect 27746 26650 27754 26658
rect 27774 26650 27782 26658
rect 27785 26656 27798 26658
rect 27802 26650 27810 26658
rect 27830 26650 27838 26658
rect 27843 26656 27854 26658
rect 27858 26650 27866 26658
rect 27886 26650 27894 26658
rect 27914 26650 27922 26658
rect 27942 26650 27950 26658
rect 27970 26650 27978 26658
rect 27998 26656 28016 26658
rect 27998 26650 28006 26656
rect 28062 26650 28070 26661
rect 28090 26650 28098 26661
rect 28110 26653 28118 26661
rect 28122 26653 28130 26661
rect 28138 26653 28146 26661
rect 28150 26653 28158 26661
rect 28166 26653 28174 26661
rect 28178 26653 28186 26661
rect 28194 26653 28202 26661
rect 28206 26653 28214 26661
rect 28222 26653 28230 26661
rect 28234 26653 28242 26661
rect 28250 26653 28258 26661
rect 28262 26653 28270 26661
rect 28278 26653 28286 26661
rect 28290 26653 28298 26661
rect 28306 26653 28314 26661
rect 28318 26653 28334 26658
rect 28350 26653 28362 26658
rect 28378 26653 28390 26658
rect 28122 26652 28138 26653
rect 28150 26652 28166 26653
rect 28178 26652 28194 26653
rect 28206 26652 28222 26653
rect 28234 26652 28250 26653
rect 28262 26652 28278 26653
rect 28290 26652 28306 26653
rect 28318 26652 28326 26653
rect 27480 26642 27488 26650
rect 27516 26639 27518 26650
rect 27528 26642 27532 26650
rect 27540 26639 27542 26650
rect 27556 26642 27560 26650
rect 27564 26639 27566 26650
rect 27620 26642 27630 26650
rect 27648 26642 27658 26650
rect 27698 26642 27706 26650
rect 27726 26642 27734 26650
rect 27754 26642 27762 26650
rect 27782 26642 27790 26650
rect 27810 26642 27818 26650
rect 27838 26642 27846 26650
rect 27866 26642 27874 26650
rect 27894 26642 27902 26650
rect 27922 26642 27930 26650
rect 27950 26642 27958 26650
rect 27978 26642 27986 26650
rect 28006 26642 28014 26650
rect 28054 26645 28062 26650
rect 28082 26645 28090 26650
rect 28130 26645 28138 26652
rect 28158 26645 28166 26652
rect 28186 26645 28194 26652
rect 28214 26645 28222 26652
rect 28242 26645 28250 26652
rect 28270 26645 28278 26652
rect 28298 26645 28306 26652
rect 28346 26642 28350 26653
rect 28374 26642 28378 26653
rect 28410 26650 28418 26658
rect 28438 26650 28446 26658
rect 28466 26650 28474 26658
rect 28494 26650 28502 26658
rect 28505 26656 28518 26658
rect 28522 26650 28530 26658
rect 28550 26650 28558 26658
rect 28563 26656 28574 26658
rect 28578 26650 28586 26658
rect 28606 26650 28614 26658
rect 28634 26650 28642 26658
rect 28662 26650 28670 26658
rect 28690 26650 28698 26658
rect 28718 26656 28736 26658
rect 28718 26650 28726 26656
rect 28782 26650 28790 26661
rect 28810 26650 28818 26661
rect 28830 26653 28838 26661
rect 28842 26653 28850 26661
rect 28858 26653 28866 26661
rect 28870 26653 28878 26661
rect 28886 26653 28894 26661
rect 28898 26653 28906 26661
rect 28914 26653 28922 26661
rect 28926 26653 28934 26661
rect 28942 26653 28950 26661
rect 28954 26653 28962 26661
rect 28970 26653 28978 26661
rect 28982 26653 28990 26661
rect 28998 26653 29006 26661
rect 29010 26653 29018 26661
rect 29026 26653 29034 26661
rect 29038 26653 29054 26658
rect 29070 26653 29082 26658
rect 29098 26653 29110 26658
rect 28842 26652 28858 26653
rect 28870 26652 28886 26653
rect 28898 26652 28914 26653
rect 28926 26652 28942 26653
rect 28954 26652 28970 26653
rect 28982 26652 28998 26653
rect 29010 26652 29026 26653
rect 29038 26652 29046 26653
rect 28418 26642 28426 26650
rect 28446 26642 28454 26650
rect 28474 26642 28482 26650
rect 28502 26642 28510 26650
rect 28530 26642 28538 26650
rect 28558 26642 28566 26650
rect 28586 26642 28594 26650
rect 28614 26642 28622 26650
rect 28642 26642 28650 26650
rect 28670 26642 28678 26650
rect 28698 26642 28706 26650
rect 28726 26642 28734 26650
rect 28774 26645 28782 26650
rect 28802 26645 28810 26650
rect 28850 26645 28858 26652
rect 28878 26645 28886 26652
rect 28906 26645 28914 26652
rect 28934 26645 28942 26652
rect 28962 26645 28970 26652
rect 28990 26645 28998 26652
rect 29018 26645 29026 26652
rect 29066 26642 29070 26653
rect 29094 26642 29098 26653
rect 29130 26650 29138 26658
rect 29158 26650 29166 26658
rect 29186 26650 29194 26658
rect 29214 26650 29222 26658
rect 29225 26656 29238 26658
rect 29242 26650 29250 26658
rect 29270 26650 29278 26658
rect 29283 26656 29294 26658
rect 29298 26650 29306 26658
rect 29326 26650 29334 26658
rect 29354 26650 29362 26658
rect 29382 26650 29390 26658
rect 29410 26650 29418 26658
rect 29438 26656 29456 26658
rect 29438 26650 29446 26656
rect 29502 26650 29510 26661
rect 29530 26650 29538 26661
rect 29550 26653 29558 26661
rect 29562 26653 29570 26661
rect 29578 26653 29586 26661
rect 29590 26653 29598 26661
rect 29606 26653 29614 26661
rect 29618 26653 29626 26661
rect 29634 26653 29642 26661
rect 29646 26653 29654 26661
rect 29662 26653 29670 26661
rect 29674 26653 29682 26661
rect 29690 26653 29698 26661
rect 29702 26653 29710 26661
rect 29718 26653 29726 26661
rect 29730 26653 29738 26661
rect 29746 26653 29754 26661
rect 29758 26653 29774 26658
rect 29790 26653 29802 26658
rect 29818 26653 29830 26658
rect 29562 26652 29578 26653
rect 29590 26652 29606 26653
rect 29618 26652 29634 26653
rect 29646 26652 29662 26653
rect 29674 26652 29690 26653
rect 29702 26652 29718 26653
rect 29730 26652 29746 26653
rect 29758 26652 29766 26653
rect 29138 26642 29146 26650
rect 29166 26642 29174 26650
rect 29194 26642 29202 26650
rect 29222 26642 29230 26650
rect 29250 26642 29258 26650
rect 29278 26642 29286 26650
rect 29306 26642 29314 26650
rect 29334 26642 29342 26650
rect 29362 26642 29370 26650
rect 29390 26642 29398 26650
rect 29418 26642 29426 26650
rect 29446 26642 29454 26650
rect 29494 26645 29502 26650
rect 29522 26645 29530 26650
rect 29570 26645 29578 26652
rect 29598 26645 29606 26652
rect 29626 26645 29634 26652
rect 29654 26645 29662 26652
rect 29682 26645 29690 26652
rect 29710 26645 29718 26652
rect 29738 26645 29746 26652
rect 29786 26642 29790 26653
rect 29814 26642 29818 26653
rect 29850 26650 29858 26658
rect 29878 26650 29886 26658
rect 29906 26650 29914 26658
rect 29934 26650 29942 26658
rect 29945 26656 29958 26658
rect 29962 26650 29970 26658
rect 29990 26650 29998 26658
rect 30003 26656 30014 26658
rect 30018 26650 30026 26658
rect 30046 26650 30054 26658
rect 30074 26650 30082 26658
rect 30102 26650 30110 26658
rect 30130 26650 30138 26658
rect 30158 26656 30176 26658
rect 30158 26650 30166 26656
rect 30222 26650 30230 26661
rect 30250 26650 30258 26661
rect 30270 26653 30278 26661
rect 30282 26653 30290 26661
rect 30298 26653 30306 26661
rect 30310 26653 30318 26661
rect 30326 26653 30334 26661
rect 30338 26653 30346 26661
rect 30354 26653 30362 26661
rect 30366 26653 30374 26661
rect 30382 26653 30390 26661
rect 30394 26653 30402 26661
rect 30410 26653 30418 26661
rect 30422 26653 30430 26661
rect 30438 26653 30446 26661
rect 30450 26653 30458 26661
rect 30466 26653 30474 26661
rect 30478 26653 30490 26658
rect 30492 26653 30494 26791
rect 30521 26787 30528 26817
rect 30520 26783 30528 26787
rect 30520 26767 30523 26783
rect 30520 26709 30526 26767
rect 30540 26658 30542 26937
rect 30599 26903 30604 26913
rect 30612 26903 30614 26964
rect 30628 26945 30631 26979
rect 30636 26969 30638 26979
rect 30636 26945 30640 26969
rect 30555 26895 30557 26899
rect 30565 26881 30567 26895
rect 30609 26889 30614 26903
rect 30547 26791 30551 26827
rect 30569 26791 30573 26849
rect 30612 26841 30614 26889
rect 30628 26851 30631 26929
rect 30625 26841 30631 26851
rect 30636 26891 30638 26945
rect 30641 26891 30645 26979
rect 30636 26841 30645 26891
rect 30655 26841 30658 26979
rect 30586 26831 30590 26839
rect 30612 26831 30621 26841
rect 30635 26831 30648 26841
rect 30660 26831 30662 26979
rect 30704 26978 30710 26979
rect 30697 26841 30700 26851
rect 30708 26841 30710 26978
rect 30743 26903 30748 26913
rect 30756 26903 30758 26979
rect 30753 26889 30758 26903
rect 30756 26841 30758 26889
rect 30772 26851 30775 26970
rect 30769 26841 30775 26851
rect 30780 26891 30782 26979
rect 30785 26891 30789 26979
rect 30780 26841 30789 26891
rect 30799 26841 30802 26979
rect 30676 26833 30680 26841
rect 30704 26833 30710 26841
rect 30730 26833 30734 26841
rect 30756 26833 30765 26841
rect 30779 26833 30792 26841
rect 30804 26833 30806 26979
rect 30848 26978 30854 26979
rect 30841 26841 30844 26851
rect 30852 26841 30854 26978
rect 30887 26903 30892 26913
rect 30900 26903 30902 26979
rect 30897 26889 30902 26903
rect 30900 26841 30902 26889
rect 30916 26851 30919 26970
rect 30913 26841 30919 26851
rect 30924 26891 30926 26979
rect 30929 26891 30933 26979
rect 30924 26841 30933 26891
rect 30943 26841 30946 26979
rect 30820 26833 30824 26841
rect 30848 26833 30854 26841
rect 30874 26833 30878 26841
rect 30900 26833 30909 26841
rect 30923 26833 30936 26841
rect 30948 26833 30950 26979
rect 30992 26978 30998 26979
rect 30985 26841 30988 26851
rect 30996 26841 30998 26978
rect 31031 26903 31036 26913
rect 31044 26903 31046 26979
rect 31041 26889 31046 26903
rect 31044 26841 31046 26889
rect 31060 26851 31063 26970
rect 31057 26841 31063 26851
rect 31068 26891 31070 26979
rect 31073 26891 31077 26979
rect 31068 26841 31077 26891
rect 31087 26841 31090 26979
rect 30964 26833 30968 26841
rect 30992 26833 30998 26841
rect 31018 26833 31022 26841
rect 31044 26833 31053 26841
rect 31067 26833 31080 26841
rect 31092 26833 31094 26979
rect 31136 26978 31142 26979
rect 31129 26841 31132 26851
rect 31140 26841 31142 26978
rect 31108 26833 31112 26841
rect 31136 26833 31142 26841
rect 31162 26833 31166 26841
rect 30574 26791 30585 26831
rect 30587 26791 30590 26831
rect 30610 26793 30621 26831
rect 30623 26793 30626 26831
rect 30628 26793 30639 26831
rect 30641 26793 30648 26831
rect 30650 26793 30653 26831
rect 30569 26783 30572 26791
rect 30596 26667 30600 26791
rect 30506 26653 30518 26658
rect 30534 26653 30546 26658
rect 30282 26652 30298 26653
rect 30310 26652 30326 26653
rect 30338 26652 30354 26653
rect 30366 26652 30382 26653
rect 30394 26652 30410 26653
rect 30422 26652 30438 26653
rect 30450 26652 30466 26653
rect 30478 26652 30486 26653
rect 29858 26642 29866 26650
rect 29886 26642 29894 26650
rect 29914 26642 29922 26650
rect 29942 26642 29950 26650
rect 29970 26642 29978 26650
rect 29998 26642 30006 26650
rect 30026 26642 30034 26650
rect 30054 26642 30062 26650
rect 30082 26642 30090 26650
rect 30110 26642 30118 26650
rect 30138 26642 30146 26650
rect 30166 26642 30174 26650
rect 30214 26645 30222 26650
rect 30242 26645 30250 26650
rect 30290 26645 30298 26652
rect 30318 26645 30326 26652
rect 30346 26645 30354 26652
rect 30374 26645 30382 26652
rect 30402 26645 30410 26652
rect 30430 26645 30438 26652
rect 30458 26645 30466 26652
rect 30490 26642 30494 26653
rect 30518 26642 30522 26653
rect 27696 26639 27732 26642
rect 28058 26639 28092 26640
rect -19052 26634 -15710 26639
rect -15670 26634 -10166 26639
rect -10126 26634 9346 26639
rect 9386 26634 14770 26639
rect 14810 26634 17794 26639
rect 17834 26634 22714 26639
rect 22754 26634 26122 26639
rect 26162 26634 26746 26639
rect 26786 26634 28092 26639
rect 28122 26639 28156 26641
rect 28416 26639 28452 26642
rect 28778 26639 28812 26640
rect 28122 26634 28812 26639
rect 28842 26639 28876 26641
rect 29136 26639 29172 26642
rect 29498 26639 29532 26640
rect 28842 26634 29532 26639
rect 29562 26639 29596 26641
rect 29856 26639 29892 26642
rect 30218 26639 30252 26640
rect 29562 26634 30252 26639
rect 30282 26639 30316 26641
rect 30492 26639 30494 26642
rect 30540 26639 30542 26653
rect 30546 26642 30550 26653
rect 30566 26650 30574 26658
rect 30594 26650 30608 26658
rect 30574 26642 30582 26650
rect 30608 26642 30610 26650
rect 30612 26639 30614 26793
rect 30628 26785 30635 26793
rect 30636 26658 30638 26793
rect 30655 26785 30662 26831
rect 30664 26793 30666 26831
rect 30660 26658 30662 26785
rect 30686 26667 30690 26833
rect 30691 26793 30702 26833
rect 30704 26793 30711 26833
rect 30713 26793 30716 26833
rect 30718 26793 30729 26833
rect 30731 26793 30734 26833
rect 30754 26793 30765 26833
rect 30767 26793 30770 26833
rect 30772 26793 30783 26833
rect 30785 26793 30792 26833
rect 30794 26793 30797 26833
rect 30624 26650 30638 26658
rect 30652 26650 30664 26658
rect 30684 26650 30692 26658
rect 30622 26642 30624 26650
rect 30636 26639 30638 26650
rect 30650 26642 30652 26650
rect 30660 26639 30662 26650
rect 30664 26642 30666 26650
rect 30692 26642 30700 26650
rect 30708 26639 30710 26793
rect 30711 26785 30716 26793
rect 30740 26667 30744 26793
rect 30712 26650 30720 26658
rect 30740 26650 30752 26658
rect 30756 26650 30758 26793
rect 30772 26785 30779 26793
rect 30780 26658 30782 26793
rect 30799 26785 30806 26833
rect 30808 26793 30810 26833
rect 30804 26658 30806 26785
rect 30830 26667 30834 26833
rect 30835 26793 30846 26833
rect 30848 26793 30855 26833
rect 30857 26793 30860 26833
rect 30862 26793 30873 26833
rect 30875 26793 30878 26833
rect 30898 26793 30909 26833
rect 30911 26793 30914 26833
rect 30916 26793 30927 26833
rect 30929 26793 30936 26833
rect 30938 26793 30941 26833
rect 30768 26650 30782 26658
rect 30796 26650 30808 26658
rect 30828 26650 30836 26658
rect 30720 26642 30728 26650
rect 30752 26642 30758 26650
rect 30756 26639 30758 26642
rect 30780 26642 30784 26650
rect 30780 26639 30782 26642
rect 30804 26639 30806 26650
rect 30808 26642 30812 26650
rect 30836 26642 30844 26650
rect 30852 26639 30854 26793
rect 30855 26785 30860 26793
rect 30884 26667 30888 26793
rect 30856 26650 30864 26658
rect 30884 26650 30896 26658
rect 30900 26650 30902 26793
rect 30916 26785 30923 26793
rect 30924 26658 30926 26793
rect 30943 26785 30950 26833
rect 30952 26793 30954 26833
rect 30948 26658 30950 26785
rect 30974 26667 30978 26833
rect 30979 26793 30990 26833
rect 30992 26793 30999 26833
rect 31001 26793 31004 26833
rect 31006 26793 31017 26833
rect 31019 26793 31022 26833
rect 31042 26793 31053 26833
rect 31055 26793 31058 26833
rect 31060 26793 31071 26833
rect 31073 26793 31080 26833
rect 31082 26793 31085 26833
rect 30912 26650 30926 26658
rect 30940 26650 30952 26658
rect 30972 26650 30980 26658
rect 30864 26642 30872 26650
rect 30896 26642 30902 26650
rect 30900 26639 30902 26642
rect 30924 26642 30928 26650
rect 30924 26639 30926 26642
rect 30948 26639 30950 26650
rect 30952 26642 30956 26650
rect 30980 26642 30988 26650
rect 30996 26639 30998 26793
rect 30999 26785 31004 26793
rect 31028 26667 31032 26793
rect 31000 26650 31008 26658
rect 31028 26650 31040 26658
rect 31044 26650 31046 26793
rect 31060 26785 31067 26793
rect 31068 26658 31070 26793
rect 31087 26785 31094 26833
rect 31096 26793 31098 26833
rect 31092 26658 31094 26785
rect 31118 26667 31122 26833
rect 31123 26793 31134 26833
rect 31136 26793 31143 26833
rect 31145 26793 31148 26833
rect 31150 26793 31161 26833
rect 31163 26793 31166 26833
rect 31056 26650 31070 26658
rect 31084 26650 31096 26658
rect 31116 26650 31124 26658
rect 31008 26642 31016 26650
rect 31040 26642 31046 26650
rect 31044 26639 31046 26642
rect 31068 26642 31072 26650
rect 31068 26639 31070 26642
rect 31092 26639 31094 26650
rect 31096 26642 31100 26650
rect 31124 26642 31132 26650
rect 31140 26639 31142 26793
rect 31143 26785 31148 26793
rect 31172 26667 31176 26793
rect 31144 26650 31152 26658
rect 31172 26650 31186 26658
rect 31188 26650 31190 26979
rect 31206 26970 31207 26974
rect 31191 26916 31197 26964
rect 31217 26916 31219 26964
rect 31236 26658 31238 26979
rect 31267 26916 31279 26956
rect 31342 26908 31349 26956
rect 31418 26882 31425 26979
rect 31468 26976 31471 26979
rect 31544 26968 31547 26979
rect 31585 26970 31588 26979
rect 31603 26978 31689 26979
rect 31638 26960 31641 26961
rect 31448 26952 31454 26960
rect 31461 26952 31475 26960
rect 31535 26952 31544 26953
rect 31604 26952 31606 26960
rect 31613 26952 31647 26960
rect 31468 26950 31471 26952
rect 31544 26950 31547 26952
rect 31454 26902 31461 26950
rect 31464 26902 31465 26942
rect 31449 26894 31458 26902
rect 31468 26894 31475 26942
rect 31486 26902 31493 26950
rect 31537 26947 31551 26950
rect 31544 26942 31551 26947
rect 31525 26902 31528 26942
rect 31480 26894 31525 26902
rect 31530 26894 31537 26942
rect 31545 26894 31551 26942
rect 31602 26902 31604 26942
rect 31606 26902 31613 26950
rect 31633 26947 31654 26950
rect 31647 26942 31654 26947
rect 31700 26942 31704 26978
rect 31621 26902 31622 26942
rect 31571 26894 31578 26902
rect 31624 26894 31631 26942
rect 31635 26902 31639 26942
rect 31647 26902 31651 26942
rect 31678 26902 31679 26942
rect 31654 26894 31661 26902
rect 31687 26894 31694 26942
rect 31468 26882 31471 26894
rect 31544 26892 31551 26894
rect 31544 26882 31547 26892
rect 31408 26874 31480 26882
rect 31525 26874 31602 26882
rect 31418 26872 31425 26874
rect 31428 26856 31432 26862
rect 31418 26816 31425 26856
rect 31468 26841 31471 26874
rect 31472 26864 31475 26874
rect 31482 26854 31485 26864
rect 31482 26848 31498 26854
rect 31526 26848 31538 26854
rect 31440 26824 31444 26834
rect 31454 26826 31476 26834
rect 31454 26825 31470 26826
rect 31544 26824 31547 26874
rect 31570 26854 31692 26859
rect 31596 26839 31614 26846
rect 31551 26826 31571 26834
rect 31700 26826 31704 26894
rect 31450 26820 31468 26824
rect 31410 26768 31417 26816
rect 31450 26776 31456 26820
rect 31486 26776 31493 26824
rect 31544 26816 31552 26824
rect 31606 26816 31613 26824
rect 31526 26776 31528 26816
rect 31428 26768 31444 26775
rect 31450 26768 31454 26776
rect 31530 26768 31537 26816
rect 31545 26768 31552 26816
rect 31588 26777 31596 26816
rect 31588 26776 31604 26777
rect 31418 26705 31425 26768
rect 31544 26765 31552 26768
rect 31571 26765 31578 26776
rect 31596 26768 31604 26776
rect 31624 26768 31631 26816
rect 31633 26776 31637 26816
rect 31647 26776 31649 26824
rect 31654 26768 31661 26816
rect 31666 26778 31672 26816
rect 31700 26778 31707 26826
rect 31709 26778 31713 26816
rect 31687 26768 31694 26778
rect 31770 26771 31774 26818
rect 31843 26815 31846 26841
rect 31854 26815 31860 26979
rect 31884 26824 31891 26979
rect 31960 26932 31967 26979
rect 32020 26948 32029 26979
rect 32068 26947 32071 26979
rect 32076 26971 32078 26979
rect 32076 26947 32080 26971
rect 32006 26934 32008 26939
rect 32018 26934 32020 26939
rect 32020 26929 32028 26934
rect 32030 26924 32038 26929
rect 32049 26921 32054 26934
rect 31788 26783 31789 26813
rect 31835 26805 31837 26815
rect 31854 26805 31861 26815
rect 31874 26805 31881 26824
rect 31897 26823 31909 26824
rect 31896 26807 31909 26823
rect 31845 26789 31847 26805
rect 31864 26789 31881 26805
rect 31770 26770 31787 26771
rect 31656 26767 31659 26768
rect 31700 26767 31704 26768
rect 31432 26747 31468 26755
rect 31544 26753 31547 26765
rect 31854 26763 31860 26789
rect 31866 26776 31881 26789
rect 31901 26776 31908 26807
rect 31933 26789 31937 26837
rect 31960 26826 31967 26916
rect 32059 26911 32063 26913
rect 32068 26911 32071 26931
rect 32027 26883 32033 26909
rect 32049 26908 32054 26911
rect 32063 26903 32071 26911
rect 32068 26851 32071 26903
rect 31942 26789 31949 26816
rect 31951 26781 31958 26816
rect 31520 26747 31568 26753
rect 31626 26747 31637 26755
rect 31467 26737 31468 26747
rect 31492 26745 31493 26747
rect 31486 26737 31493 26745
rect 31544 26743 31547 26747
rect 31418 26697 31434 26705
rect 31408 26685 31416 26695
rect 31418 26689 31427 26697
rect 31442 26687 31444 26715
rect 31467 26689 31475 26737
rect 31492 26697 31493 26737
rect 31513 26689 31520 26737
rect 31530 26727 31546 26737
rect 31606 26735 31613 26745
rect 31656 26735 31662 26755
rect 31670 26737 31679 26745
rect 31682 26737 31689 26755
rect 31734 26747 31751 26755
rect 31761 26747 31774 26755
rect 31772 26746 31774 26747
rect 31606 26719 31622 26735
rect 31584 26693 31590 26699
rect 31682 26697 31691 26737
rect 31744 26697 31755 26737
rect 31773 26697 31774 26746
rect 31827 26737 31833 26755
rect 31839 26747 31847 26759
rect 31884 26755 31891 26776
rect 31960 26768 31968 26826
rect 31969 26789 31976 26816
rect 31978 26781 31985 26816
rect 31987 26789 31995 26826
rect 32008 26819 32013 26847
rect 32065 26841 32071 26851
rect 32076 26891 32078 26947
rect 32081 26891 32085 26979
rect 32095 26891 32098 26979
rect 32076 26841 32085 26891
rect 32100 26885 32102 26979
rect 32144 26978 32150 26979
rect 32095 26841 32098 26875
rect 32100 26861 32109 26885
rect 32026 26829 32030 26837
rect 32009 26789 32013 26819
rect 32014 26789 32025 26829
rect 32027 26789 32030 26829
rect 32050 26793 32052 26829
rect 32054 26793 32061 26841
rect 32075 26829 32088 26841
rect 32100 26829 32102 26861
rect 32137 26841 32140 26851
rect 32148 26841 32150 26978
rect 32116 26833 32120 26841
rect 32144 26833 32150 26841
rect 32170 26833 32174 26841
rect 32063 26793 32066 26829
rect 32068 26793 32079 26829
rect 32081 26793 32088 26829
rect 32090 26793 32093 26829
rect 32009 26781 32012 26789
rect 31850 26751 31874 26755
rect 31881 26751 31892 26755
rect 31850 26747 31863 26751
rect 31839 26745 31849 26747
rect 31854 26745 31860 26747
rect 31884 26745 31891 26751
rect 31902 26745 31909 26747
rect 31843 26742 31854 26745
rect 31861 26742 31868 26745
rect 31843 26737 31852 26742
rect 31873 26737 31882 26745
rect 31901 26737 31909 26745
rect 31915 26737 31919 26751
rect 31820 26697 31823 26737
rect 31825 26697 31832 26737
rect 31836 26697 31840 26737
rect 31843 26697 31850 26737
rect 31855 26697 31862 26737
rect 31866 26697 31871 26737
rect 31874 26697 31881 26737
rect 31883 26697 31892 26737
rect 31893 26697 31899 26737
rect 31901 26697 31908 26737
rect 31580 26689 31584 26693
rect 31646 26685 31652 26695
rect 31682 26689 31689 26697
rect 31820 26689 31840 26697
rect 31854 26689 31861 26697
rect 31883 26689 31891 26697
rect 31912 26689 31919 26737
rect 31960 26689 31968 26747
rect 31418 26677 31426 26685
rect 31656 26677 31662 26685
rect 31886 26677 31889 26689
rect 31418 26669 31534 26677
rect 31656 26669 31663 26677
rect 31679 26669 31697 26677
rect 31713 26669 31728 26677
rect 31886 26669 31893 26677
rect 31909 26669 31955 26677
rect 31960 26669 31965 26689
rect 32036 26667 32040 26789
rect 32068 26785 32075 26793
rect 31202 26650 31214 26658
rect 31230 26650 31242 26658
rect 31262 26650 31270 26658
rect 31326 26650 31334 26658
rect 31354 26650 31362 26658
rect 31386 26650 31394 26658
rect 31414 26650 31422 26658
rect 31442 26650 31450 26658
rect 31470 26650 31478 26658
rect 31481 26656 31494 26658
rect 31498 26650 31506 26658
rect 31526 26650 31534 26658
rect 31539 26656 31550 26658
rect 31554 26650 31562 26658
rect 31582 26650 31590 26658
rect 31610 26650 31618 26658
rect 31638 26650 31646 26658
rect 31666 26650 31674 26658
rect 31694 26656 31712 26658
rect 31694 26650 31702 26656
rect 31750 26650 31756 26661
rect 31778 26650 31784 26661
rect 31820 26653 31828 26661
rect 31832 26653 31840 26661
rect 31848 26653 31856 26661
rect 31860 26653 31868 26661
rect 31876 26653 31884 26661
rect 31888 26653 31896 26661
rect 31904 26653 31912 26661
rect 32076 26658 32078 26793
rect 32095 26785 32102 26829
rect 32104 26793 32106 26829
rect 32100 26658 32102 26785
rect 32126 26667 32130 26833
rect 32131 26793 32142 26833
rect 32144 26793 32151 26833
rect 32153 26793 32156 26833
rect 32158 26793 32169 26833
rect 32171 26793 32174 26833
rect 31934 26653 31944 26658
rect 31950 26653 31960 26658
rect 31962 26653 31972 26658
rect 31978 26653 31988 26658
rect 31832 26652 31848 26653
rect 31860 26652 31876 26653
rect 31888 26652 31904 26653
rect 31916 26652 31924 26653
rect 31934 26652 31950 26653
rect 31962 26652 31978 26653
rect 31990 26652 32000 26658
rect 31152 26642 31160 26650
rect 31186 26642 31190 26650
rect 31200 26642 31202 26650
rect 31214 26642 31216 26650
rect 31228 26642 31230 26650
rect 31188 26639 31190 26642
rect 31236 26639 31238 26650
rect 31242 26642 31244 26650
rect 31270 26642 31278 26650
rect 31318 26642 31326 26650
rect 31346 26642 31354 26650
rect 31394 26642 31402 26650
rect 31422 26642 31430 26650
rect 31450 26642 31458 26650
rect 31478 26642 31486 26650
rect 31506 26642 31514 26650
rect 31534 26642 31542 26650
rect 31562 26642 31570 26650
rect 31590 26642 31598 26650
rect 31618 26642 31626 26650
rect 31646 26642 31654 26650
rect 31674 26642 31682 26650
rect 31702 26642 31710 26650
rect 31756 26645 31766 26650
rect 31784 26645 31794 26650
rect 31840 26645 31848 26652
rect 31868 26645 31876 26652
rect 31896 26645 31904 26652
rect 31944 26642 31950 26652
rect 31972 26642 31978 26652
rect 32010 26650 32018 26658
rect 32038 26650 32048 26658
rect 32066 26650 32078 26658
rect 32094 26650 32104 26658
rect 32124 26650 32132 26658
rect 32018 26642 32026 26650
rect 32048 26642 32054 26650
rect 32076 26642 32082 26650
rect 31392 26639 31428 26642
rect 31778 26639 31812 26641
rect 32076 26639 32078 26642
rect 32100 26639 32102 26650
rect 32104 26642 32110 26650
rect 32132 26642 32140 26650
rect 32148 26639 32150 26793
rect 32151 26785 32156 26793
rect 32180 26667 32184 26793
rect 32152 26650 32160 26658
rect 32160 26642 32168 26650
rect 30282 26634 31738 26639
rect 31778 26634 32194 26639
rect -17916 26616 -17914 26634
rect -17868 26616 -17866 26634
rect -17820 26616 -17818 26634
rect -17772 26616 -17770 26634
rect -17652 26616 -17650 26634
rect -17532 26616 -17530 26634
rect -17436 26616 -17434 26634
rect -17412 26616 -17410 26634
rect -17364 26616 -17362 26634
rect -17316 26616 -17314 26634
rect -17220 26616 -17218 26634
rect -17196 26616 -17194 26634
rect -17124 26616 -17122 26634
rect -17028 26616 -17026 26634
rect -16980 26616 -16978 26634
rect -16884 26616 -16882 26634
rect -16860 26616 -16858 26634
rect -16812 26616 -16810 26634
rect -16788 26616 -16786 26634
rect -16764 26616 -16762 26634
rect -16716 26616 -16714 26634
rect -16692 26616 -16690 26634
rect -16668 26616 -16666 26634
rect -16596 26616 -16594 26634
rect -16500 26616 -16498 26634
rect -16404 26616 -16402 26634
rect -16380 26616 -16378 26634
rect -16332 26616 -16330 26634
rect -16308 26616 -16306 26634
rect -16284 26616 -16282 26634
rect -16236 26616 -16234 26634
rect -16212 26616 -16210 26634
rect -16188 26616 -16186 26634
rect -15420 26616 -15418 26634
rect -15396 26616 -15394 26634
rect -15372 26616 -15370 26634
rect -15300 26616 -15298 26634
rect -15084 26616 -15082 26634
rect -15036 26616 -15034 26634
rect -14940 26616 -14938 26634
rect -14916 26616 -14914 26634
rect -14868 26616 -14866 26634
rect -14820 26616 -14818 26634
rect -14724 26616 -14722 26634
rect -14700 26616 -14698 26634
rect -14652 26616 -14650 26634
rect -14604 26616 -14602 26634
rect -14508 26616 -14506 26634
rect -14484 26616 -14482 26634
rect -14436 26616 -14434 26634
rect -14388 26616 -14386 26634
rect -14268 26616 -14266 26634
rect -14172 26616 -14170 26634
rect -14076 26616 -14074 26634
rect -14028 26616 -14026 26634
rect -13980 26616 -13978 26634
rect -13956 26616 -13954 26634
rect -13932 26616 -13930 26634
rect -13860 26616 -13858 26634
rect -13764 26616 -13762 26634
rect -13716 26616 -13714 26634
rect -13644 26616 -13642 26634
rect -13596 26616 -13594 26634
rect -13500 26616 -13498 26634
rect -13404 26616 -13402 26634
rect -13356 26616 -13354 26634
rect -13284 26616 -13282 26634
rect -12828 26616 -12826 26634
rect -12780 26616 -12778 26634
rect -12684 26616 -12682 26634
rect -12660 26616 -12658 26634
rect -12612 26616 -12610 26634
rect -12588 26616 -12586 26634
rect -12564 26616 -12562 26634
rect -12492 26616 -12490 26634
rect -12396 26616 -12394 26634
rect -12348 26616 -12346 26634
rect -12276 26616 -12274 26634
rect -12252 26616 -12250 26634
rect -12228 26616 -12226 26634
rect -12156 26616 -12154 26634
rect -12060 26616 -12058 26634
rect -12012 26616 -12010 26634
rect -11916 26616 -11914 26634
rect -11892 26616 -11890 26634
rect -11844 26616 -11842 26634
rect -11796 26616 -11794 26634
rect -11676 26616 -11674 26634
rect -11580 26616 -11578 26634
rect -11556 26616 -11554 26634
rect -11484 26616 -11482 26634
rect -11460 26616 -11458 26634
rect -11436 26616 -11434 26634
rect -11388 26616 -11386 26634
rect -11364 26616 -11362 26634
rect -11340 26616 -11338 26634
rect -11268 26616 -11266 26634
rect -11172 26616 -11170 26634
rect -11124 26616 -11122 26634
rect -11076 26616 -11074 26634
rect -11028 26616 -11026 26634
rect -10932 26616 -10930 26634
rect -10836 26616 -10834 26634
rect -10788 26616 -10786 26634
rect -10668 26616 -10666 26634
rect -9876 26616 -9874 26634
rect -9828 26616 -9826 26634
rect -9732 26616 -9730 26634
rect -9708 26616 -9706 26634
rect -9612 26616 -9610 26634
rect -9516 26616 -9514 26634
rect -9468 26616 -9466 26634
rect -9420 26616 -9418 26634
rect -9396 26616 -9394 26634
rect -9372 26616 -9370 26634
rect -9300 26616 -9298 26634
rect -9252 26616 -9250 26634
rect -9156 26616 -9154 26634
rect -9132 26616 -9130 26634
rect -9084 26616 -9082 26634
rect -9060 26616 -9058 26634
rect -9036 26616 -9034 26634
rect -8988 26616 -8986 26634
rect -8964 26616 -8962 26634
rect -8940 26616 -8938 26634
rect -8892 26616 -8890 26634
rect -8844 26616 -8842 26634
rect -8796 26616 -8794 26634
rect -8700 26616 -8698 26634
rect -8604 26616 -8602 26634
rect -8556 26616 -8554 26634
rect -8508 26616 -8506 26634
rect -8484 26616 -8482 26634
rect -8460 26616 -8458 26634
rect -8412 26616 -8410 26634
rect -8388 26616 -8386 26634
rect -8364 26616 -8362 26634
rect -8316 26616 -8314 26634
rect -8292 26616 -8290 26634
rect -8268 26616 -8266 26634
rect -8196 26616 -8194 26634
rect -8100 26616 -8098 26634
rect -8052 26616 -8050 26634
rect -7932 26616 -7930 26634
rect -7836 26616 -7834 26634
rect -7740 26616 -7738 26634
rect -7692 26616 -7690 26634
rect -7620 26616 -7618 26634
rect -7356 26616 -7354 26634
rect -7284 26616 -7282 26634
rect -7212 26616 -7210 26634
rect -7188 26616 -7186 26634
rect -7116 26616 -7114 26634
rect -7092 26616 -7090 26634
rect -7068 26616 -7066 26634
rect -6996 26616 -6994 26634
rect -6972 26616 -6970 26634
rect -6948 26616 -6946 26634
rect -6900 26616 -6898 26634
rect -6876 26616 -6874 26634
rect -6852 26616 -6850 26634
rect -6804 26616 -6802 26634
rect -6780 26616 -6778 26634
rect -6756 26616 -6754 26634
rect -6708 26616 -6706 26634
rect -6684 26616 -6682 26634
rect -6660 26616 -6658 26634
rect -6612 26616 -6610 26634
rect -6588 26616 -6586 26634
rect -6564 26616 -6562 26634
rect -6516 26616 -6514 26634
rect -6492 26616 -6490 26634
rect -6468 26616 -6466 26634
rect -6420 26616 -6418 26634
rect -6396 26616 -6394 26634
rect -6372 26616 -6370 26634
rect -6324 26616 -6322 26634
rect -6300 26616 -6298 26634
rect -6276 26616 -6274 26634
rect -6228 26616 -6226 26634
rect -6180 26616 -6178 26634
rect -6060 26616 -6058 26634
rect -5964 26616 -5962 26634
rect -5940 26616 -5938 26634
rect -5868 26616 -5866 26634
rect -5796 26616 -5794 26634
rect -5652 26616 -5650 26634
rect -5316 26616 -5314 26634
rect -5268 26616 -5266 26634
rect -5220 26616 -5218 26634
rect -5196 26616 -5194 26634
rect -5172 26616 -5170 26634
rect -5124 26616 -5122 26634
rect -5100 26616 -5098 26634
rect -5076 26616 -5074 26634
rect -5028 26616 -5026 26634
rect -4980 26616 -4978 26634
rect -4884 26616 -4882 26634
rect -4860 26616 -4858 26634
rect -4788 26616 -4786 26634
rect -4692 26616 -4690 26634
rect -4644 26616 -4642 26634
rect -4596 26616 -4594 26634
rect -4548 26616 -4546 26634
rect -4428 26616 -4426 26634
rect -4332 26616 -4330 26634
rect -4308 26616 -4306 26634
rect -4260 26616 -4258 26634
rect -4212 26616 -4210 26634
rect -4116 26616 -4114 26634
rect -4092 26616 -4090 26634
rect -4020 26616 -4018 26634
rect -3876 26616 -3874 26634
rect -3804 26616 -3802 26634
rect -3732 26616 -3730 26634
rect -3588 26616 -3586 26634
rect -3564 26616 -3562 26634
rect -3516 26616 -3514 26634
rect -3492 26616 -3490 26634
rect -3468 26616 -3466 26634
rect -3420 26616 -3418 26634
rect -3372 26616 -3370 26634
rect -3252 26616 -3250 26634
rect -3156 26616 -3154 26634
rect -3132 26616 -3130 26634
rect -3060 26616 -3058 26634
rect -3012 26616 -3010 26634
rect -2916 26616 -2914 26634
rect -2892 26616 -2890 26634
rect -2844 26616 -2842 26634
rect -2820 26616 -2818 26634
rect -2796 26616 -2794 26634
rect -2748 26616 -2746 26634
rect -2700 26616 -2698 26634
rect -2604 26616 -2602 26634
rect -2580 26616 -2578 26634
rect -2508 26616 -2506 26634
rect -2412 26616 -2410 26634
rect -2364 26616 -2362 26634
rect -2292 26616 -2290 26634
rect -2268 26616 -2266 26634
rect -2244 26616 -2242 26634
rect -2196 26616 -2194 26634
rect -2172 26616 -2170 26634
rect -2148 26616 -2146 26634
rect -2100 26616 -2098 26634
rect -2076 26616 -2074 26634
rect -2052 26616 -2050 26634
rect -1980 26616 -1978 26634
rect -1884 26616 -1882 26634
rect -1836 26616 -1834 26634
rect -1716 26616 -1714 26634
rect -1596 26616 -1594 26634
rect -1476 26616 -1474 26634
rect -1380 26616 -1378 26634
rect -1356 26616 -1354 26634
rect -1308 26616 -1306 26634
rect -1260 26616 -1258 26634
rect -1164 26616 -1162 26634
rect -1140 26616 -1138 26634
rect -1068 26616 -1066 26634
rect -852 26616 -850 26634
rect -804 26616 -802 26634
rect -756 26616 -754 26634
rect -708 26616 -706 26634
rect -612 26616 -610 26634
rect -588 26616 -586 26634
rect -540 26616 -538 26634
rect -516 26616 -514 26634
rect -492 26616 -490 26634
rect -444 26616 -442 26634
rect -396 26616 -394 26634
rect -300 26616 -298 26634
rect -276 26616 -274 26634
rect -204 26616 -202 26634
rect -108 26616 -106 26634
rect -60 26616 -58 26634
rect 12 26616 14 26634
rect 108 26616 110 26634
rect 156 26616 158 26634
rect 204 26616 206 26634
rect 228 26616 230 26634
rect 252 26616 254 26634
rect 300 26616 302 26634
rect 348 26616 350 26634
rect 468 26616 470 26634
rect 564 26616 566 26634
rect 588 26616 590 26634
rect 636 26616 638 26634
rect 660 26616 662 26634
rect 684 26616 686 26634
rect 732 26616 734 26634
rect 756 26616 758 26634
rect 780 26616 782 26634
rect 876 26616 878 26634
rect 972 26616 974 26634
rect 1020 26616 1022 26634
rect 1068 26616 1070 26634
rect 1092 26616 1094 26634
rect 1116 26616 1118 26634
rect 1164 26616 1166 26634
rect 1212 26616 1214 26634
rect 1308 26616 1310 26634
rect 1332 26616 1334 26634
rect 1380 26616 1382 26634
rect 1428 26616 1430 26634
rect 1524 26616 1526 26634
rect 1548 26616 1550 26634
rect 1596 26616 1598 26634
rect 1620 26616 1622 26634
rect 1644 26616 1646 26634
rect 1692 26616 1694 26634
rect 1716 26616 1718 26634
rect 1740 26616 1742 26634
rect 1788 26616 1790 26634
rect 1812 26616 1814 26634
rect 1836 26616 1838 26634
rect 1884 26616 1886 26634
rect 1908 26616 1910 26634
rect 1932 26616 1934 26634
rect 1980 26616 1982 26634
rect 2004 26616 2006 26634
rect 2028 26616 2030 26634
rect 2076 26616 2078 26634
rect 2100 26616 2102 26634
rect 2124 26616 2126 26634
rect 2172 26616 2174 26634
rect 2196 26616 2198 26634
rect 2220 26616 2222 26634
rect 2268 26616 2270 26634
rect 2292 26616 2294 26634
rect 2316 26616 2318 26634
rect 2364 26616 2366 26634
rect 2388 26616 2390 26634
rect 2412 26616 2414 26634
rect 2460 26616 2462 26634
rect 2484 26616 2486 26634
rect 2508 26616 2510 26634
rect 2556 26616 2558 26634
rect 2580 26616 2582 26634
rect 2604 26616 2606 26634
rect 2652 26616 2654 26634
rect 2676 26616 2678 26634
rect 2700 26616 2702 26634
rect 2748 26616 2750 26634
rect 2772 26616 2774 26634
rect 2796 26616 2798 26634
rect 2844 26616 2846 26634
rect 2868 26616 2870 26634
rect 2892 26616 2894 26634
rect 2940 26616 2942 26634
rect 3012 26616 3014 26634
rect 3108 26616 3110 26634
rect 3156 26616 3158 26634
rect 3252 26616 3254 26634
rect 3348 26616 3350 26634
rect 3396 26616 3398 26634
rect 3468 26616 3470 26634
rect 3492 26616 3494 26634
rect 3516 26616 3518 26634
rect 3588 26616 3590 26634
rect 3612 26616 3614 26634
rect 3636 26616 3638 26634
rect 3708 26616 3710 26634
rect 3732 26616 3734 26634
rect 3756 26616 3758 26634
rect 3804 26616 3806 26634
rect 3828 26616 3830 26634
rect 3852 26616 3854 26634
rect 3900 26616 3902 26634
rect 3924 26616 3926 26634
rect 3948 26616 3950 26634
rect 3996 26616 3998 26634
rect 4020 26616 4022 26634
rect 4044 26616 4046 26634
rect 4092 26616 4094 26634
rect 4116 26616 4118 26634
rect 4140 26616 4142 26634
rect 4188 26616 4190 26634
rect 4212 26616 4214 26634
rect 4236 26616 4238 26634
rect 4284 26616 4286 26634
rect 4308 26616 4310 26634
rect 4332 26616 4334 26634
rect 4380 26616 4382 26634
rect 4404 26616 4406 26634
rect 4428 26616 4430 26634
rect 4476 26616 4478 26634
rect 4500 26616 4502 26634
rect 4524 26616 4526 26634
rect 4596 26616 4598 26634
rect 4812 26616 4814 26634
rect 4860 26616 4862 26634
rect 4908 26616 4910 26634
rect 4956 26616 4958 26634
rect 4980 26616 4982 26634
rect 5004 26616 5006 26634
rect 5076 26616 5078 26634
rect 5100 26616 5102 26634
rect 5124 26616 5126 26634
rect 5172 26616 5174 26634
rect 5196 26616 5198 26634
rect 5220 26616 5222 26634
rect 5268 26616 5270 26634
rect 5292 26616 5294 26634
rect 5316 26616 5318 26634
rect 5388 26616 5390 26634
rect 5412 26616 5414 26634
rect 5436 26616 5438 26634
rect 5484 26616 5486 26634
rect 5508 26616 5510 26634
rect 5532 26616 5534 26634
rect 5580 26616 5582 26634
rect 5628 26616 5630 26634
rect 5724 26616 5726 26634
rect 5748 26616 5750 26634
rect 5796 26616 5798 26634
rect 5820 26616 5822 26634
rect 5844 26616 5846 26634
rect 5916 26616 5918 26634
rect 6132 26616 6134 26634
rect 6180 26616 6182 26634
rect 6228 26616 6230 26634
rect 6252 26616 6254 26634
rect 6276 26616 6278 26634
rect 6324 26616 6326 26634
rect 6372 26616 6374 26634
rect 6468 26616 6470 26634
rect 6492 26616 6494 26634
rect 6564 26616 6566 26634
rect 6588 26616 6590 26634
rect 6612 26616 6614 26634
rect 6660 26616 6662 26634
rect 6684 26616 6686 26634
rect 6708 26616 6710 26634
rect 6780 26616 6782 26634
rect 6804 26616 6806 26634
rect 6828 26616 6830 26634
rect 6876 26616 6878 26634
rect 6900 26616 6902 26634
rect 6924 26616 6926 26634
rect 6972 26616 6974 26634
rect 7020 26616 7022 26634
rect 7140 26616 7142 26634
rect 7236 26616 7238 26634
rect 7260 26616 7262 26634
rect 7332 26616 7334 26634
rect 7356 26616 7358 26634
rect 7380 26616 7382 26634
rect 7428 26616 7430 26634
rect 7452 26616 7454 26634
rect 7476 26616 7478 26634
rect 7524 26616 7526 26634
rect 7548 26616 7550 26634
rect 7572 26616 7574 26634
rect 7620 26616 7622 26634
rect 7644 26616 7646 26634
rect 7668 26616 7670 26634
rect 7716 26616 7718 26634
rect 7740 26616 7742 26634
rect 7764 26616 7766 26634
rect 7836 26616 7838 26634
rect 7860 26616 7862 26634
rect 7884 26616 7886 26634
rect 7932 26616 7934 26634
rect 7956 26616 7958 26634
rect 7980 26616 7982 26634
rect 8052 26616 8054 26634
rect 8148 26616 8150 26634
rect 8196 26616 8198 26634
rect 8244 26616 8246 26634
rect 8268 26616 8270 26634
rect 8292 26616 8294 26634
rect 8340 26616 8342 26634
rect 8364 26616 8366 26634
rect 8388 26616 8390 26634
rect 8436 26616 8438 26634
rect 8460 26616 8462 26634
rect 8484 26616 8486 26634
rect 8556 26616 8558 26634
rect 8580 26616 8582 26634
rect 8604 26616 8606 26634
rect 8676 26616 8678 26634
rect 8700 26616 8702 26634
rect 8724 26616 8726 26634
rect 8772 26616 8774 26634
rect 8820 26616 8822 26634
rect 8844 26616 8846 26634
rect 8868 26616 8870 26634
rect 9660 26616 9662 26634
rect 9684 26616 9686 26634
rect 9708 26616 9710 26634
rect 9756 26616 9758 26634
rect 9780 26616 9782 26634
rect 9804 26616 9806 26634
rect 9852 26616 9854 26634
rect 9876 26616 9878 26634
rect 9900 26616 9902 26634
rect 9948 26616 9950 26634
rect 9972 26616 9974 26634
rect 9996 26616 9998 26634
rect 10068 26616 10070 26634
rect 10092 26616 10094 26634
rect 10116 26616 10118 26634
rect 10164 26616 10166 26634
rect 10188 26616 10190 26634
rect 10212 26616 10214 26634
rect 10260 26616 10262 26634
rect 10284 26616 10286 26634
rect 10308 26616 10310 26634
rect 10380 26616 10382 26634
rect 10404 26616 10406 26634
rect 10428 26616 10430 26634
rect 10476 26616 10478 26634
rect 10500 26616 10502 26634
rect 10524 26616 10526 26634
rect 10572 26616 10574 26634
rect 10596 26616 10598 26634
rect 10620 26616 10622 26634
rect 10668 26616 10670 26634
rect 10692 26616 10694 26634
rect 10716 26616 10718 26634
rect 10788 26616 10790 26634
rect 10836 26616 10838 26634
rect 10956 26616 10958 26634
rect 11052 26616 11054 26634
rect 11076 26616 11078 26634
rect 11124 26616 11126 26634
rect 11172 26616 11174 26634
rect 11220 26616 11222 26634
rect 11340 26616 11342 26634
rect 11436 26616 11438 26634
rect 11532 26616 11534 26634
rect 11580 26616 11582 26634
rect 11628 26616 11630 26634
rect 11652 26616 11654 26634
rect 11676 26616 11678 26634
rect 11748 26616 11750 26634
rect 11772 26616 11774 26634
rect 11796 26616 11798 26634
rect 11844 26616 11846 26634
rect 11892 26616 11894 26634
rect 11988 26616 11990 26634
rect 12012 26616 12014 26634
rect 12084 26616 12086 26634
rect 12132 26616 12134 26634
rect 12228 26616 12230 26634
rect 12252 26616 12254 26634
rect 12300 26616 12302 26634
rect 12324 26616 12326 26634
rect 12348 26616 12350 26634
rect 12396 26616 12398 26634
rect 12420 26616 12422 26634
rect 12444 26616 12446 26634
rect 12492 26616 12494 26634
rect 12516 26616 12518 26634
rect 12540 26616 12542 26634
rect 12588 26616 12590 26634
rect 12636 26616 12638 26634
rect 12732 26616 12734 26634
rect 12756 26616 12758 26634
rect 12804 26616 12806 26634
rect 12828 26616 12830 26634
rect 12852 26616 12854 26634
rect 12900 26616 12902 26634
rect 12924 26616 12926 26634
rect 12948 26616 12950 26634
rect 13020 26616 13022 26634
rect 13044 26616 13046 26634
rect 13068 26616 13070 26634
rect 13116 26616 13118 26634
rect 13188 26616 13190 26634
rect 13284 26616 13286 26634
rect 13332 26616 13334 26634
rect 13428 26616 13430 26634
rect 13524 26616 13526 26634
rect 13572 26616 13574 26634
rect 13644 26616 13646 26634
rect 13668 26616 13670 26634
rect 13692 26616 13694 26634
rect 13764 26616 13766 26634
rect 13788 26616 13790 26634
rect 13812 26616 13814 26634
rect 13860 26616 13862 26634
rect 13884 26616 13886 26634
rect 13908 26616 13910 26634
rect 13956 26616 13958 26634
rect 14004 26616 14006 26634
rect 14100 26616 14102 26634
rect 14196 26616 14198 26634
rect 14244 26616 14246 26634
rect 14292 26616 14294 26634
rect 15132 26616 15134 26634
rect 15228 26616 15230 26634
rect 15252 26616 15254 26634
rect 15300 26616 15302 26634
rect 15324 26616 15326 26634
rect 15348 26616 15350 26634
rect 15396 26616 15398 26634
rect 15420 26616 15422 26634
rect 15444 26616 15446 26634
rect 15492 26616 15494 26634
rect 15540 26616 15542 26634
rect 15636 26616 15638 26634
rect 15660 26616 15662 26634
rect 15708 26616 15710 26634
rect 15732 26616 15734 26634
rect 15756 26616 15758 26634
rect 15804 26616 15806 26634
rect 15828 26616 15830 26634
rect 15852 26616 15854 26634
rect 15900 26616 15902 26634
rect 15924 26616 15926 26634
rect 15948 26616 15950 26634
rect 15996 26616 15998 26634
rect 16020 26616 16022 26634
rect 16044 26616 16046 26634
rect 16092 26616 16094 26634
rect 16140 26616 16142 26634
rect 16236 26616 16238 26634
rect 16260 26616 16262 26634
rect 16308 26616 16310 26634
rect 16332 26616 16334 26634
rect 16356 26616 16358 26634
rect 16404 26616 16406 26634
rect 16452 26616 16454 26634
rect 16548 26616 16550 26634
rect 16572 26616 16574 26634
rect 16620 26616 16622 26634
rect 16644 26616 16646 26634
rect 16668 26616 16670 26634
rect 16716 26616 16718 26634
rect 16740 26616 16742 26634
rect 16764 26616 16766 26634
rect 16836 26616 16838 26634
rect 16884 26616 16886 26634
rect 16980 26616 16982 26634
rect 17004 26616 17006 26634
rect 17052 26616 17054 26634
rect 17100 26616 17102 26634
rect 17196 26616 17198 26634
rect 17220 26616 17222 26634
rect 17268 26616 17270 26634
rect 17292 26616 17294 26634
rect 17316 26616 17318 26634
rect 18084 26616 18086 26634
rect 18108 26616 18110 26634
rect 18132 26616 18134 26634
rect 18180 26616 18182 26634
rect 18252 26616 18254 26634
rect 18348 26616 18350 26634
rect 18396 26616 18398 26634
rect 18492 26616 18494 26634
rect 18516 26616 18518 26634
rect 18564 26616 18566 26634
rect 18588 26616 18590 26634
rect 18612 26616 18614 26634
rect 18660 26616 18662 26634
rect 18684 26616 18686 26634
rect 18708 26616 18710 26634
rect 18756 26616 18758 26634
rect 18780 26616 18782 26634
rect 18804 26616 18806 26634
rect 18852 26616 18854 26634
rect 18876 26616 18878 26634
rect 18900 26616 18902 26634
rect 18948 26616 18950 26634
rect 18996 26616 18998 26634
rect 19020 26616 19022 26634
rect 19044 26616 19046 26634
rect 19092 26616 19094 26634
rect 19116 26616 19118 26634
rect 19140 26616 19142 26634
rect 19188 26616 19190 26634
rect 19236 26616 19238 26634
rect 19332 26616 19334 26634
rect 19428 26616 19430 26634
rect 19476 26616 19478 26634
rect 19524 26616 19526 26634
rect 19572 26616 19574 26634
rect 19596 26616 19598 26634
rect 19620 26616 19622 26634
rect 19668 26616 19670 26634
rect 19692 26616 19694 26634
rect 19716 26616 19718 26634
rect 19764 26616 19766 26634
rect 19812 26616 19814 26634
rect 19836 26616 19838 26634
rect 19860 26616 19862 26634
rect 19932 26616 19934 26634
rect 19956 26616 19958 26634
rect 19980 26616 19982 26634
rect 20028 26616 20030 26634
rect 20052 26616 20054 26634
rect 20076 26616 20078 26634
rect 20148 26616 20150 26634
rect 20172 26616 20174 26634
rect 20196 26616 20198 26634
rect 20244 26616 20246 26634
rect 20268 26616 20270 26634
rect 20292 26616 20294 26634
rect 20340 26616 20342 26634
rect 20388 26616 20390 26634
rect 20484 26616 20486 26634
rect 20508 26616 20510 26634
rect 20556 26616 20558 26634
rect 20580 26616 20582 26634
rect 20604 26616 20606 26634
rect 20700 26616 20702 26634
rect 20916 26616 20918 26634
rect 20964 26616 20966 26634
rect 21012 26616 21014 26634
rect 21060 26616 21062 26634
rect 21084 26616 21086 26634
rect 21108 26616 21110 26634
rect 21156 26616 21158 26634
rect 21204 26616 21206 26634
rect 21300 26616 21302 26634
rect 21324 26616 21326 26634
rect 21372 26616 21374 26634
rect 21420 26616 21422 26634
rect 21444 26616 21446 26634
rect 21468 26616 21470 26634
rect 21516 26616 21518 26634
rect 21540 26616 21542 26634
rect 21564 26616 21566 26634
rect 21612 26616 21614 26634
rect 21660 26616 21662 26634
rect 21684 26616 21686 26634
rect 21708 26616 21710 26634
rect 21780 26616 21782 26634
rect 21804 26616 21806 26634
rect 21828 26616 21830 26634
rect 21900 26616 21902 26634
rect 21924 26616 21926 26634
rect 21948 26616 21950 26634
rect 22020 26616 22022 26634
rect 22044 26616 22046 26634
rect 22068 26616 22070 26634
rect 22116 26616 22118 26634
rect 22164 26616 22166 26634
rect 22188 26616 22190 26634
rect 22212 26616 22214 26634
rect 23004 26616 23006 26634
rect 23052 26616 23054 26634
rect 23076 26616 23078 26634
rect 23100 26616 23102 26634
rect 23148 26616 23150 26634
rect 23196 26616 23198 26634
rect 23220 26616 23222 26634
rect 23244 26616 23246 26634
rect 23292 26616 23294 26634
rect 23316 26616 23318 26634
rect 23340 26616 23342 26634
rect 23388 26616 23390 26634
rect 23412 26616 23414 26634
rect 23436 26616 23438 26634
rect 23484 26616 23486 26634
rect 23532 26616 23534 26634
rect 23556 26616 23558 26634
rect 23580 26616 23582 26634
rect 23628 26616 23630 26634
rect 23652 26616 23654 26634
rect 23676 26616 23678 26634
rect 23724 26616 23726 26634
rect 23748 26616 23750 26634
rect 23772 26616 23774 26634
rect 23820 26616 23822 26634
rect 23868 26616 23870 26634
rect 23892 26616 23894 26634
rect 23916 26616 23918 26634
rect 23988 26616 23990 26634
rect 24012 26616 24014 26634
rect 24036 26616 24038 26634
rect 24084 26616 24086 26634
rect 24132 26616 24134 26634
rect 24228 26616 24230 26634
rect 24252 26616 24254 26634
rect 24300 26616 24302 26634
rect 24348 26616 24350 26634
rect 24372 26616 24374 26634
rect 24396 26616 24398 26634
rect 24468 26616 24470 26634
rect 24492 26616 24494 26634
rect 24516 26616 24518 26634
rect 24564 26616 24566 26634
rect 24588 26616 24590 26634
rect 24612 26616 24614 26634
rect 24660 26616 24662 26634
rect 24708 26616 24710 26634
rect 24732 26616 24734 26634
rect 24756 26616 24758 26634
rect 24828 26616 24830 26634
rect 24852 26616 24854 26634
rect 24876 26616 24878 26634
rect 24948 26616 24950 26634
rect 24972 26616 24974 26634
rect 24996 26616 24998 26634
rect 25044 26616 25046 26634
rect 25092 26616 25094 26634
rect 25140 26616 25142 26634
rect 25260 26616 25262 26634
rect 25356 26616 25358 26634
rect 25380 26616 25382 26634
rect 25452 26616 25454 26634
rect 25476 26616 25478 26634
rect 25500 26616 25502 26634
rect 25548 26616 25550 26634
rect 25572 26616 25574 26634
rect 25596 26616 25598 26634
rect 25644 26616 25646 26634
rect 27060 26616 27062 26634
rect 27108 26616 27110 26634
rect 27180 26616 27182 26634
rect 27276 26616 27278 26634
rect 27324 26616 27326 26634
rect 27372 26616 27374 26634
rect 27396 26616 27398 26634
rect 27420 26616 27422 26634
rect 27468 26616 27470 26634
rect 27516 26616 27518 26634
rect 27540 26616 27542 26634
rect 27564 26616 27566 26634
rect 28146 26622 28158 26631
rect 28866 26622 28878 26631
rect 29586 26622 29598 26631
rect 30306 26622 30318 26631
rect 28144 26617 28146 26622
rect 28864 26617 28866 26622
rect 29584 26617 29586 26622
rect 30304 26617 30306 26622
rect 30492 26616 30494 26634
rect 30540 26616 30542 26634
rect 30612 26616 30614 26634
rect 30636 26616 30638 26634
rect 30660 26616 30662 26634
rect 30708 26616 30710 26634
rect 30756 26616 30758 26634
rect 30780 26616 30782 26634
rect 30804 26616 30806 26634
rect 30852 26616 30854 26634
rect 30900 26616 30902 26634
rect 30924 26616 30926 26634
rect 30948 26616 30950 26634
rect 30996 26616 30998 26634
rect 31044 26616 31046 26634
rect 31068 26616 31070 26634
rect 31092 26616 31094 26634
rect 31140 26616 31142 26634
rect 31188 26616 31190 26634
rect 31236 26616 31238 26634
rect 32076 26616 32078 26634
rect 32100 26616 32102 26634
rect 32148 26616 32150 26634
rect -19052 26611 -15644 26616
rect -15584 26611 -10100 26616
rect -10040 26611 9412 26616
rect 9472 26611 14836 26616
rect 14896 26611 17860 26616
rect 17920 26611 22780 26616
rect 22840 26611 26188 26616
rect 26248 26611 26812 26616
rect 26872 26611 28158 26616
rect -18839 26558 -18835 26566
rect -18849 26552 -18839 26558
rect -18836 26544 -18835 26551
rect -18777 26544 -18774 26551
rect -18764 26544 -18763 26551
rect -18815 26527 -18798 26528
rect -18767 26527 -18709 26528
rect -18407 26527 -18349 26528
rect -18047 26527 -17989 26528
rect -17916 26527 -17914 26611
rect -17868 26527 -17866 26611
rect -17820 26527 -17818 26611
rect -17772 26527 -17770 26611
rect -17652 26589 -17650 26611
rect -17532 26527 -17530 26611
rect -17436 26527 -17434 26611
rect -17412 26527 -17410 26611
rect -17364 26527 -17362 26611
rect -17316 26527 -17314 26611
rect -17220 26527 -17218 26611
rect -17196 26527 -17194 26611
rect -17124 26527 -17122 26611
rect -17028 26527 -17026 26611
rect -16980 26589 -16978 26611
rect -16884 26581 -16882 26611
rect -16860 26527 -16858 26611
rect -16812 26527 -16810 26611
rect -16788 26527 -16786 26611
rect -16764 26527 -16762 26611
rect -16716 26527 -16714 26611
rect -16692 26527 -16690 26611
rect -16668 26527 -16666 26611
rect -16596 26527 -16594 26611
rect -16500 26527 -16498 26611
rect -16404 26527 -16402 26611
rect -16380 26527 -16378 26611
rect -16332 26527 -16330 26611
rect -16308 26527 -16306 26611
rect -16284 26527 -16282 26611
rect -16236 26527 -16234 26611
rect -16212 26527 -16210 26611
rect -16188 26527 -16186 26611
rect -15970 26608 -15954 26611
rect -15584 26609 -15570 26611
rect -15420 26581 -15418 26611
rect -15396 26581 -15394 26611
rect -15372 26527 -15370 26611
rect -15300 26527 -15298 26611
rect -15084 26527 -15082 26611
rect -15036 26527 -15034 26611
rect -14940 26589 -14938 26611
rect -14927 26566 -14924 26576
rect -14916 26568 -14914 26611
rect -14916 26566 -14913 26568
rect -14917 26552 -14913 26566
rect -14937 26544 -14934 26551
rect -14924 26544 -14923 26551
rect -14914 26544 -14913 26552
rect -14868 26527 -14866 26611
rect -14820 26568 -14818 26611
rect -14841 26544 -14838 26551
rect -14828 26544 -14827 26551
rect -14820 26544 -14817 26568
rect -14724 26527 -14722 26611
rect -14700 26528 -14698 26611
rect -14711 26527 -14677 26528
rect -14652 26527 -14650 26611
rect -14604 26527 -14602 26611
rect -14508 26527 -14506 26611
rect -14484 26581 -14482 26611
rect -14436 26527 -14434 26611
rect -14388 26527 -14386 26611
rect -14268 26527 -14266 26611
rect -14172 26527 -14170 26611
rect -14076 26527 -14074 26611
rect -14028 26527 -14026 26611
rect -13980 26527 -13978 26611
rect -13956 26527 -13954 26611
rect -13932 26527 -13930 26611
rect -13860 26527 -13858 26611
rect -13764 26527 -13762 26611
rect -13716 26527 -13714 26611
rect -13644 26527 -13642 26611
rect -13596 26527 -13594 26611
rect -13500 26527 -13498 26611
rect -13404 26527 -13402 26611
rect -13356 26527 -13354 26611
rect -13284 26527 -13282 26611
rect -12828 26527 -12826 26611
rect -12780 26527 -12778 26611
rect -12684 26527 -12682 26611
rect -12660 26527 -12658 26611
rect -12612 26527 -12610 26611
rect -12588 26527 -12586 26611
rect -12564 26527 -12562 26611
rect -12492 26527 -12490 26611
rect -12396 26527 -12394 26611
rect -12348 26527 -12346 26611
rect -12335 26527 -12301 26528
rect -12276 26527 -12274 26611
rect -12252 26527 -12250 26611
rect -12228 26527 -12226 26611
rect -12156 26527 -12154 26611
rect -12060 26527 -12058 26611
rect -12012 26527 -12010 26611
rect -11916 26527 -11914 26611
rect -11892 26527 -11890 26611
rect -11844 26527 -11842 26611
rect -11796 26527 -11794 26611
rect -11676 26527 -11674 26611
rect -11580 26527 -11578 26611
rect -11556 26527 -11554 26611
rect -11484 26527 -11482 26611
rect -11460 26527 -11458 26611
rect -11436 26527 -11434 26611
rect -11388 26527 -11386 26611
rect -11364 26527 -11362 26611
rect -11340 26527 -11338 26611
rect -11268 26527 -11266 26611
rect -11172 26527 -11170 26611
rect -11124 26527 -11122 26611
rect -11076 26527 -11074 26611
rect -11073 26544 -11070 26551
rect -11060 26544 -11059 26551
rect -11028 26527 -11026 26611
rect -10932 26589 -10930 26611
rect -10836 26581 -10834 26611
rect -10788 26527 -10786 26611
rect -10668 26527 -10666 26611
rect -10426 26608 -10410 26611
rect -10040 26609 -10026 26611
rect -9876 26527 -9874 26611
rect -9828 26527 -9826 26611
rect -9732 26527 -9730 26611
rect -9708 26527 -9706 26611
rect -9612 26527 -9610 26611
rect -9516 26527 -9514 26611
rect -9468 26527 -9466 26611
rect -9420 26527 -9418 26611
rect -9396 26527 -9394 26611
rect -9372 26527 -9370 26611
rect -9300 26527 -9298 26611
rect -9252 26527 -9250 26611
rect -9167 26566 -9164 26576
rect -9156 26566 -9154 26611
rect -9157 26552 -9154 26566
rect -9132 26527 -9130 26611
rect -9084 26527 -9082 26611
rect -9060 26568 -9058 26611
rect -9081 26544 -9078 26551
rect -9068 26544 -9067 26551
rect -9060 26544 -9057 26568
rect -9071 26527 -9037 26528
rect -9036 26527 -9034 26611
rect -8988 26527 -8986 26611
rect -8964 26589 -8962 26611
rect -8940 26527 -8938 26611
rect -8892 26527 -8890 26611
rect -8844 26527 -8842 26611
rect -8796 26527 -8794 26611
rect -8700 26527 -8698 26611
rect -8604 26527 -8602 26611
rect -8567 26566 -8564 26576
rect -8556 26566 -8554 26611
rect -8557 26552 -8554 26566
rect -8508 26527 -8506 26611
rect -8484 26527 -8482 26611
rect -8460 26568 -8458 26611
rect -8481 26544 -8478 26551
rect -8468 26544 -8467 26551
rect -8460 26544 -8457 26568
rect -8412 26527 -8410 26611
rect -8388 26527 -8386 26611
rect -8364 26527 -8362 26611
rect -8316 26527 -8314 26611
rect -8292 26527 -8290 26611
rect -8268 26527 -8266 26611
rect -8196 26527 -8194 26611
rect -8100 26527 -8098 26611
rect -8052 26527 -8050 26611
rect -7932 26527 -7930 26611
rect -7836 26527 -7834 26611
rect -7740 26527 -7738 26611
rect -7692 26527 -7690 26611
rect -7620 26527 -7618 26611
rect -7356 26527 -7354 26611
rect -7284 26527 -7282 26611
rect -7212 26527 -7210 26611
rect -7188 26527 -7186 26611
rect -7116 26527 -7114 26611
rect -7092 26589 -7090 26611
rect -7068 26527 -7066 26611
rect -6996 26589 -6994 26611
rect -6972 26527 -6970 26611
rect -6948 26527 -6946 26611
rect -6900 26581 -6898 26611
rect -6876 26527 -6874 26611
rect -6852 26527 -6850 26611
rect -6804 26527 -6802 26611
rect -6780 26527 -6778 26611
rect -6756 26527 -6754 26611
rect -6708 26527 -6706 26611
rect -6684 26527 -6682 26611
rect -6660 26527 -6658 26611
rect -6612 26527 -6610 26611
rect -6588 26527 -6586 26611
rect -6564 26527 -6562 26611
rect -6516 26527 -6514 26611
rect -6492 26527 -6490 26611
rect -6468 26527 -6466 26611
rect -6420 26527 -6418 26611
rect -6396 26527 -6394 26611
rect -6372 26527 -6370 26611
rect -6324 26527 -6322 26611
rect -6300 26527 -6298 26611
rect -6276 26527 -6274 26611
rect -6228 26527 -6226 26611
rect -6180 26527 -6178 26611
rect -6060 26527 -6058 26611
rect -5964 26527 -5962 26611
rect -5940 26527 -5938 26611
rect -5868 26527 -5866 26611
rect -5796 26589 -5794 26611
rect -5652 26527 -5650 26611
rect -5316 26527 -5314 26611
rect -5268 26527 -5266 26611
rect -5220 26589 -5218 26611
rect -5196 26527 -5194 26611
rect -5172 26527 -5170 26611
rect -5124 26589 -5122 26611
rect -5100 26527 -5098 26611
rect -5076 26527 -5074 26611
rect -5028 26581 -5026 26611
rect -4980 26527 -4978 26611
rect -4953 26544 -4950 26551
rect -4940 26544 -4939 26551
rect -18846 26523 -18798 26527
rect -18774 26523 -4963 26527
rect -18407 26518 -18404 26523
rect -18047 26518 -18044 26523
rect -17916 26520 -17914 26523
rect -18733 26504 -18730 26518
rect -18719 26510 -18715 26518
rect -18729 26504 -18719 26510
rect -18397 26504 -18394 26518
rect -18037 26504 -18034 26518
rect -18396 26503 -18394 26504
rect -18119 26503 -18061 26504
rect -18036 26503 -18034 26504
rect -17916 26503 -17913 26520
rect -17868 26504 -17866 26523
rect -17879 26503 -17845 26504
rect -17820 26503 -17818 26523
rect -17772 26503 -17770 26523
rect -17532 26503 -17530 26523
rect -17436 26503 -17434 26523
rect -17412 26503 -17410 26523
rect -17364 26503 -17362 26523
rect -17316 26503 -17314 26523
rect -17220 26504 -17218 26523
rect -17231 26503 -17197 26504
rect -17196 26503 -17194 26523
rect -17124 26503 -17122 26523
rect -17028 26503 -17026 26523
rect -16860 26503 -16858 26523
rect -16812 26503 -16810 26523
rect -16788 26504 -16786 26523
rect -16799 26503 -16765 26504
rect -16764 26503 -16762 26523
rect -16716 26503 -16714 26523
rect -16692 26503 -16690 26523
rect -16668 26503 -16666 26523
rect -16596 26503 -16594 26523
rect -16500 26503 -16498 26523
rect -16463 26503 -16405 26504
rect -16404 26503 -16402 26523
rect -16380 26503 -16378 26523
rect -16332 26503 -16330 26523
rect -16308 26503 -16306 26523
rect -16284 26503 -16282 26523
rect -16236 26503 -16234 26523
rect -16212 26503 -16210 26523
rect -16188 26503 -16186 26523
rect -15372 26503 -15370 26523
rect -15300 26503 -15298 26523
rect -15084 26503 -15082 26523
rect -15036 26503 -15034 26523
rect -14868 26503 -14866 26523
rect -14724 26503 -14722 26523
rect -14711 26518 -14708 26523
rect -14700 26518 -14698 26523
rect -14701 26504 -14698 26518
rect -14652 26503 -14650 26523
rect -14604 26520 -14602 26523
rect -14604 26503 -14601 26520
rect -14508 26503 -14506 26523
rect -14436 26503 -14434 26523
rect -14388 26503 -14386 26523
rect -14268 26503 -14266 26523
rect -14172 26503 -14170 26523
rect -14076 26503 -14074 26523
rect -14028 26503 -14026 26523
rect -13980 26503 -13978 26523
rect -13956 26503 -13954 26523
rect -13932 26503 -13930 26523
rect -13860 26503 -13858 26523
rect -13764 26503 -13762 26523
rect -13716 26503 -13714 26523
rect -13644 26503 -13642 26523
rect -13596 26503 -13594 26523
rect -13500 26503 -13498 26523
rect -13404 26503 -13402 26523
rect -13356 26503 -13354 26523
rect -13284 26503 -13282 26523
rect -12828 26503 -12826 26523
rect -12780 26503 -12778 26523
rect -12684 26503 -12682 26523
rect -12660 26503 -12658 26523
rect -12612 26504 -12610 26523
rect -12647 26503 -12589 26504
rect -12588 26503 -12586 26523
rect -12564 26503 -12562 26523
rect -12492 26503 -12490 26523
rect -12396 26503 -12394 26523
rect -12348 26503 -12346 26523
rect -12276 26503 -12274 26523
rect -12252 26503 -12250 26523
rect -12228 26520 -12226 26523
rect -12228 26503 -12225 26520
rect -12156 26503 -12154 26523
rect -12060 26503 -12058 26523
rect -12012 26503 -12010 26523
rect -11916 26503 -11914 26523
rect -11892 26503 -11890 26523
rect -11844 26503 -11842 26523
rect -11796 26503 -11794 26523
rect -11676 26503 -11674 26523
rect -11580 26503 -11578 26523
rect -11556 26503 -11554 26523
rect -11484 26503 -11482 26523
rect -11460 26503 -11458 26523
rect -11436 26503 -11434 26523
rect -11388 26503 -11386 26523
rect -11364 26503 -11362 26523
rect -11340 26503 -11338 26523
rect -11268 26503 -11266 26523
rect -11172 26503 -11170 26523
rect -11124 26503 -11122 26523
rect -11076 26503 -11074 26523
rect -11028 26503 -11026 26523
rect -10788 26503 -10786 26523
rect -10668 26503 -10666 26523
rect -9876 26503 -9874 26523
rect -9828 26503 -9826 26523
rect -9732 26503 -9730 26523
rect -9708 26503 -9706 26523
rect -9612 26503 -9610 26523
rect -9516 26503 -9514 26523
rect -9468 26503 -9466 26523
rect -9420 26503 -9418 26523
rect -9396 26503 -9394 26523
rect -9372 26503 -9370 26523
rect -9300 26503 -9298 26523
rect -9252 26503 -9250 26523
rect -9132 26503 -9130 26523
rect -9084 26503 -9082 26523
rect -9036 26503 -9034 26523
rect -8988 26503 -8986 26523
rect -8940 26503 -8938 26523
rect -8892 26503 -8890 26523
rect -8844 26503 -8842 26523
rect -8796 26503 -8794 26523
rect -8700 26503 -8698 26523
rect -8604 26503 -8602 26523
rect -8508 26503 -8506 26523
rect -8484 26503 -8482 26523
rect -8412 26504 -8410 26523
rect -8447 26503 -8389 26504
rect -8388 26503 -8386 26523
rect -8364 26503 -8362 26523
rect -8316 26503 -8314 26523
rect -8292 26503 -8290 26523
rect -8268 26503 -8266 26523
rect -8196 26503 -8194 26523
rect -8100 26503 -8098 26523
rect -8052 26503 -8050 26523
rect -7932 26503 -7930 26523
rect -7836 26503 -7834 26523
rect -7740 26503 -7738 26523
rect -7692 26503 -7690 26523
rect -7620 26503 -7618 26523
rect -7356 26503 -7354 26523
rect -7284 26503 -7282 26523
rect -7212 26503 -7210 26523
rect -7188 26503 -7186 26523
rect -7116 26503 -7114 26523
rect -7068 26503 -7066 26523
rect -6972 26503 -6970 26523
rect -6948 26503 -6946 26523
rect -6876 26503 -6874 26523
rect -6852 26503 -6850 26523
rect -6804 26503 -6802 26523
rect -6780 26503 -6778 26523
rect -6756 26503 -6754 26523
rect -6708 26503 -6706 26523
rect -6684 26503 -6682 26523
rect -6660 26503 -6658 26523
rect -6612 26503 -6610 26523
rect -6588 26503 -6586 26523
rect -6564 26503 -6562 26523
rect -6516 26503 -6514 26523
rect -6492 26503 -6490 26523
rect -6468 26503 -6466 26523
rect -6420 26503 -6418 26523
rect -6396 26503 -6394 26523
rect -6372 26503 -6370 26523
rect -6324 26503 -6322 26523
rect -6300 26503 -6298 26523
rect -6276 26503 -6274 26523
rect -6228 26503 -6226 26523
rect -6180 26503 -6178 26523
rect -6060 26503 -6058 26523
rect -5964 26503 -5962 26523
rect -5940 26503 -5938 26523
rect -5868 26503 -5866 26523
rect -5652 26503 -5650 26523
rect -5495 26503 -5461 26504
rect -5316 26503 -5314 26523
rect -5268 26503 -5266 26523
rect -5196 26503 -5194 26523
rect -5172 26503 -5170 26523
rect -5100 26503 -5098 26523
rect -5076 26503 -5074 26523
rect -4980 26503 -4978 26523
rect -4977 26520 -4963 26523
rect -4956 26520 -4953 26544
rect -4884 26527 -4882 26611
rect -4860 26527 -4858 26611
rect -4788 26527 -4786 26611
rect -4692 26527 -4690 26611
rect -4644 26527 -4642 26611
rect -4596 26527 -4594 26611
rect -4548 26527 -4546 26611
rect -4428 26527 -4426 26611
rect -4332 26527 -4330 26611
rect -4308 26527 -4306 26611
rect -4260 26527 -4258 26611
rect -4212 26527 -4210 26611
rect -4116 26527 -4114 26611
rect -4092 26527 -4090 26611
rect -4020 26527 -4018 26611
rect -3876 26527 -3874 26611
rect -3804 26528 -3802 26611
rect -3815 26527 -3781 26528
rect -3732 26527 -3730 26611
rect -3588 26527 -3586 26611
rect -3564 26527 -3562 26611
rect -3516 26527 -3514 26611
rect -3492 26527 -3490 26611
rect -3468 26527 -3466 26611
rect -3420 26527 -3418 26611
rect -3372 26589 -3370 26611
rect -3252 26527 -3250 26611
rect -3156 26527 -3154 26611
rect -3132 26527 -3130 26611
rect -3060 26527 -3058 26611
rect -3012 26527 -3010 26611
rect -2916 26527 -2914 26611
rect -2892 26527 -2890 26611
rect -2844 26527 -2842 26611
rect -2820 26527 -2818 26611
rect -2796 26527 -2794 26611
rect -2748 26527 -2746 26611
rect -2700 26527 -2698 26611
rect -2604 26527 -2602 26611
rect -2580 26527 -2578 26611
rect -2508 26589 -2506 26611
rect -2412 26581 -2410 26611
rect -2364 26527 -2362 26611
rect -2292 26527 -2290 26611
rect -2268 26527 -2266 26611
rect -2244 26527 -2242 26611
rect -2196 26589 -2194 26611
rect -2172 26527 -2170 26611
rect -2148 26527 -2146 26611
rect -2100 26581 -2098 26611
rect -2076 26527 -2074 26611
rect -2052 26527 -2050 26611
rect -1980 26527 -1978 26611
rect -1884 26527 -1882 26611
rect -1836 26527 -1834 26611
rect -1716 26527 -1714 26611
rect -1596 26527 -1594 26611
rect -1476 26527 -1474 26611
rect -1380 26527 -1378 26611
rect -1356 26527 -1354 26611
rect -1308 26527 -1306 26611
rect -1260 26527 -1258 26611
rect -1164 26589 -1162 26611
rect -1140 26527 -1138 26611
rect -1068 26581 -1066 26611
rect -852 26527 -850 26611
rect -804 26527 -802 26611
rect -756 26527 -754 26611
rect -708 26527 -706 26611
rect -612 26527 -610 26611
rect -588 26527 -586 26611
rect -540 26527 -538 26611
rect -516 26527 -514 26611
rect -492 26527 -490 26611
rect -444 26527 -442 26611
rect -396 26527 -394 26611
rect -300 26527 -298 26611
rect -276 26527 -274 26611
rect -204 26527 -202 26611
rect -108 26527 -106 26611
rect -60 26581 -58 26611
rect 12 26527 14 26611
rect 108 26527 110 26611
rect 156 26527 158 26611
rect 204 26527 206 26611
rect 228 26527 230 26611
rect 252 26527 254 26611
rect 300 26589 302 26611
rect 348 26527 350 26611
rect 468 26527 470 26611
rect 564 26527 566 26611
rect 588 26527 590 26611
rect 636 26527 638 26611
rect 660 26527 662 26611
rect 684 26527 686 26611
rect 732 26527 734 26611
rect 756 26527 758 26611
rect 780 26527 782 26611
rect 876 26527 878 26611
rect 972 26527 974 26611
rect 1020 26527 1022 26611
rect 1068 26527 1070 26611
rect 1092 26527 1094 26611
rect 1116 26527 1118 26611
rect 1164 26527 1166 26611
rect 1212 26527 1214 26611
rect 1308 26527 1310 26611
rect 1332 26527 1334 26611
rect 1380 26527 1382 26611
rect 1428 26527 1430 26611
rect 1524 26527 1526 26611
rect 1548 26527 1550 26611
rect 1596 26527 1598 26611
rect 1620 26527 1622 26611
rect 1644 26527 1646 26611
rect 1692 26527 1694 26611
rect 1716 26527 1718 26611
rect 1740 26527 1742 26611
rect 1788 26527 1790 26611
rect 1812 26589 1814 26611
rect 1836 26527 1838 26611
rect 1884 26527 1886 26611
rect 1908 26589 1910 26611
rect 1932 26527 1934 26611
rect 1980 26527 1982 26611
rect 2004 26581 2006 26611
rect 2028 26527 2030 26611
rect 2076 26527 2078 26611
rect 2100 26527 2102 26611
rect 2124 26527 2126 26611
rect 2172 26527 2174 26611
rect 2196 26527 2198 26611
rect 2220 26527 2222 26611
rect 2268 26527 2270 26611
rect 2292 26527 2294 26611
rect 2316 26527 2318 26611
rect 2364 26527 2366 26611
rect 2388 26589 2390 26611
rect 2412 26527 2414 26611
rect 2460 26527 2462 26611
rect 2484 26581 2486 26611
rect 2508 26527 2510 26611
rect 2556 26527 2558 26611
rect 2580 26527 2582 26611
rect 2604 26527 2606 26611
rect 2652 26527 2654 26611
rect 2676 26527 2678 26611
rect 2700 26527 2702 26611
rect 2748 26527 2750 26611
rect 2772 26527 2774 26611
rect 2796 26527 2798 26611
rect 2844 26527 2846 26611
rect 2868 26527 2870 26611
rect 2892 26527 2894 26611
rect 2940 26527 2942 26611
rect 3012 26527 3014 26611
rect 3108 26527 3110 26611
rect 3156 26527 3158 26611
rect 3252 26527 3254 26611
rect 3348 26527 3350 26611
rect 3396 26527 3398 26611
rect 3468 26527 3470 26611
rect 3492 26527 3494 26611
rect 3516 26581 3518 26611
rect 3588 26527 3590 26611
rect 3612 26527 3614 26611
rect 3636 26527 3638 26611
rect 3708 26527 3710 26611
rect 3732 26527 3734 26611
rect 3756 26527 3758 26611
rect 3804 26527 3806 26611
rect 3828 26527 3830 26611
rect 3852 26527 3854 26611
rect 3900 26589 3902 26611
rect 3924 26527 3926 26611
rect 3948 26527 3950 26611
rect 3996 26581 3998 26611
rect 4020 26527 4022 26611
rect 4044 26527 4046 26611
rect 4092 26527 4094 26611
rect 4116 26527 4118 26611
rect 4140 26527 4142 26611
rect 4188 26527 4190 26611
rect 4212 26527 4214 26611
rect 4236 26527 4238 26611
rect 4284 26589 4286 26611
rect 4308 26527 4310 26611
rect 4332 26527 4334 26611
rect 4380 26589 4382 26611
rect 4404 26527 4406 26611
rect 4428 26527 4430 26611
rect 4476 26589 4478 26611
rect 4500 26527 4502 26611
rect 4524 26527 4526 26611
rect 4596 26527 4598 26611
rect 4812 26589 4814 26611
rect 4860 26527 4862 26611
rect 4908 26581 4910 26611
rect 4956 26527 4958 26611
rect 4980 26527 4982 26611
rect 5004 26527 5006 26611
rect 5076 26527 5078 26611
rect 5100 26527 5102 26611
rect 5124 26527 5126 26611
rect 5172 26527 5174 26611
rect 5196 26527 5198 26611
rect 5220 26527 5222 26611
rect 5268 26527 5270 26611
rect 5292 26527 5294 26611
rect 5316 26589 5318 26611
rect 5388 26527 5390 26611
rect 5412 26581 5414 26611
rect 5436 26581 5438 26611
rect 5484 26527 5486 26611
rect 5508 26527 5510 26611
rect 5532 26527 5534 26611
rect 5580 26527 5582 26611
rect 5628 26527 5630 26611
rect 5724 26527 5726 26611
rect 5748 26527 5750 26611
rect 5796 26527 5798 26611
rect 5820 26527 5822 26611
rect 5844 26527 5846 26611
rect 5916 26527 5918 26611
rect 6132 26527 6134 26611
rect 6180 26527 6182 26611
rect 6228 26527 6230 26611
rect 6252 26527 6254 26611
rect 6276 26527 6278 26611
rect 6324 26527 6326 26611
rect 6372 26527 6374 26611
rect 6468 26589 6470 26611
rect 6492 26527 6494 26611
rect 6564 26581 6566 26611
rect 6588 26527 6590 26611
rect 6612 26527 6614 26611
rect 6660 26527 6662 26611
rect 6684 26527 6686 26611
rect 6708 26527 6710 26611
rect 6780 26527 6782 26611
rect 6804 26527 6806 26611
rect 6828 26527 6830 26611
rect 6876 26589 6878 26611
rect 6900 26527 6902 26611
rect 6924 26527 6926 26611
rect 6972 26581 6974 26611
rect 7020 26527 7022 26611
rect 7140 26527 7142 26611
rect 7236 26527 7238 26611
rect 7260 26527 7262 26611
rect 7332 26527 7334 26611
rect 7356 26527 7358 26611
rect 7380 26527 7382 26611
rect 7428 26527 7430 26611
rect 7452 26527 7454 26611
rect 7476 26527 7478 26611
rect 7524 26527 7526 26611
rect 7548 26527 7550 26611
rect 7572 26527 7574 26611
rect 7620 26527 7622 26611
rect 7644 26527 7646 26611
rect 7668 26527 7670 26611
rect 7716 26527 7718 26611
rect 7740 26527 7742 26611
rect 7764 26527 7766 26611
rect 7836 26527 7838 26611
rect 7860 26527 7862 26611
rect 7884 26527 7886 26611
rect 7932 26527 7934 26611
rect 7956 26527 7958 26611
rect 7980 26527 7982 26611
rect 8052 26527 8054 26611
rect 8148 26527 8150 26611
rect 8196 26527 8198 26611
rect 8244 26527 8246 26611
rect 8268 26527 8270 26611
rect 8292 26527 8294 26611
rect 8340 26527 8342 26611
rect 8364 26527 8366 26611
rect 8388 26527 8390 26611
rect 8436 26527 8438 26611
rect 8460 26527 8462 26611
rect 8484 26527 8486 26611
rect 8556 26527 8558 26611
rect 8580 26527 8582 26611
rect 8604 26527 8606 26611
rect 8676 26527 8678 26611
rect 8700 26527 8702 26611
rect 8724 26527 8726 26611
rect 8772 26527 8774 26611
rect 8820 26527 8822 26611
rect 8844 26527 8846 26611
rect 8868 26527 8870 26611
rect 9086 26608 9102 26611
rect 9472 26609 9486 26611
rect 9660 26527 9662 26611
rect 9684 26527 9686 26611
rect 9708 26527 9710 26611
rect 9756 26527 9758 26611
rect 9780 26527 9782 26611
rect 9804 26527 9806 26611
rect 9852 26527 9854 26611
rect 9876 26527 9878 26611
rect 9900 26527 9902 26611
rect 9948 26527 9950 26611
rect 9972 26527 9974 26611
rect 9996 26527 9998 26611
rect 10068 26527 10070 26611
rect 10092 26527 10094 26611
rect 10116 26527 10118 26611
rect 10164 26527 10166 26611
rect 10188 26527 10190 26611
rect 10212 26527 10214 26611
rect 10260 26527 10262 26611
rect 10284 26527 10286 26611
rect 10308 26527 10310 26611
rect 10380 26527 10382 26611
rect 10404 26527 10406 26611
rect 10428 26527 10430 26611
rect 10476 26527 10478 26611
rect 10500 26527 10502 26611
rect 10524 26527 10526 26611
rect 10572 26527 10574 26611
rect 10596 26527 10598 26611
rect 10620 26527 10622 26611
rect 10668 26527 10670 26611
rect 10692 26527 10694 26611
rect 10716 26527 10718 26611
rect 10788 26527 10790 26611
rect 10836 26527 10838 26611
rect 10956 26527 10958 26611
rect 11052 26527 11054 26611
rect 11076 26527 11078 26611
rect 11124 26527 11126 26611
rect 11172 26527 11174 26611
rect 11220 26527 11222 26611
rect 11340 26527 11342 26611
rect 11436 26527 11438 26611
rect 11532 26527 11534 26611
rect 11580 26527 11582 26611
rect 11628 26527 11630 26611
rect 11652 26589 11654 26611
rect 11676 26527 11678 26611
rect 11748 26581 11750 26611
rect 11772 26527 11774 26611
rect 11796 26527 11798 26611
rect 11844 26527 11846 26611
rect 11892 26527 11894 26611
rect 11988 26527 11990 26611
rect 12012 26581 12014 26611
rect 12084 26527 12086 26611
rect 12132 26527 12134 26611
rect 12228 26527 12230 26611
rect 12252 26527 12254 26611
rect 12300 26527 12302 26611
rect 12324 26527 12326 26611
rect 12348 26527 12350 26611
rect 12396 26527 12398 26611
rect 12420 26527 12422 26611
rect 12444 26527 12446 26611
rect 12492 26527 12494 26611
rect 12516 26527 12518 26611
rect 12540 26527 12542 26611
rect 12588 26527 12590 26611
rect 12636 26527 12638 26611
rect 12732 26527 12734 26611
rect 12756 26527 12758 26611
rect 12804 26527 12806 26611
rect 12828 26527 12830 26611
rect 12852 26527 12854 26611
rect 12900 26527 12902 26611
rect 12924 26589 12926 26611
rect 12948 26527 12950 26611
rect 13020 26581 13022 26611
rect 13044 26527 13046 26611
rect 13068 26527 13070 26611
rect 13116 26527 13118 26611
rect 13188 26581 13190 26611
rect 13284 26527 13286 26611
rect 13332 26527 13334 26611
rect 13428 26527 13430 26611
rect 13524 26527 13526 26611
rect 13572 26527 13574 26611
rect 13644 26527 13646 26611
rect 13668 26527 13670 26611
rect 13692 26581 13694 26611
rect 13764 26527 13766 26611
rect 13788 26589 13790 26611
rect 13812 26527 13814 26611
rect 13860 26527 13862 26611
rect 13884 26581 13886 26611
rect 13908 26527 13910 26611
rect 13956 26527 13958 26611
rect 14004 26527 14006 26611
rect 14100 26527 14102 26611
rect 14196 26527 14198 26611
rect 14209 26527 14243 26528
rect 14244 26527 14246 26611
rect 14292 26527 14294 26611
rect 14510 26608 14526 26611
rect 14896 26609 14910 26611
rect 15132 26527 15134 26611
rect 15228 26527 15230 26611
rect 15252 26527 15254 26611
rect 15300 26527 15302 26611
rect 15324 26527 15326 26611
rect 15348 26589 15350 26611
rect 15396 26527 15398 26611
rect 15420 26527 15422 26611
rect 15444 26581 15446 26611
rect 15492 26527 15494 26611
rect 15540 26527 15542 26611
rect 15636 26527 15638 26611
rect 15660 26527 15662 26611
rect 15708 26527 15710 26611
rect 15732 26527 15734 26611
rect 15756 26527 15758 26611
rect 15804 26527 15806 26611
rect 15828 26527 15830 26611
rect 15852 26527 15854 26611
rect 15900 26527 15902 26611
rect 15924 26589 15926 26611
rect 15948 26527 15950 26611
rect 15996 26527 15998 26611
rect 16020 26581 16022 26611
rect 16044 26527 16046 26611
rect 16092 26527 16094 26611
rect 16140 26527 16142 26611
rect 16236 26527 16238 26611
rect 16260 26527 16262 26611
rect 16308 26527 16310 26611
rect 16332 26527 16334 26611
rect 16356 26527 16358 26611
rect 16404 26527 16406 26611
rect 16452 26527 16454 26611
rect 16548 26527 16550 26611
rect 16572 26527 16574 26611
rect 16620 26527 16622 26611
rect 16644 26589 16646 26611
rect 16668 26527 16670 26611
rect 16716 26527 16718 26611
rect 16740 26581 16742 26611
rect 16764 26527 16766 26611
rect 16836 26527 16838 26611
rect 16884 26527 16886 26611
rect 16980 26527 16982 26611
rect 17004 26527 17006 26611
rect 17052 26527 17054 26611
rect 17100 26527 17102 26611
rect 17196 26527 17198 26611
rect 17220 26527 17222 26611
rect 17268 26589 17270 26611
rect 17292 26527 17294 26611
rect 17316 26527 17318 26611
rect 17534 26608 17550 26611
rect 17920 26609 17934 26611
rect 18084 26527 18086 26611
rect 18108 26589 18110 26611
rect 18132 26527 18134 26611
rect 18180 26589 18182 26611
rect 18145 26527 18179 26528
rect 18252 26527 18254 26611
rect 18348 26589 18350 26611
rect 18396 26527 18398 26611
rect 18492 26527 18494 26611
rect 18516 26527 18518 26611
rect 18564 26527 18566 26611
rect 18588 26528 18590 26611
rect 18577 26527 18611 26528
rect 18612 26527 18614 26611
rect 18660 26527 18662 26611
rect 18684 26527 18686 26611
rect 18708 26527 18710 26611
rect 18756 26527 18758 26611
rect 18780 26589 18782 26611
rect 18804 26527 18806 26611
rect 18852 26527 18854 26611
rect 18876 26581 18878 26611
rect 18900 26527 18902 26611
rect 18948 26589 18950 26611
rect 18996 26527 18998 26611
rect 19020 26527 19022 26611
rect 19044 26581 19046 26611
rect 19092 26527 19094 26611
rect 19116 26527 19118 26611
rect 19140 26527 19142 26611
rect 19188 26527 19190 26611
rect 19236 26527 19238 26611
rect 19332 26527 19334 26611
rect 19428 26589 19430 26611
rect 19476 26527 19478 26611
rect 19524 26581 19526 26611
rect 19572 26589 19574 26611
rect 19596 26589 19598 26611
rect 19620 26527 19622 26611
rect 19668 26589 19670 26611
rect 19692 26581 19694 26611
rect 19716 26527 19718 26611
rect 19764 26581 19766 26611
rect 19812 26528 19814 26611
rect 19777 26527 19835 26528
rect 19836 26527 19838 26611
rect 19860 26527 19862 26611
rect 19932 26527 19934 26611
rect 19956 26527 19958 26611
rect 19980 26527 19982 26611
rect 20028 26527 20030 26611
rect 20052 26527 20054 26611
rect 20076 26527 20078 26611
rect 20148 26527 20150 26611
rect 20172 26527 20174 26611
rect 20196 26527 20198 26611
rect 20244 26589 20246 26611
rect 20268 26527 20270 26611
rect 20292 26527 20294 26611
rect 20340 26581 20342 26611
rect 20388 26527 20390 26611
rect 20484 26589 20486 26611
rect 20415 26544 20418 26551
rect 20428 26544 20429 26551
rect -4950 26523 20405 26527
rect -4956 26503 -4954 26520
rect -4884 26503 -4882 26523
rect -4860 26503 -4858 26523
rect -4788 26503 -4786 26523
rect -4692 26503 -4690 26523
rect -4644 26503 -4642 26523
rect -4596 26503 -4594 26523
rect -4548 26503 -4546 26523
rect -4428 26503 -4426 26523
rect -4332 26503 -4330 26523
rect -4308 26503 -4306 26523
rect -4260 26503 -4258 26523
rect -4212 26503 -4210 26523
rect -4116 26503 -4114 26523
rect -4092 26503 -4090 26523
rect -4020 26503 -4018 26523
rect -3876 26503 -3874 26523
rect -3815 26518 -3812 26523
rect -3804 26518 -3802 26523
rect -3805 26504 -3802 26518
rect -3732 26503 -3730 26523
rect -3588 26503 -3586 26523
rect -3564 26503 -3562 26523
rect -3516 26503 -3514 26523
rect -3492 26503 -3490 26523
rect -3468 26503 -3466 26523
rect -3420 26503 -3418 26523
rect -3252 26503 -3250 26523
rect -3156 26503 -3154 26523
rect -3132 26503 -3130 26523
rect -3060 26503 -3058 26523
rect -3012 26503 -3010 26523
rect -2975 26503 -2917 26504
rect -2916 26503 -2914 26523
rect -2892 26503 -2890 26523
rect -2844 26503 -2842 26523
rect -2820 26503 -2818 26523
rect -2796 26503 -2794 26523
rect -2748 26503 -2746 26523
rect -2700 26503 -2698 26523
rect -2604 26503 -2602 26523
rect -2580 26503 -2578 26523
rect -2364 26503 -2362 26523
rect -2292 26503 -2290 26523
rect -2268 26503 -2266 26523
rect -2244 26503 -2242 26523
rect -2172 26503 -2170 26523
rect -2148 26503 -2146 26523
rect -2076 26503 -2074 26523
rect -2052 26503 -2050 26523
rect -1980 26503 -1978 26523
rect -1884 26503 -1882 26523
rect -1836 26503 -1834 26523
rect -1716 26503 -1714 26523
rect -1596 26503 -1594 26523
rect -1476 26503 -1474 26523
rect -1380 26503 -1378 26523
rect -1356 26503 -1354 26523
rect -1308 26503 -1306 26523
rect -1260 26503 -1258 26523
rect -1140 26503 -1138 26523
rect -1103 26503 -1045 26504
rect -852 26503 -850 26523
rect -804 26503 -802 26523
rect -756 26503 -754 26523
rect -708 26503 -706 26523
rect -612 26503 -610 26523
rect -588 26503 -586 26523
rect -540 26503 -538 26523
rect -516 26503 -514 26523
rect -492 26503 -490 26523
rect -444 26503 -442 26523
rect -396 26503 -394 26523
rect -300 26503 -298 26523
rect -276 26503 -274 26523
rect -204 26503 -202 26523
rect -108 26503 -106 26523
rect 12 26503 14 26523
rect 108 26503 110 26523
rect 156 26503 158 26523
rect 204 26503 206 26523
rect 228 26503 230 26523
rect 252 26503 254 26523
rect 348 26503 350 26523
rect 468 26503 470 26523
rect 564 26503 566 26523
rect 588 26503 590 26523
rect 636 26503 638 26523
rect 660 26503 662 26523
rect 684 26503 686 26523
rect 732 26503 734 26523
rect 756 26503 758 26523
rect 780 26503 782 26523
rect 876 26503 878 26523
rect 972 26503 974 26523
rect 1020 26503 1022 26523
rect 1068 26503 1070 26523
rect 1092 26503 1094 26523
rect 1116 26503 1118 26523
rect 1164 26503 1166 26523
rect 1212 26503 1214 26523
rect 1308 26503 1310 26523
rect 1332 26503 1334 26523
rect 1380 26503 1382 26523
rect 1428 26503 1430 26523
rect 1524 26503 1526 26523
rect 1548 26503 1550 26523
rect 1596 26503 1598 26523
rect 1620 26503 1622 26523
rect 1644 26503 1646 26523
rect 1692 26503 1694 26523
rect 1716 26503 1718 26523
rect 1740 26503 1742 26523
rect 1788 26503 1790 26523
rect 1836 26503 1838 26523
rect 1884 26503 1886 26523
rect 1932 26503 1934 26523
rect 1980 26503 1982 26523
rect 2028 26503 2030 26523
rect 2076 26503 2078 26523
rect 2100 26503 2102 26523
rect 2124 26503 2126 26523
rect 2172 26503 2174 26523
rect 2196 26503 2198 26523
rect 2220 26503 2222 26523
rect 2268 26503 2270 26523
rect 2292 26503 2294 26523
rect 2316 26503 2318 26523
rect 2364 26503 2366 26523
rect 2412 26503 2414 26523
rect 2460 26503 2462 26523
rect 2508 26503 2510 26523
rect 2556 26503 2558 26523
rect 2580 26503 2582 26523
rect 2604 26503 2606 26523
rect 2652 26503 2654 26523
rect 2676 26503 2678 26523
rect 2700 26503 2702 26523
rect 2748 26503 2750 26523
rect 2772 26503 2774 26523
rect 2796 26503 2798 26523
rect 2844 26503 2846 26523
rect 2868 26503 2870 26523
rect 2892 26503 2894 26523
rect 2940 26503 2942 26523
rect 3012 26503 3014 26523
rect 3108 26503 3110 26523
rect 3156 26503 3158 26523
rect 3252 26503 3254 26523
rect 3348 26503 3350 26523
rect 3396 26503 3398 26523
rect 3468 26503 3470 26523
rect 3492 26503 3494 26523
rect 3588 26503 3590 26523
rect 3612 26503 3614 26523
rect 3636 26503 3638 26523
rect 3708 26503 3710 26523
rect 3732 26503 3734 26523
rect 3756 26504 3758 26523
rect 3745 26503 3779 26504
rect 3804 26503 3806 26523
rect 3828 26503 3830 26523
rect 3852 26504 3854 26523
rect 3841 26503 3875 26504
rect 3924 26503 3926 26523
rect 3948 26503 3950 26523
rect 4020 26503 4022 26523
rect 4044 26503 4046 26523
rect 4092 26503 4094 26523
rect 4116 26503 4118 26523
rect 4140 26503 4142 26523
rect 4188 26503 4190 26523
rect 4212 26503 4214 26523
rect 4236 26503 4238 26523
rect 4308 26503 4310 26523
rect 4332 26503 4334 26523
rect 4404 26503 4406 26523
rect 4428 26504 4430 26523
rect 4417 26503 4451 26504
rect 4500 26503 4502 26523
rect 4524 26503 4526 26523
rect 4596 26503 4598 26523
rect 4860 26503 4862 26523
rect 4956 26503 4958 26523
rect 4980 26503 4982 26523
rect 5004 26503 5006 26523
rect 5076 26503 5078 26523
rect 5100 26503 5102 26523
rect 5124 26503 5126 26523
rect 5172 26503 5174 26523
rect 5196 26503 5198 26523
rect 5220 26503 5222 26523
rect 5268 26503 5270 26523
rect 5292 26503 5294 26523
rect 5388 26503 5390 26523
rect 5484 26503 5486 26523
rect 5508 26503 5510 26523
rect 5532 26503 5534 26523
rect 5580 26503 5582 26523
rect 5628 26503 5630 26523
rect 5724 26503 5726 26523
rect 5748 26503 5750 26523
rect 5796 26503 5798 26523
rect 5820 26503 5822 26523
rect 5844 26503 5846 26523
rect 5916 26503 5918 26523
rect 6132 26503 6134 26523
rect 6180 26503 6182 26523
rect 6228 26503 6230 26523
rect 6252 26503 6254 26523
rect 6276 26503 6278 26523
rect 6324 26503 6326 26523
rect 6372 26503 6374 26523
rect 6492 26503 6494 26523
rect 6588 26503 6590 26523
rect 6612 26503 6614 26523
rect 6660 26503 6662 26523
rect 6684 26503 6686 26523
rect 6708 26503 6710 26523
rect 6780 26503 6782 26523
rect 6804 26503 6806 26523
rect 6828 26503 6830 26523
rect 6900 26503 6902 26523
rect 6924 26503 6926 26523
rect 7020 26503 7022 26523
rect 7140 26503 7142 26523
rect 7236 26503 7238 26523
rect 7260 26504 7262 26523
rect 7249 26503 7283 26504
rect 7332 26503 7334 26523
rect 7356 26503 7358 26523
rect 7380 26503 7382 26523
rect 7428 26503 7430 26523
rect 7452 26503 7454 26523
rect 7476 26503 7478 26523
rect 7524 26503 7526 26523
rect 7548 26503 7550 26523
rect 7572 26503 7574 26523
rect 7620 26503 7622 26523
rect 7644 26503 7646 26523
rect 7668 26503 7670 26523
rect 7716 26503 7718 26523
rect 7740 26503 7742 26523
rect 7764 26504 7766 26523
rect 7753 26503 7787 26504
rect 7836 26503 7838 26523
rect 7860 26503 7862 26523
rect 7884 26503 7886 26523
rect 7932 26503 7934 26523
rect 7956 26503 7958 26523
rect 7980 26503 7982 26523
rect 8052 26503 8054 26523
rect 8148 26503 8150 26523
rect 8196 26503 8198 26523
rect 8244 26503 8246 26523
rect 8268 26503 8270 26523
rect 8292 26503 8294 26523
rect 8340 26503 8342 26523
rect 8364 26503 8366 26523
rect 8388 26503 8390 26523
rect 8436 26503 8438 26523
rect 8460 26503 8462 26523
rect 8484 26504 8486 26523
rect 8473 26503 8507 26504
rect 8556 26503 8558 26523
rect 8580 26503 8582 26523
rect 8604 26503 8606 26523
rect 8676 26503 8678 26523
rect 8700 26503 8702 26523
rect 8724 26503 8726 26523
rect 8772 26503 8774 26523
rect 8820 26503 8822 26523
rect 8844 26503 8846 26523
rect 8868 26503 8870 26523
rect 9505 26503 9563 26504
rect 9660 26503 9662 26523
rect 9684 26503 9686 26523
rect 9708 26503 9710 26523
rect 9756 26503 9758 26523
rect 9780 26503 9782 26523
rect 9804 26503 9806 26523
rect 9852 26503 9854 26523
rect 9876 26503 9878 26523
rect 9900 26503 9902 26523
rect 9948 26503 9950 26523
rect 9972 26503 9974 26523
rect 9996 26503 9998 26523
rect 10068 26503 10070 26523
rect 10092 26503 10094 26523
rect 10116 26503 10118 26523
rect 10164 26503 10166 26523
rect 10188 26503 10190 26523
rect 10212 26503 10214 26523
rect 10260 26503 10262 26523
rect 10284 26503 10286 26523
rect 10308 26503 10310 26523
rect 10380 26503 10382 26523
rect 10404 26503 10406 26523
rect 10428 26503 10430 26523
rect 10476 26503 10478 26523
rect 10500 26503 10502 26523
rect 10524 26503 10526 26523
rect 10572 26503 10574 26523
rect 10596 26503 10598 26523
rect 10620 26503 10622 26523
rect 10668 26503 10670 26523
rect 10692 26503 10694 26523
rect 10716 26503 10718 26523
rect 10788 26503 10790 26523
rect 10836 26503 10838 26523
rect 10956 26503 10958 26523
rect 11052 26503 11054 26523
rect 11076 26503 11078 26523
rect 11124 26503 11126 26523
rect 11172 26503 11174 26523
rect 11220 26503 11222 26523
rect 11340 26503 11342 26523
rect 11436 26503 11438 26523
rect 11532 26503 11534 26523
rect 11580 26503 11582 26523
rect 11628 26503 11630 26523
rect 11676 26503 11678 26523
rect 11772 26503 11774 26523
rect 11796 26503 11798 26523
rect 11844 26503 11846 26523
rect 11892 26503 11894 26523
rect 11988 26503 11990 26523
rect 12084 26503 12086 26523
rect 12132 26503 12134 26523
rect 12228 26503 12230 26523
rect 12252 26503 12254 26523
rect 12300 26503 12302 26523
rect 12324 26503 12326 26523
rect 12348 26503 12350 26523
rect 12396 26503 12398 26523
rect 12420 26503 12422 26523
rect 12444 26503 12446 26523
rect 12492 26503 12494 26523
rect 12516 26503 12518 26523
rect 12540 26503 12542 26523
rect 12588 26503 12590 26523
rect 12636 26503 12638 26523
rect 12732 26503 12734 26523
rect 12756 26503 12758 26523
rect 12804 26503 12806 26523
rect 12828 26503 12830 26523
rect 12852 26503 12854 26523
rect 12900 26503 12902 26523
rect 12948 26503 12950 26523
rect 13044 26503 13046 26523
rect 13068 26503 13070 26523
rect 13116 26503 13118 26523
rect 13284 26503 13286 26523
rect 13332 26503 13334 26523
rect 13428 26503 13430 26523
rect 13524 26503 13526 26523
rect 13572 26503 13574 26523
rect 13644 26503 13646 26523
rect 13668 26503 13670 26523
rect 13764 26503 13766 26523
rect 13812 26503 13814 26523
rect 13860 26503 13862 26523
rect 13908 26503 13910 26523
rect 13956 26503 13958 26523
rect 14004 26503 14006 26523
rect 14100 26503 14102 26523
rect 14196 26503 14198 26523
rect 14244 26503 14246 26523
rect 14292 26503 14294 26523
rect 15132 26503 15134 26523
rect 15228 26503 15230 26523
rect 15252 26503 15254 26523
rect 15300 26503 15302 26523
rect 15324 26503 15326 26523
rect 15396 26503 15398 26523
rect 15420 26503 15422 26523
rect 15492 26503 15494 26523
rect 15540 26503 15542 26523
rect 15636 26503 15638 26523
rect 15660 26503 15662 26523
rect 15708 26503 15710 26523
rect 15732 26503 15734 26523
rect 15756 26503 15758 26523
rect 15804 26503 15806 26523
rect 15828 26503 15830 26523
rect 15852 26503 15854 26523
rect 15900 26503 15902 26523
rect 15948 26503 15950 26523
rect 15996 26503 15998 26523
rect 16044 26503 16046 26523
rect 16092 26503 16094 26523
rect 16140 26503 16142 26523
rect 16236 26503 16238 26523
rect 16260 26503 16262 26523
rect 16308 26503 16310 26523
rect 16332 26503 16334 26523
rect 16356 26503 16358 26523
rect 16404 26503 16406 26523
rect 16452 26503 16454 26523
rect 16548 26503 16550 26523
rect 16572 26503 16574 26523
rect 16620 26503 16622 26523
rect 16668 26503 16670 26523
rect 16716 26503 16718 26523
rect 16764 26503 16766 26523
rect 16836 26503 16838 26523
rect 16884 26503 16886 26523
rect 16980 26503 16982 26523
rect 17004 26503 17006 26523
rect 17052 26503 17054 26523
rect 17100 26503 17102 26523
rect 17196 26503 17198 26523
rect 17220 26503 17222 26523
rect 17292 26503 17294 26523
rect 17316 26503 17318 26523
rect 18084 26503 18086 26523
rect 18132 26503 18134 26523
rect 18252 26520 18254 26523
rect 18252 26503 18255 26520
rect 18396 26503 18398 26523
rect 18492 26503 18494 26523
rect 18516 26503 18518 26523
rect 18564 26503 18566 26523
rect 18577 26518 18580 26523
rect 18588 26518 18590 26523
rect 18587 26504 18590 26518
rect 18612 26503 18614 26523
rect 18660 26503 18662 26523
rect 18684 26520 18686 26523
rect 18684 26503 18687 26520
rect 18708 26503 18710 26523
rect 18756 26503 18758 26523
rect 18804 26503 18806 26523
rect 18852 26503 18854 26523
rect 18900 26503 18902 26523
rect 18996 26503 18998 26523
rect 19020 26503 19022 26523
rect 19092 26503 19094 26523
rect 19116 26503 19118 26523
rect 19140 26503 19142 26523
rect 19188 26503 19190 26523
rect 19236 26503 19238 26523
rect 19332 26503 19334 26523
rect 19476 26503 19478 26523
rect 19620 26503 19622 26523
rect 19716 26503 19718 26523
rect 19777 26518 19780 26523
rect 19801 26518 19804 26523
rect 19812 26518 19814 26523
rect 19787 26504 19790 26518
rect 19811 26504 19814 26518
rect 19788 26503 19790 26504
rect 19836 26503 19838 26523
rect 19860 26503 19862 26523
rect 19884 26503 19887 26520
rect 19932 26503 19934 26523
rect 19956 26503 19958 26523
rect 19980 26503 19982 26523
rect 20028 26503 20030 26523
rect 20052 26503 20054 26523
rect 20076 26503 20078 26523
rect 20148 26503 20150 26523
rect 20172 26503 20174 26523
rect 20196 26503 20198 26523
rect 20268 26503 20270 26523
rect 20292 26503 20294 26523
rect 20388 26503 20390 26523
rect 20391 26520 20405 26523
rect 20412 26520 20415 26544
rect 20508 26527 20510 26611
rect 20556 26527 20558 26611
rect 20580 26581 20582 26611
rect 20604 26527 20606 26611
rect 20700 26589 20702 26611
rect 20916 26527 20918 26611
rect 20964 26527 20966 26611
rect 21012 26527 21014 26611
rect 21060 26527 21062 26611
rect 21084 26527 21086 26611
rect 21108 26527 21110 26611
rect 21156 26589 21158 26611
rect 21204 26527 21206 26611
rect 21300 26527 21302 26611
rect 21324 26527 21326 26611
rect 21372 26581 21374 26611
rect 21420 26589 21422 26611
rect 21444 26527 21446 26611
rect 21468 26527 21470 26611
rect 21516 26581 21518 26611
rect 21540 26589 21542 26611
rect 21564 26527 21566 26611
rect 21612 26527 21614 26611
rect 21660 26589 21662 26611
rect 21684 26527 21686 26611
rect 21708 26527 21710 26611
rect 21780 26589 21782 26611
rect 21804 26527 21806 26611
rect 21828 26527 21830 26611
rect 21900 26589 21902 26611
rect 21924 26527 21926 26611
rect 21948 26527 21950 26611
rect 22020 26589 22022 26611
rect 22044 26527 22046 26611
rect 22068 26527 22070 26611
rect 22116 26581 22118 26611
rect 22164 26589 22166 26611
rect 22188 26527 22190 26611
rect 22212 26527 22214 26611
rect 22454 26608 22470 26611
rect 22840 26609 22854 26611
rect 23004 26527 23006 26611
rect 23052 26527 23054 26611
rect 23076 26527 23078 26611
rect 23100 26527 23102 26611
rect 23148 26527 23150 26611
rect 23196 26589 23198 26611
rect 23220 26527 23222 26611
rect 23244 26527 23246 26611
rect 23292 26589 23294 26611
rect 23316 26527 23318 26611
rect 23340 26527 23342 26611
rect 23388 26581 23390 26611
rect 23412 26527 23414 26611
rect 23436 26589 23438 26611
rect 23484 26589 23486 26611
rect 23532 26581 23534 26611
rect 23556 26527 23558 26611
rect 23580 26581 23582 26611
rect 23628 26527 23630 26611
rect 23652 26527 23654 26611
rect 23676 26527 23678 26611
rect 23724 26527 23726 26611
rect 23748 26527 23750 26611
rect 23772 26527 23774 26611
rect 23820 26527 23822 26611
rect 23868 26527 23870 26611
rect 23892 26527 23894 26611
rect 23916 26527 23918 26611
rect 23988 26527 23990 26611
rect 24012 26527 24014 26611
rect 24036 26581 24038 26611
rect 24084 26527 24086 26611
rect 24132 26589 24134 26611
rect 24228 26581 24230 26611
rect 24252 26528 24254 26611
rect 24300 26581 24302 26611
rect 24348 26589 24350 26611
rect 24241 26527 24275 26528
rect 24372 26527 24374 26611
rect 24396 26527 24398 26611
rect 24468 26589 24470 26611
rect 24492 26527 24494 26611
rect 24516 26527 24518 26611
rect 24564 26589 24566 26611
rect 24588 26527 24590 26611
rect 24612 26527 24614 26611
rect 24660 26581 24662 26611
rect 24708 26527 24710 26611
rect 24732 26527 24734 26611
rect 24756 26527 24758 26611
rect 24828 26589 24830 26611
rect 24852 26527 24854 26611
rect 24876 26527 24878 26611
rect 24948 26589 24950 26611
rect 24972 26527 24974 26611
rect 24996 26527 24998 26611
rect 25044 26581 25046 26611
rect 25092 26527 25094 26611
rect 25140 26589 25142 26611
rect 25095 26544 25098 26551
rect 25108 26544 25109 26551
rect 25260 26527 25262 26611
rect 25356 26527 25358 26611
rect 25380 26527 25382 26611
rect 25452 26527 25454 26611
rect 25476 26527 25478 26611
rect 25500 26527 25502 26611
rect 25548 26589 25550 26611
rect 25572 26527 25574 26611
rect 25596 26527 25598 26611
rect 25644 26581 25646 26611
rect 25862 26608 25878 26611
rect 26248 26609 26262 26611
rect 26486 26608 26502 26611
rect 26872 26609 26886 26611
rect 27060 26527 27062 26611
rect 27108 26527 27110 26611
rect 27180 26527 27182 26611
rect 27276 26589 27278 26611
rect 27324 26527 27326 26611
rect 27372 26589 27374 26611
rect 27396 26527 27398 26611
rect 27420 26527 27422 26611
rect 27468 26581 27470 26611
rect 27516 26589 27518 26611
rect 27540 26527 27542 26611
rect 27564 26527 27566 26611
rect 27782 26608 27798 26611
rect 28144 26608 28158 26611
rect 28208 26611 28878 26616
rect 28208 26609 28222 26611
rect 28502 26608 28518 26611
rect 28864 26608 28878 26611
rect 28928 26611 29598 26616
rect 28928 26609 28942 26611
rect 29222 26608 29238 26611
rect 29584 26608 29598 26611
rect 29648 26611 30318 26616
rect 29648 26609 29662 26611
rect 29942 26608 29958 26611
rect 30304 26608 30318 26611
rect 30368 26611 31804 26616
rect 31864 26611 32194 26616
rect 30368 26609 30382 26611
rect 30492 26581 30494 26611
rect 30540 26581 30542 26611
rect 30612 26589 30614 26611
rect 30636 26527 30638 26611
rect 30660 26527 30662 26611
rect 30708 26581 30710 26611
rect 30756 26589 30758 26611
rect 30780 26527 30782 26611
rect 30804 26527 30806 26611
rect 30852 26581 30854 26611
rect 30900 26589 30902 26611
rect 30924 26527 30926 26611
rect 30948 26527 30950 26611
rect 30996 26581 30998 26611
rect 31044 26589 31046 26611
rect 31068 26527 31070 26611
rect 31092 26527 31094 26611
rect 31140 26581 31142 26611
rect 31188 26527 31190 26611
rect 31236 26527 31238 26611
rect 31478 26608 31494 26611
rect 31864 26609 31878 26611
rect 32076 26527 32078 26611
rect 32100 26527 32102 26611
rect 32148 26581 32150 26611
rect 32113 26527 32147 26528
rect 20418 26523 32147 26527
rect 20412 26503 20414 26520
rect 20508 26503 20510 26523
rect 20556 26503 20558 26523
rect 20604 26503 20606 26523
rect 20916 26503 20918 26523
rect 20964 26503 20966 26523
rect 21012 26503 21014 26523
rect 21060 26503 21062 26523
rect 21084 26503 21086 26523
rect 21108 26503 21110 26523
rect 21204 26503 21206 26523
rect 21300 26503 21302 26523
rect 21324 26503 21326 26523
rect 21444 26503 21446 26523
rect 21468 26503 21470 26523
rect 21564 26503 21566 26523
rect 21612 26503 21614 26523
rect 21684 26503 21686 26523
rect 21708 26503 21710 26523
rect 21804 26503 21806 26523
rect 21828 26503 21830 26523
rect 21924 26503 21926 26523
rect 21948 26503 21950 26523
rect 22044 26503 22046 26523
rect 22068 26503 22070 26523
rect 22188 26503 22190 26523
rect 22212 26503 22214 26523
rect 23004 26503 23006 26523
rect 23052 26503 23054 26523
rect 23076 26503 23078 26523
rect 23100 26503 23102 26523
rect 23148 26503 23150 26523
rect 23220 26503 23222 26523
rect 23244 26503 23246 26523
rect 23316 26503 23318 26523
rect 23340 26503 23342 26523
rect 23412 26503 23414 26523
rect 23556 26503 23558 26523
rect 23628 26503 23630 26523
rect 23652 26503 23654 26523
rect 23676 26503 23678 26523
rect 23724 26503 23726 26523
rect 23748 26504 23750 26523
rect 23737 26503 23771 26504
rect 23772 26503 23774 26523
rect 23820 26503 23822 26523
rect 23868 26503 23870 26523
rect 23892 26503 23894 26523
rect 23916 26503 23918 26523
rect 23988 26503 23990 26523
rect 24012 26503 24014 26523
rect 24084 26503 24086 26523
rect 24241 26518 24244 26523
rect 24252 26518 24254 26523
rect 24251 26504 24254 26518
rect 24372 26503 24374 26523
rect 24396 26503 24398 26523
rect 24492 26503 24494 26523
rect 24516 26503 24518 26523
rect 24588 26503 24590 26523
rect 24612 26503 24614 26523
rect 24708 26503 24710 26523
rect 24732 26503 24734 26523
rect 24756 26503 24758 26523
rect 24852 26503 24854 26523
rect 24876 26503 24878 26523
rect 24972 26503 24974 26523
rect 24996 26503 24998 26523
rect 25092 26503 25094 26523
rect 25260 26503 25262 26523
rect 25356 26503 25358 26523
rect 25380 26503 25382 26523
rect 25452 26503 25454 26523
rect 25476 26503 25478 26523
rect 25500 26503 25502 26523
rect 25572 26503 25574 26523
rect 25596 26503 25598 26523
rect 27060 26503 27062 26523
rect 27108 26503 27110 26523
rect 27180 26503 27182 26523
rect 27324 26503 27326 26523
rect 27396 26503 27398 26523
rect 27420 26503 27422 26523
rect 27540 26503 27542 26523
rect 27564 26503 27566 26523
rect 30636 26503 30638 26523
rect 30660 26503 30662 26523
rect 30780 26503 30782 26523
rect 30804 26503 30806 26523
rect 30924 26503 30926 26523
rect 30948 26503 30950 26523
rect 31068 26503 31070 26523
rect 31092 26503 31094 26523
rect 31188 26503 31190 26523
rect 31236 26503 31238 26523
rect 31897 26503 31955 26504
rect 32076 26503 32078 26523
rect 32100 26504 32102 26523
rect 32089 26503 32123 26504
rect -18798 26499 -18750 26503
rect -18729 26499 -18667 26503
rect -18729 26496 -18715 26499
rect -18681 26496 -18667 26499
rect -18657 26499 -18307 26503
rect -18657 26496 -18643 26499
rect -18750 26479 -18733 26480
rect -18527 26479 -18469 26480
rect -18396 26479 -18394 26499
rect -18321 26496 -18307 26499
rect -18297 26499 -17947 26503
rect -18297 26496 -18283 26499
rect -18119 26494 -18116 26499
rect -18109 26480 -18106 26494
rect -18108 26479 -18106 26480
rect -18036 26479 -18034 26499
rect -17961 26496 -17947 26499
rect -17937 26499 19877 26503
rect -17937 26496 -17923 26499
rect -17916 26496 -17913 26499
rect -17879 26494 -17876 26499
rect -17868 26494 -17866 26499
rect -17869 26480 -17866 26494
rect -17820 26479 -17818 26499
rect -17772 26496 -17770 26499
rect -17772 26479 -17769 26496
rect -17532 26479 -17530 26499
rect -17436 26479 -17434 26499
rect -17412 26479 -17410 26499
rect -17364 26479 -17362 26499
rect -17316 26479 -17314 26499
rect -17231 26494 -17228 26499
rect -17220 26494 -17218 26499
rect -17221 26480 -17218 26494
rect -17279 26479 -17221 26480
rect -17196 26479 -17194 26499
rect -17124 26496 -17122 26499
rect -17124 26479 -17121 26496
rect -17028 26479 -17026 26499
rect -16860 26479 -16858 26499
rect -16812 26479 -16810 26499
rect -16799 26494 -16796 26499
rect -16788 26494 -16786 26499
rect -16789 26480 -16786 26494
rect -16764 26479 -16762 26499
rect -16716 26479 -16714 26499
rect -16692 26496 -16690 26499
rect -16692 26479 -16689 26496
rect -16668 26479 -16666 26499
rect -16596 26479 -16594 26499
rect -16500 26479 -16498 26499
rect -16404 26479 -16402 26499
rect -16380 26479 -16378 26499
rect -16332 26496 -16330 26499
rect -16332 26479 -16329 26496
rect -16308 26479 -16306 26499
rect -16284 26479 -16282 26499
rect -16236 26479 -16234 26499
rect -16212 26479 -16210 26499
rect -16188 26479 -16186 26499
rect -15372 26479 -15370 26499
rect -15300 26479 -15298 26499
rect -15263 26479 -15229 26480
rect -15084 26479 -15082 26499
rect -15036 26479 -15034 26499
rect -14868 26479 -14866 26499
rect -14724 26479 -14722 26499
rect -14652 26479 -14650 26499
rect -14625 26496 -14611 26499
rect -14604 26496 -14601 26499
rect -14508 26479 -14506 26499
rect -14436 26479 -14434 26499
rect -14388 26479 -14386 26499
rect -14268 26479 -14266 26499
rect -14172 26479 -14170 26499
rect -14076 26479 -14074 26499
rect -14028 26479 -14026 26499
rect -13980 26479 -13978 26499
rect -13956 26479 -13954 26499
rect -13932 26479 -13930 26499
rect -13860 26479 -13858 26499
rect -13764 26479 -13762 26499
rect -13716 26479 -13714 26499
rect -13644 26479 -13642 26499
rect -13596 26479 -13594 26499
rect -13500 26479 -13498 26499
rect -13404 26479 -13402 26499
rect -13356 26479 -13354 26499
rect -13284 26479 -13282 26499
rect -12828 26479 -12826 26499
rect -12780 26479 -12778 26499
rect -12684 26479 -12682 26499
rect -12660 26479 -12658 26499
rect -12623 26494 -12620 26499
rect -12612 26494 -12610 26499
rect -12613 26480 -12610 26494
rect -12588 26479 -12586 26499
rect -12564 26479 -12562 26499
rect -12492 26479 -12490 26499
rect -12396 26479 -12394 26499
rect -12348 26479 -12346 26499
rect -12276 26479 -12274 26499
rect -12252 26479 -12250 26499
rect -12249 26496 -12235 26499
rect -12228 26496 -12225 26499
rect -12156 26479 -12154 26499
rect -12060 26479 -12058 26499
rect -12012 26479 -12010 26499
rect -11916 26479 -11914 26499
rect -11892 26479 -11890 26499
rect -11844 26479 -11842 26499
rect -11796 26479 -11794 26499
rect -11676 26479 -11674 26499
rect -11580 26479 -11578 26499
rect -11556 26479 -11554 26499
rect -11484 26479 -11482 26499
rect -11460 26479 -11458 26499
rect -11436 26479 -11434 26499
rect -11388 26479 -11386 26499
rect -11364 26479 -11362 26499
rect -11340 26479 -11338 26499
rect -11268 26479 -11266 26499
rect -11172 26479 -11170 26499
rect -11124 26479 -11122 26499
rect -11076 26479 -11074 26499
rect -11028 26479 -11026 26499
rect -10788 26479 -10786 26499
rect -10668 26479 -10666 26499
rect -9876 26479 -9874 26499
rect -9828 26479 -9826 26499
rect -9732 26479 -9730 26499
rect -9708 26479 -9706 26499
rect -9612 26479 -9610 26499
rect -9516 26479 -9514 26499
rect -9468 26479 -9466 26499
rect -9420 26479 -9418 26499
rect -9396 26479 -9394 26499
rect -9372 26479 -9370 26499
rect -9300 26479 -9298 26499
rect -9252 26479 -9250 26499
rect -9132 26479 -9130 26499
rect -9084 26479 -9082 26499
rect -9036 26479 -9034 26499
rect -8988 26479 -8986 26499
rect -8985 26496 -8971 26499
rect -8940 26479 -8938 26499
rect -8892 26479 -8890 26499
rect -8844 26479 -8842 26499
rect -8796 26479 -8794 26499
rect -8700 26479 -8698 26499
rect -8604 26479 -8602 26499
rect -8508 26479 -8506 26499
rect -8484 26479 -8482 26499
rect -8423 26494 -8420 26499
rect -8412 26494 -8410 26499
rect -8413 26480 -8410 26494
rect -8388 26479 -8386 26499
rect -8364 26479 -8362 26499
rect -8316 26496 -8314 26499
rect -8316 26479 -8313 26496
rect -8292 26479 -8290 26499
rect -8268 26479 -8266 26499
rect -8196 26479 -8194 26499
rect -8100 26479 -8098 26499
rect -8052 26479 -8050 26499
rect -7932 26479 -7930 26499
rect -7836 26479 -7834 26499
rect -7740 26479 -7738 26499
rect -7692 26479 -7690 26499
rect -7620 26479 -7618 26499
rect -7356 26479 -7354 26499
rect -7284 26479 -7282 26499
rect -7212 26479 -7210 26499
rect -7188 26479 -7186 26499
rect -7116 26479 -7114 26499
rect -7068 26479 -7066 26499
rect -6972 26479 -6970 26499
rect -6948 26479 -6946 26499
rect -6876 26479 -6874 26499
rect -6852 26479 -6850 26499
rect -6804 26479 -6802 26499
rect -6780 26479 -6778 26499
rect -6756 26479 -6754 26499
rect -6708 26479 -6706 26499
rect -6684 26479 -6682 26499
rect -6660 26479 -6658 26499
rect -6612 26479 -6610 26499
rect -6588 26479 -6586 26499
rect -6564 26479 -6562 26499
rect -6516 26479 -6514 26499
rect -6492 26479 -6490 26499
rect -6468 26479 -6466 26499
rect -6420 26479 -6418 26499
rect -6396 26479 -6394 26499
rect -6372 26479 -6370 26499
rect -6324 26479 -6322 26499
rect -6300 26479 -6298 26499
rect -6276 26479 -6274 26499
rect -6228 26479 -6226 26499
rect -6180 26479 -6178 26499
rect -6060 26479 -6058 26499
rect -5964 26479 -5962 26499
rect -5940 26479 -5938 26499
rect -5868 26479 -5866 26499
rect -5652 26479 -5650 26499
rect -5316 26479 -5314 26499
rect -5268 26479 -5266 26499
rect -5196 26479 -5194 26499
rect -5172 26479 -5170 26499
rect -5100 26479 -5098 26499
rect -5076 26479 -5074 26499
rect -4980 26479 -4978 26499
rect -4956 26479 -4954 26499
rect -4884 26479 -4882 26499
rect -4860 26479 -4858 26499
rect -4788 26479 -4786 26499
rect -4692 26479 -4690 26499
rect -4644 26479 -4642 26499
rect -4596 26479 -4594 26499
rect -4548 26479 -4546 26499
rect -4428 26479 -4426 26499
rect -4332 26479 -4330 26499
rect -4308 26479 -4306 26499
rect -4260 26479 -4258 26499
rect -4212 26479 -4210 26499
rect -4116 26479 -4114 26499
rect -4092 26479 -4090 26499
rect -4020 26479 -4018 26499
rect -3876 26479 -3874 26499
rect -3732 26479 -3730 26499
rect -3729 26496 -3715 26499
rect -3588 26479 -3586 26499
rect -3564 26479 -3562 26499
rect -3516 26479 -3514 26499
rect -3492 26479 -3490 26499
rect -3468 26479 -3466 26499
rect -3420 26479 -3418 26499
rect -3252 26479 -3250 26499
rect -3156 26479 -3154 26499
rect -3132 26479 -3130 26499
rect -3060 26479 -3058 26499
rect -3012 26479 -3010 26499
rect -2975 26494 -2972 26499
rect -2965 26480 -2962 26494
rect -2964 26479 -2962 26480
rect -2916 26479 -2914 26499
rect -2892 26479 -2890 26499
rect -2844 26496 -2842 26499
rect -2844 26479 -2841 26496
rect -2820 26479 -2818 26499
rect -2796 26479 -2794 26499
rect -2748 26479 -2746 26499
rect -2700 26479 -2698 26499
rect -2604 26479 -2602 26499
rect -2580 26479 -2578 26499
rect -2364 26479 -2362 26499
rect -2292 26479 -2290 26499
rect -2268 26479 -2266 26499
rect -2244 26479 -2242 26499
rect -2172 26479 -2170 26499
rect -2148 26479 -2146 26499
rect -2076 26479 -2074 26499
rect -2052 26479 -2050 26499
rect -1980 26479 -1978 26499
rect -1884 26479 -1882 26499
rect -1836 26479 -1834 26499
rect -1716 26479 -1714 26499
rect -1596 26479 -1594 26499
rect -1476 26479 -1474 26499
rect -1380 26479 -1378 26499
rect -1356 26479 -1354 26499
rect -1308 26479 -1306 26499
rect -1260 26479 -1258 26499
rect -1140 26479 -1138 26499
rect -852 26479 -850 26499
rect -804 26479 -802 26499
rect -756 26479 -754 26499
rect -708 26479 -706 26499
rect -612 26479 -610 26499
rect -588 26479 -586 26499
rect -540 26479 -538 26499
rect -516 26479 -514 26499
rect -492 26479 -490 26499
rect -444 26479 -442 26499
rect -396 26479 -394 26499
rect -300 26479 -298 26499
rect -276 26479 -274 26499
rect -204 26479 -202 26499
rect -108 26479 -106 26499
rect 12 26479 14 26499
rect 108 26479 110 26499
rect 156 26479 158 26499
rect 204 26479 206 26499
rect 228 26479 230 26499
rect 252 26479 254 26499
rect 348 26479 350 26499
rect 468 26479 470 26499
rect 564 26479 566 26499
rect 588 26479 590 26499
rect 636 26479 638 26499
rect 660 26479 662 26499
rect 684 26479 686 26499
rect 732 26479 734 26499
rect 756 26479 758 26499
rect 780 26479 782 26499
rect 876 26479 878 26499
rect 972 26479 974 26499
rect 1020 26479 1022 26499
rect 1068 26479 1070 26499
rect 1092 26479 1094 26499
rect 1116 26479 1118 26499
rect 1164 26479 1166 26499
rect 1212 26479 1214 26499
rect 1308 26479 1310 26499
rect 1332 26479 1334 26499
rect 1380 26479 1382 26499
rect 1428 26479 1430 26499
rect 1524 26479 1526 26499
rect 1548 26479 1550 26499
rect 1596 26479 1598 26499
rect 1620 26479 1622 26499
rect 1644 26479 1646 26499
rect 1692 26479 1694 26499
rect 1716 26479 1718 26499
rect 1740 26479 1742 26499
rect 1788 26479 1790 26499
rect 1836 26479 1838 26499
rect 1884 26479 1886 26499
rect 1932 26479 1934 26499
rect 1980 26479 1982 26499
rect 2028 26479 2030 26499
rect 2076 26479 2078 26499
rect 2100 26479 2102 26499
rect 2124 26479 2126 26499
rect 2172 26479 2174 26499
rect 2196 26479 2198 26499
rect 2220 26479 2222 26499
rect 2268 26479 2270 26499
rect 2292 26479 2294 26499
rect 2316 26479 2318 26499
rect 2364 26479 2366 26499
rect 2412 26479 2414 26499
rect 2460 26479 2462 26499
rect 2508 26479 2510 26499
rect 2556 26479 2558 26499
rect 2580 26479 2582 26499
rect 2604 26479 2606 26499
rect 2652 26479 2654 26499
rect 2676 26479 2678 26499
rect 2700 26479 2702 26499
rect 2748 26479 2750 26499
rect 2772 26479 2774 26499
rect 2796 26479 2798 26499
rect 2844 26479 2846 26499
rect 2868 26479 2870 26499
rect 2892 26479 2894 26499
rect 2940 26479 2942 26499
rect 3012 26479 3014 26499
rect 3108 26479 3110 26499
rect 3156 26479 3158 26499
rect 3252 26479 3254 26499
rect 3348 26479 3350 26499
rect 3396 26479 3398 26499
rect 3468 26479 3470 26499
rect 3492 26479 3494 26499
rect 3588 26479 3590 26499
rect 3612 26479 3614 26499
rect 3636 26479 3638 26499
rect 3708 26479 3710 26499
rect 3732 26479 3734 26499
rect 3745 26494 3748 26499
rect 3756 26494 3758 26499
rect 3755 26480 3758 26494
rect 3804 26479 3806 26499
rect 3828 26479 3830 26499
rect 3841 26494 3844 26499
rect 3852 26496 3854 26499
rect 3852 26494 3855 26496
rect 3851 26480 3855 26494
rect 3924 26479 3926 26499
rect 3948 26496 3950 26499
rect 3948 26479 3951 26496
rect 4020 26479 4022 26499
rect 4044 26479 4046 26499
rect 4092 26479 4094 26499
rect 4116 26479 4118 26499
rect 4140 26479 4142 26499
rect 4188 26479 4190 26499
rect 4212 26479 4214 26499
rect 4236 26479 4238 26499
rect 4308 26479 4310 26499
rect 4332 26479 4334 26499
rect 4404 26479 4406 26499
rect 4417 26494 4420 26499
rect 4428 26494 4430 26499
rect 4427 26480 4430 26494
rect 4500 26479 4502 26499
rect 4524 26496 4526 26499
rect 4524 26479 4527 26496
rect 4596 26479 4598 26499
rect 4860 26479 4862 26499
rect 4956 26479 4958 26499
rect 4980 26479 4982 26499
rect 5004 26479 5006 26499
rect 5076 26479 5078 26499
rect 5100 26479 5102 26499
rect 5124 26479 5126 26499
rect 5172 26479 5174 26499
rect 5196 26479 5198 26499
rect 5220 26479 5222 26499
rect 5268 26479 5270 26499
rect 5292 26479 5294 26499
rect 5388 26479 5390 26499
rect 5484 26479 5486 26499
rect 5508 26479 5510 26499
rect 5532 26479 5534 26499
rect 5580 26479 5582 26499
rect 5628 26479 5630 26499
rect 5724 26479 5726 26499
rect 5748 26479 5750 26499
rect 5796 26479 5798 26499
rect 5820 26479 5822 26499
rect 5844 26479 5846 26499
rect 5916 26480 5918 26499
rect 5881 26479 5939 26480
rect 6132 26479 6134 26499
rect 6180 26479 6182 26499
rect 6228 26479 6230 26499
rect 6252 26479 6254 26499
rect 6276 26479 6278 26499
rect 6324 26479 6326 26499
rect 6372 26479 6374 26499
rect 6492 26479 6494 26499
rect 6588 26479 6590 26499
rect 6612 26479 6614 26499
rect 6660 26479 6662 26499
rect 6684 26479 6686 26499
rect 6708 26479 6710 26499
rect 6780 26479 6782 26499
rect 6804 26479 6806 26499
rect 6828 26479 6830 26499
rect 6900 26479 6902 26499
rect 6924 26479 6926 26499
rect 7020 26479 7022 26499
rect 7140 26479 7142 26499
rect 7236 26479 7238 26499
rect 7249 26494 7252 26499
rect 7260 26494 7262 26499
rect 7259 26480 7262 26494
rect 7332 26479 7334 26499
rect 7356 26496 7358 26499
rect 7356 26479 7359 26496
rect 7380 26479 7382 26499
rect 7428 26479 7430 26499
rect 7452 26479 7454 26499
rect 7476 26479 7478 26499
rect 7524 26479 7526 26499
rect 7548 26479 7550 26499
rect 7572 26479 7574 26499
rect 7620 26479 7622 26499
rect 7644 26479 7646 26499
rect 7668 26479 7670 26499
rect 7716 26479 7718 26499
rect 7740 26479 7742 26499
rect 7753 26494 7756 26499
rect 7764 26494 7766 26499
rect 7763 26480 7766 26494
rect 7836 26479 7838 26499
rect 7860 26496 7862 26499
rect 7860 26479 7863 26496
rect 7884 26479 7886 26499
rect 7932 26479 7934 26499
rect 7956 26479 7958 26499
rect 7980 26479 7982 26499
rect 8052 26479 8054 26499
rect 8148 26479 8150 26499
rect 8196 26479 8198 26499
rect 8244 26479 8246 26499
rect 8268 26479 8270 26499
rect 8292 26479 8294 26499
rect 8340 26479 8342 26499
rect 8364 26479 8366 26499
rect 8388 26479 8390 26499
rect 8436 26479 8438 26499
rect 8460 26479 8462 26499
rect 8473 26494 8476 26499
rect 8484 26494 8486 26499
rect 8483 26480 8486 26494
rect 8556 26479 8558 26499
rect 8580 26496 8582 26499
rect 8580 26479 8583 26496
rect 8604 26479 8606 26499
rect 8676 26479 8678 26499
rect 8700 26479 8702 26499
rect 8724 26479 8726 26499
rect 8772 26479 8774 26499
rect 8820 26479 8822 26499
rect 8844 26479 8846 26499
rect 8868 26479 8870 26499
rect 9505 26494 9508 26499
rect 9515 26480 9518 26494
rect 9516 26479 9518 26480
rect 9612 26479 9615 26496
rect 9660 26479 9662 26499
rect 9684 26479 9686 26499
rect 9708 26479 9710 26499
rect 9756 26479 9758 26499
rect 9780 26479 9782 26499
rect 9804 26479 9806 26499
rect 9852 26479 9854 26499
rect 9876 26479 9878 26499
rect 9900 26479 9902 26499
rect 9948 26479 9950 26499
rect 9972 26479 9974 26499
rect 9996 26479 9998 26499
rect 10068 26479 10070 26499
rect 10092 26479 10094 26499
rect 10116 26479 10118 26499
rect 10164 26479 10166 26499
rect 10188 26479 10190 26499
rect 10212 26479 10214 26499
rect 10260 26479 10262 26499
rect 10284 26479 10286 26499
rect 10308 26479 10310 26499
rect 10380 26479 10382 26499
rect 10404 26479 10406 26499
rect 10428 26479 10430 26499
rect 10476 26479 10478 26499
rect 10500 26479 10502 26499
rect 10524 26479 10526 26499
rect 10572 26479 10574 26499
rect 10596 26479 10598 26499
rect 10620 26479 10622 26499
rect 10668 26479 10670 26499
rect 10692 26479 10694 26499
rect 10716 26479 10718 26499
rect 10788 26479 10790 26499
rect 10836 26479 10838 26499
rect 10956 26479 10958 26499
rect 11052 26479 11054 26499
rect 11076 26479 11078 26499
rect 11124 26479 11126 26499
rect 11172 26479 11174 26499
rect 11220 26479 11222 26499
rect 11340 26479 11342 26499
rect 11436 26479 11438 26499
rect 11532 26479 11534 26499
rect 11580 26479 11582 26499
rect 11628 26479 11630 26499
rect 11676 26479 11678 26499
rect 11772 26479 11774 26499
rect 11796 26479 11798 26499
rect 11844 26479 11846 26499
rect 11892 26479 11894 26499
rect 11988 26479 11990 26499
rect 12084 26479 12086 26499
rect 12132 26479 12134 26499
rect 12145 26479 12179 26480
rect 12228 26479 12230 26499
rect 12252 26480 12254 26499
rect 12300 26480 12302 26499
rect 12241 26479 12323 26480
rect 12324 26479 12326 26499
rect 12348 26479 12350 26499
rect 12396 26479 12398 26499
rect 12420 26479 12422 26499
rect 12444 26479 12446 26499
rect 12492 26479 12494 26499
rect 12516 26479 12518 26499
rect 12540 26479 12542 26499
rect 12588 26479 12590 26499
rect 12636 26479 12638 26499
rect 12732 26479 12734 26499
rect 12756 26479 12758 26499
rect 12804 26479 12806 26499
rect 12828 26479 12830 26499
rect 12852 26479 12854 26499
rect 12900 26479 12902 26499
rect 12948 26479 12950 26499
rect 13044 26479 13046 26499
rect 13068 26479 13070 26499
rect 13116 26479 13118 26499
rect 13284 26479 13286 26499
rect 13332 26479 13334 26499
rect 13428 26479 13430 26499
rect 13524 26479 13526 26499
rect 13572 26479 13574 26499
rect 13644 26479 13646 26499
rect 13668 26479 13670 26499
rect 13764 26479 13766 26499
rect 13812 26479 13814 26499
rect 13860 26479 13862 26499
rect 13908 26479 13910 26499
rect 13956 26479 13958 26499
rect 14004 26479 14006 26499
rect 14100 26479 14102 26499
rect 14196 26479 14198 26499
rect 14244 26479 14246 26499
rect 14292 26479 14294 26499
rect 14295 26496 14309 26499
rect 15132 26479 15134 26499
rect 15228 26479 15230 26499
rect 15252 26479 15254 26499
rect 15300 26479 15302 26499
rect 15324 26479 15326 26499
rect 15396 26479 15398 26499
rect 15420 26479 15422 26499
rect 15492 26479 15494 26499
rect 15540 26479 15542 26499
rect 15636 26479 15638 26499
rect 15660 26479 15662 26499
rect 15708 26479 15710 26499
rect 15732 26479 15734 26499
rect 15756 26479 15758 26499
rect 15804 26479 15806 26499
rect 15828 26479 15830 26499
rect 15852 26479 15854 26499
rect 15900 26479 15902 26499
rect 15948 26479 15950 26499
rect 15996 26479 15998 26499
rect 16044 26479 16046 26499
rect 16092 26479 16094 26499
rect 16140 26479 16142 26499
rect 16236 26479 16238 26499
rect 16260 26479 16262 26499
rect 16308 26479 16310 26499
rect 16332 26479 16334 26499
rect 16356 26479 16358 26499
rect 16404 26479 16406 26499
rect 16452 26479 16454 26499
rect 16548 26479 16550 26499
rect 16572 26479 16574 26499
rect 16620 26479 16622 26499
rect 16668 26479 16670 26499
rect 16716 26479 16718 26499
rect 16764 26479 16766 26499
rect 16836 26479 16838 26499
rect 16884 26479 16886 26499
rect 16980 26479 16982 26499
rect 17004 26480 17006 26499
rect 16993 26479 17027 26480
rect 17052 26479 17054 26499
rect 17100 26479 17102 26499
rect 17196 26479 17198 26499
rect 17220 26479 17222 26499
rect 17292 26479 17294 26499
rect 17316 26479 17318 26499
rect 18084 26479 18086 26499
rect 18132 26479 18134 26499
rect 18231 26496 18245 26499
rect 18252 26496 18255 26499
rect 18396 26479 18398 26499
rect 18492 26479 18494 26499
rect 18516 26479 18518 26499
rect 18564 26479 18566 26499
rect 18612 26479 18614 26499
rect 18660 26479 18662 26499
rect 18663 26496 18677 26499
rect 18684 26496 18687 26499
rect 18708 26479 18710 26499
rect 18756 26479 18758 26499
rect 18804 26479 18806 26499
rect 18852 26479 18854 26499
rect 18900 26479 18902 26499
rect 18996 26479 18998 26499
rect 19020 26479 19022 26499
rect 19092 26479 19094 26499
rect 19116 26479 19118 26499
rect 19140 26479 19142 26499
rect 19188 26479 19190 26499
rect 19236 26479 19238 26499
rect 19332 26479 19334 26499
rect 19476 26479 19478 26499
rect 19620 26479 19622 26499
rect 19716 26479 19718 26499
rect 19788 26479 19790 26499
rect 19836 26479 19838 26499
rect 19860 26479 19862 26499
rect 19863 26496 19877 26499
rect 19884 26499 32123 26503
rect 19884 26496 19901 26499
rect 19884 26479 19886 26496
rect 19932 26479 19934 26499
rect 19956 26479 19958 26499
rect 19980 26479 19982 26499
rect 20028 26479 20030 26499
rect 20052 26479 20054 26499
rect 20076 26479 20078 26499
rect 20148 26479 20150 26499
rect 20172 26479 20174 26499
rect 20196 26479 20198 26499
rect 20268 26479 20270 26499
rect 20292 26479 20294 26499
rect 20388 26479 20390 26499
rect 20412 26479 20414 26499
rect 20508 26479 20510 26499
rect 20556 26479 20558 26499
rect 20604 26479 20606 26499
rect 20916 26479 20918 26499
rect 20964 26479 20966 26499
rect 21012 26479 21014 26499
rect 21060 26479 21062 26499
rect 21084 26479 21086 26499
rect 21108 26479 21110 26499
rect 21204 26479 21206 26499
rect 21300 26479 21302 26499
rect 21324 26479 21326 26499
rect 21444 26479 21446 26499
rect 21468 26479 21470 26499
rect 21564 26479 21566 26499
rect 21612 26479 21614 26499
rect 21684 26479 21686 26499
rect 21708 26479 21710 26499
rect 21804 26479 21806 26499
rect 21828 26479 21830 26499
rect 21924 26479 21926 26499
rect 21948 26479 21950 26499
rect 22044 26479 22046 26499
rect 22068 26479 22070 26499
rect 22188 26479 22190 26499
rect 22212 26479 22214 26499
rect 23004 26479 23006 26499
rect 23052 26479 23054 26499
rect 23076 26479 23078 26499
rect 23100 26479 23102 26499
rect 23148 26479 23150 26499
rect 23220 26479 23222 26499
rect 23244 26479 23246 26499
rect 23316 26479 23318 26499
rect 23340 26479 23342 26499
rect 23412 26479 23414 26499
rect 23556 26479 23558 26499
rect 23628 26479 23630 26499
rect 23652 26479 23654 26499
rect 23676 26479 23678 26499
rect 23724 26479 23726 26499
rect 23737 26494 23740 26499
rect 23748 26494 23750 26499
rect 23747 26480 23750 26494
rect 23772 26479 23774 26499
rect 23820 26479 23822 26499
rect 23868 26479 23870 26499
rect 23892 26480 23894 26499
rect 23881 26479 23915 26480
rect 23916 26479 23918 26499
rect 23988 26479 23990 26499
rect 24012 26479 24014 26499
rect 24084 26479 24086 26499
rect 24327 26496 24341 26499
rect 24372 26479 24374 26499
rect 24396 26479 24398 26499
rect 24492 26479 24494 26499
rect 24516 26479 24518 26499
rect 24588 26479 24590 26499
rect 24612 26479 24614 26499
rect 24708 26479 24710 26499
rect 24732 26479 24734 26499
rect 24756 26479 24758 26499
rect 24852 26479 24854 26499
rect 24876 26479 24878 26499
rect 24972 26479 24974 26499
rect 24996 26479 24998 26499
rect 25092 26479 25094 26499
rect 25260 26479 25262 26499
rect 25356 26479 25358 26499
rect 25380 26479 25382 26499
rect 25452 26479 25454 26499
rect 25476 26479 25478 26499
rect 25500 26479 25502 26499
rect 25572 26479 25574 26499
rect 25596 26479 25598 26499
rect 27060 26479 27062 26499
rect 27108 26479 27110 26499
rect 27180 26479 27182 26499
rect 27324 26479 27326 26499
rect 27396 26479 27398 26499
rect 27420 26479 27422 26499
rect 27540 26479 27542 26499
rect 27564 26479 27566 26499
rect 30636 26479 30638 26499
rect 30660 26479 30662 26499
rect 30780 26479 30782 26499
rect 30804 26479 30806 26499
rect 30924 26479 30926 26499
rect 30948 26479 30950 26499
rect 31068 26479 31070 26499
rect 31092 26479 31094 26499
rect 31188 26479 31190 26499
rect 31236 26479 31238 26499
rect 31897 26494 31900 26499
rect 31907 26480 31910 26494
rect 31908 26479 31910 26480
rect 32004 26479 32007 26496
rect 32076 26480 32078 26499
rect 32089 26494 32092 26499
rect 32100 26494 32102 26499
rect 32099 26480 32102 26494
rect 32065 26479 32099 26480
rect -18750 26475 -18019 26479
rect -18527 26470 -18524 26475
rect -18396 26472 -18394 26475
rect -18517 26456 -18514 26470
rect -18623 26455 -18589 26456
rect -18516 26455 -18514 26456
rect -18396 26455 -18393 26472
rect -18287 26455 -18229 26456
rect -18108 26455 -18106 26475
rect -18036 26455 -18034 26475
rect -18033 26472 -18019 26475
rect -18009 26475 -16363 26479
rect -18009 26472 -17995 26475
rect -17820 26455 -17818 26475
rect -17793 26472 -17779 26475
rect -17772 26472 -17769 26475
rect -17567 26455 -17533 26456
rect -18623 26451 -18427 26455
rect -18516 26448 -18514 26451
rect -18441 26448 -18427 26451
rect -18417 26451 -17533 26455
rect -18417 26448 -18403 26451
rect -18396 26448 -18393 26451
rect -18516 26432 -18513 26448
rect -18527 26431 -18493 26432
rect -18359 26431 -18301 26432
rect -18108 26431 -18106 26451
rect -18036 26431 -18034 26451
rect -17951 26431 -17893 26432
rect -17820 26431 -17818 26451
rect -17532 26431 -17530 26475
rect -17519 26455 -17485 26456
rect -17436 26455 -17434 26475
rect -17412 26455 -17410 26475
rect -17364 26456 -17362 26475
rect -17399 26455 -17341 26456
rect -17316 26455 -17314 26475
rect -17279 26470 -17276 26475
rect -17269 26456 -17266 26470
rect -17268 26455 -17266 26456
rect -17196 26455 -17194 26475
rect -17145 26472 -17131 26475
rect -17124 26472 -17121 26475
rect -17028 26455 -17026 26475
rect -16860 26455 -16858 26475
rect -16812 26455 -16810 26475
rect -16764 26455 -16762 26475
rect -16716 26455 -16714 26475
rect -16713 26472 -16699 26475
rect -16692 26472 -16689 26475
rect -16668 26455 -16666 26475
rect -16596 26455 -16594 26475
rect -16500 26455 -16498 26475
rect -16404 26455 -16402 26475
rect -16380 26455 -16378 26475
rect -16377 26472 -16363 26475
rect -16353 26475 -12547 26479
rect -16353 26472 -16339 26475
rect -16332 26472 -16329 26475
rect -16308 26455 -16306 26475
rect -16284 26455 -16282 26475
rect -16236 26455 -16234 26475
rect -16212 26455 -16210 26475
rect -16188 26455 -16186 26475
rect -15372 26455 -15370 26475
rect -15300 26455 -15298 26475
rect -15084 26455 -15082 26475
rect -15036 26455 -15034 26475
rect -14868 26455 -14866 26475
rect -14724 26455 -14722 26475
rect -14652 26455 -14650 26475
rect -14508 26455 -14506 26475
rect -14436 26455 -14434 26475
rect -14388 26455 -14386 26475
rect -14268 26455 -14266 26475
rect -14172 26455 -14170 26475
rect -14076 26455 -14074 26475
rect -14028 26455 -14026 26475
rect -13980 26455 -13978 26475
rect -13956 26455 -13954 26475
rect -13932 26455 -13930 26475
rect -13860 26455 -13858 26475
rect -13764 26455 -13762 26475
rect -13716 26455 -13714 26475
rect -13644 26455 -13642 26475
rect -13596 26455 -13594 26475
rect -13500 26455 -13498 26475
rect -13404 26455 -13402 26475
rect -13356 26455 -13354 26475
rect -13284 26455 -13282 26475
rect -12828 26455 -12826 26475
rect -12780 26455 -12778 26475
rect -12684 26456 -12682 26475
rect -12695 26455 -12661 26456
rect -12660 26455 -12658 26475
rect -12588 26455 -12586 26475
rect -12564 26455 -12562 26475
rect -12561 26472 -12547 26475
rect -12537 26475 -8347 26479
rect -12537 26472 -12523 26475
rect -12492 26455 -12490 26475
rect -12396 26455 -12394 26475
rect -12348 26455 -12346 26475
rect -12276 26455 -12274 26475
rect -12252 26455 -12250 26475
rect -12156 26455 -12154 26475
rect -12060 26455 -12058 26475
rect -12012 26455 -12010 26475
rect -11916 26455 -11914 26475
rect -11892 26455 -11890 26475
rect -11844 26455 -11842 26475
rect -11796 26455 -11794 26475
rect -11676 26455 -11674 26475
rect -11580 26455 -11578 26475
rect -11556 26455 -11554 26475
rect -11484 26455 -11482 26475
rect -11460 26455 -11458 26475
rect -11436 26455 -11434 26475
rect -11388 26455 -11386 26475
rect -11364 26455 -11362 26475
rect -11340 26455 -11338 26475
rect -11268 26455 -11266 26475
rect -11172 26455 -11170 26475
rect -11124 26455 -11122 26475
rect -11076 26455 -11074 26475
rect -11028 26455 -11026 26475
rect -10788 26455 -10786 26475
rect -10668 26455 -10666 26475
rect -9876 26455 -9874 26475
rect -9828 26455 -9826 26475
rect -9732 26455 -9730 26475
rect -9708 26455 -9706 26475
rect -9612 26455 -9610 26475
rect -9516 26455 -9514 26475
rect -9468 26455 -9466 26475
rect -9420 26455 -9418 26475
rect -9396 26455 -9394 26475
rect -9372 26455 -9370 26475
rect -9300 26455 -9298 26475
rect -9252 26455 -9250 26475
rect -9132 26455 -9130 26475
rect -9084 26455 -9082 26475
rect -9036 26455 -9034 26475
rect -8988 26455 -8986 26475
rect -8940 26455 -8938 26475
rect -8892 26455 -8890 26475
rect -8844 26455 -8842 26475
rect -8796 26455 -8794 26475
rect -8700 26455 -8698 26475
rect -8604 26455 -8602 26475
rect -8508 26455 -8506 26475
rect -8484 26455 -8482 26475
rect -8388 26455 -8386 26475
rect -8364 26455 -8362 26475
rect -8361 26472 -8347 26475
rect -8337 26475 -2875 26479
rect -8337 26472 -8323 26475
rect -8316 26472 -8313 26475
rect -8292 26455 -8290 26475
rect -8268 26455 -8266 26475
rect -8196 26455 -8194 26475
rect -8100 26455 -8098 26475
rect -8052 26455 -8050 26475
rect -7932 26455 -7930 26475
rect -7836 26455 -7834 26475
rect -7740 26455 -7738 26475
rect -7692 26455 -7690 26475
rect -7620 26455 -7618 26475
rect -7415 26455 -7357 26456
rect -7356 26455 -7354 26475
rect -7284 26455 -7282 26475
rect -7212 26455 -7210 26475
rect -7188 26455 -7186 26475
rect -7116 26455 -7114 26475
rect -7068 26455 -7066 26475
rect -6972 26455 -6970 26475
rect -6948 26455 -6946 26475
rect -6876 26455 -6874 26475
rect -6852 26455 -6850 26475
rect -6804 26455 -6802 26475
rect -6780 26455 -6778 26475
rect -6756 26455 -6754 26475
rect -6708 26455 -6706 26475
rect -6684 26455 -6682 26475
rect -6660 26455 -6658 26475
rect -6612 26455 -6610 26475
rect -6588 26455 -6586 26475
rect -6564 26455 -6562 26475
rect -6516 26455 -6514 26475
rect -6492 26455 -6490 26475
rect -6468 26455 -6466 26475
rect -6420 26455 -6418 26475
rect -6396 26455 -6394 26475
rect -6372 26455 -6370 26475
rect -6324 26455 -6322 26475
rect -6300 26455 -6298 26475
rect -6276 26455 -6274 26475
rect -6228 26455 -6226 26475
rect -6180 26455 -6178 26475
rect -6060 26455 -6058 26475
rect -5964 26455 -5962 26475
rect -5940 26455 -5938 26475
rect -5868 26455 -5866 26475
rect -5652 26455 -5650 26475
rect -5409 26472 -5395 26475
rect -5316 26455 -5314 26475
rect -5268 26455 -5266 26475
rect -5196 26455 -5194 26475
rect -5172 26455 -5170 26475
rect -5100 26455 -5098 26475
rect -5076 26455 -5074 26475
rect -4980 26455 -4978 26475
rect -4956 26455 -4954 26475
rect -4884 26455 -4882 26475
rect -4860 26455 -4858 26475
rect -4788 26455 -4786 26475
rect -4692 26455 -4690 26475
rect -4644 26455 -4642 26475
rect -4596 26455 -4594 26475
rect -4548 26455 -4546 26475
rect -4428 26455 -4426 26475
rect -4332 26455 -4330 26475
rect -4308 26455 -4306 26475
rect -4260 26455 -4258 26475
rect -4212 26455 -4210 26475
rect -4116 26455 -4114 26475
rect -4092 26455 -4090 26475
rect -4020 26455 -4018 26475
rect -3876 26455 -3874 26475
rect -3732 26455 -3730 26475
rect -3588 26455 -3586 26475
rect -3564 26455 -3562 26475
rect -3516 26455 -3514 26475
rect -3492 26455 -3490 26475
rect -3468 26455 -3466 26475
rect -3420 26455 -3418 26475
rect -3335 26455 -3277 26456
rect -3252 26455 -3250 26475
rect -3156 26455 -3154 26475
rect -3132 26455 -3130 26475
rect -3060 26455 -3058 26475
rect -3012 26455 -3010 26475
rect -2964 26455 -2962 26475
rect -2916 26455 -2914 26475
rect -2892 26455 -2890 26475
rect -2889 26472 -2875 26475
rect -2865 26475 -1003 26479
rect -2865 26472 -2851 26475
rect -2844 26472 -2841 26475
rect -2820 26455 -2818 26475
rect -2796 26455 -2794 26475
rect -2748 26455 -2746 26475
rect -2700 26455 -2698 26475
rect -2604 26455 -2602 26475
rect -2580 26455 -2578 26475
rect -2364 26455 -2362 26475
rect -2292 26455 -2290 26475
rect -2268 26455 -2266 26475
rect -2244 26455 -2242 26475
rect -2172 26455 -2170 26475
rect -2148 26455 -2146 26475
rect -2076 26455 -2074 26475
rect -2052 26455 -2050 26475
rect -1980 26455 -1978 26475
rect -1884 26455 -1882 26475
rect -1836 26455 -1834 26475
rect -1716 26455 -1714 26475
rect -1596 26455 -1594 26475
rect -1476 26455 -1474 26475
rect -1380 26455 -1378 26475
rect -1356 26455 -1354 26475
rect -1308 26455 -1306 26475
rect -1260 26455 -1258 26475
rect -1140 26455 -1138 26475
rect -1017 26472 -1003 26475
rect -993 26475 9605 26479
rect -993 26472 -979 26475
rect -852 26455 -850 26475
rect -804 26455 -802 26475
rect -756 26455 -754 26475
rect -708 26455 -706 26475
rect -612 26455 -610 26475
rect -588 26455 -586 26475
rect -540 26455 -538 26475
rect -516 26455 -514 26475
rect -492 26455 -490 26475
rect -444 26455 -442 26475
rect -396 26455 -394 26475
rect -300 26455 -298 26475
rect -276 26455 -274 26475
rect -204 26455 -202 26475
rect -108 26455 -106 26475
rect 12 26455 14 26475
rect 108 26455 110 26475
rect 156 26455 158 26475
rect 204 26455 206 26475
rect 228 26455 230 26475
rect 252 26455 254 26475
rect 348 26455 350 26475
rect 385 26455 443 26456
rect 468 26455 470 26475
rect 564 26455 566 26475
rect 588 26455 590 26475
rect 636 26455 638 26475
rect 660 26455 662 26475
rect 684 26455 686 26475
rect 732 26455 734 26475
rect 756 26455 758 26475
rect 780 26455 782 26475
rect 876 26455 878 26475
rect 972 26455 974 26475
rect 1020 26455 1022 26475
rect 1068 26455 1070 26475
rect 1092 26455 1094 26475
rect 1116 26455 1118 26475
rect 1164 26455 1166 26475
rect 1212 26455 1214 26475
rect 1308 26455 1310 26475
rect 1332 26455 1334 26475
rect 1380 26455 1382 26475
rect 1428 26455 1430 26475
rect 1524 26455 1526 26475
rect 1548 26455 1550 26475
rect 1596 26455 1598 26475
rect 1620 26455 1622 26475
rect 1644 26455 1646 26475
rect 1692 26455 1694 26475
rect 1716 26455 1718 26475
rect 1740 26455 1742 26475
rect 1788 26455 1790 26475
rect 1836 26455 1838 26475
rect 1884 26455 1886 26475
rect 1932 26455 1934 26475
rect 1980 26455 1982 26475
rect 2028 26455 2030 26475
rect 2076 26455 2078 26475
rect 2100 26455 2102 26475
rect 2124 26455 2126 26475
rect 2172 26455 2174 26475
rect 2196 26455 2198 26475
rect 2220 26455 2222 26475
rect 2268 26455 2270 26475
rect 2292 26455 2294 26475
rect 2316 26455 2318 26475
rect 2364 26455 2366 26475
rect 2412 26455 2414 26475
rect 2460 26455 2462 26475
rect 2508 26455 2510 26475
rect 2556 26455 2558 26475
rect 2580 26455 2582 26475
rect 2604 26455 2606 26475
rect 2652 26455 2654 26475
rect 2676 26455 2678 26475
rect 2700 26455 2702 26475
rect 2748 26455 2750 26475
rect 2772 26455 2774 26475
rect 2796 26455 2798 26475
rect 2844 26455 2846 26475
rect 2868 26455 2870 26475
rect 2892 26455 2894 26475
rect 2940 26455 2942 26475
rect 3012 26455 3014 26475
rect 3108 26455 3110 26475
rect 3156 26455 3158 26475
rect 3252 26455 3254 26475
rect 3348 26455 3350 26475
rect 3396 26455 3398 26475
rect 3468 26455 3470 26475
rect 3492 26455 3494 26475
rect 3588 26455 3590 26475
rect 3612 26455 3614 26475
rect 3636 26455 3638 26475
rect 3708 26455 3710 26475
rect 3732 26455 3734 26475
rect 3804 26455 3806 26475
rect 3828 26455 3830 26475
rect 3831 26472 3845 26475
rect 3924 26455 3926 26475
rect 3927 26472 3941 26475
rect 3948 26472 3951 26475
rect 4020 26455 4022 26475
rect 4044 26455 4046 26475
rect 4092 26455 4094 26475
rect 4116 26455 4118 26475
rect 4140 26455 4142 26475
rect 4188 26455 4190 26475
rect 4212 26455 4214 26475
rect 4236 26455 4238 26475
rect 4308 26455 4310 26475
rect 4332 26455 4334 26475
rect 4404 26455 4406 26475
rect 4500 26455 4502 26475
rect 4503 26472 4517 26475
rect 4524 26472 4527 26475
rect 4596 26455 4598 26475
rect 4860 26455 4862 26475
rect 4956 26455 4958 26475
rect 4980 26455 4982 26475
rect 5004 26455 5006 26475
rect 5076 26455 5078 26475
rect 5100 26455 5102 26475
rect 5124 26455 5126 26475
rect 5172 26455 5174 26475
rect 5196 26455 5198 26475
rect 5220 26455 5222 26475
rect 5268 26455 5270 26475
rect 5292 26455 5294 26475
rect 5388 26455 5390 26475
rect 5484 26455 5486 26475
rect 5508 26455 5510 26475
rect 5532 26455 5534 26475
rect 5580 26455 5582 26475
rect 5628 26455 5630 26475
rect 5724 26455 5726 26475
rect 5748 26455 5750 26475
rect 5796 26455 5798 26475
rect 5820 26455 5822 26475
rect 5844 26455 5846 26475
rect 5881 26470 5884 26475
rect 5905 26470 5908 26475
rect 5916 26470 5918 26475
rect 5891 26456 5894 26470
rect 5915 26456 5918 26470
rect 5892 26455 5894 26456
rect 6132 26455 6134 26475
rect 6180 26455 6182 26475
rect 6228 26455 6230 26475
rect 6252 26455 6254 26475
rect 6276 26455 6278 26475
rect 6324 26455 6326 26475
rect 6372 26455 6374 26475
rect 6492 26455 6494 26475
rect 6588 26455 6590 26475
rect 6612 26455 6614 26475
rect 6660 26455 6662 26475
rect 6684 26455 6686 26475
rect 6708 26455 6710 26475
rect 6780 26455 6782 26475
rect 6804 26455 6806 26475
rect 6828 26455 6830 26475
rect 6900 26455 6902 26475
rect 6924 26455 6926 26475
rect 7020 26455 7022 26475
rect 7140 26455 7142 26475
rect 7236 26455 7238 26475
rect 7332 26455 7334 26475
rect 7335 26472 7349 26475
rect 7356 26472 7359 26475
rect 7380 26455 7382 26475
rect 7428 26455 7430 26475
rect 7452 26455 7454 26475
rect 7476 26455 7478 26475
rect 7524 26455 7526 26475
rect 7548 26455 7550 26475
rect 7572 26455 7574 26475
rect 7620 26455 7622 26475
rect 7644 26455 7646 26475
rect 7668 26455 7670 26475
rect 7716 26455 7718 26475
rect 7740 26455 7742 26475
rect 7836 26455 7838 26475
rect 7839 26472 7853 26475
rect 7860 26472 7863 26475
rect 7884 26455 7886 26475
rect 7932 26455 7934 26475
rect 7956 26455 7958 26475
rect 7980 26455 7982 26475
rect 8052 26455 8054 26475
rect 8148 26455 8150 26475
rect 8196 26455 8198 26475
rect 8244 26455 8246 26475
rect 8268 26455 8270 26475
rect 8292 26455 8294 26475
rect 8340 26455 8342 26475
rect 8364 26455 8366 26475
rect 8388 26455 8390 26475
rect 8436 26455 8438 26475
rect 8460 26455 8462 26475
rect 8556 26455 8558 26475
rect 8559 26472 8573 26475
rect 8580 26472 8583 26475
rect 8604 26455 8606 26475
rect 8676 26456 8678 26475
rect 8641 26455 8699 26456
rect 8700 26455 8702 26475
rect 8724 26455 8726 26475
rect 8772 26455 8774 26475
rect 8820 26455 8822 26475
rect 8844 26455 8846 26475
rect 8868 26455 8870 26475
rect 9516 26455 9518 26475
rect 9591 26472 9605 26475
rect 9612 26475 31997 26479
rect 9612 26472 9629 26475
rect 9612 26455 9614 26472
rect 9660 26455 9662 26475
rect 9684 26455 9686 26475
rect 9708 26455 9710 26475
rect 9756 26455 9758 26475
rect 9780 26455 9782 26475
rect 9804 26455 9806 26475
rect 9852 26455 9854 26475
rect 9876 26455 9878 26475
rect 9900 26455 9902 26475
rect 9948 26455 9950 26475
rect 9972 26455 9974 26475
rect 9996 26455 9998 26475
rect 10068 26455 10070 26475
rect 10092 26455 10094 26475
rect 10116 26455 10118 26475
rect 10164 26455 10166 26475
rect 10188 26455 10190 26475
rect 10212 26455 10214 26475
rect 10260 26455 10262 26475
rect 10284 26455 10286 26475
rect 10308 26455 10310 26475
rect 10380 26455 10382 26475
rect 10404 26455 10406 26475
rect 10428 26455 10430 26475
rect 10476 26455 10478 26475
rect 10500 26455 10502 26475
rect 10524 26455 10526 26475
rect 10572 26455 10574 26475
rect 10596 26455 10598 26475
rect 10620 26455 10622 26475
rect 10668 26455 10670 26475
rect 10692 26455 10694 26475
rect 10716 26455 10718 26475
rect 10788 26455 10790 26475
rect 10836 26455 10838 26475
rect 10956 26455 10958 26475
rect 11052 26455 11054 26475
rect 11076 26455 11078 26475
rect 11124 26455 11126 26475
rect 11172 26455 11174 26475
rect 11220 26455 11222 26475
rect 11340 26455 11342 26475
rect 11436 26455 11438 26475
rect 11532 26455 11534 26475
rect 11580 26455 11582 26475
rect 11628 26455 11630 26475
rect 11676 26455 11678 26475
rect 11772 26455 11774 26475
rect 11796 26455 11798 26475
rect 11844 26455 11846 26475
rect 11892 26455 11894 26475
rect 11988 26455 11990 26475
rect 12084 26456 12086 26475
rect 12049 26455 12107 26456
rect 12132 26455 12134 26475
rect 12228 26455 12230 26475
rect 12241 26470 12244 26475
rect 12252 26472 12254 26475
rect 12252 26470 12255 26472
rect 12289 26470 12292 26475
rect 12300 26470 12302 26475
rect 12251 26456 12255 26470
rect 12299 26456 12302 26470
rect 12324 26455 12326 26475
rect 12348 26472 12350 26475
rect 12396 26472 12398 26475
rect 12348 26455 12351 26472
rect 12396 26455 12399 26472
rect 12420 26455 12422 26475
rect 12444 26455 12446 26475
rect 12492 26455 12494 26475
rect 12516 26455 12518 26475
rect 12540 26455 12542 26475
rect 12588 26455 12590 26475
rect 12636 26455 12638 26475
rect 12732 26455 12734 26475
rect 12756 26455 12758 26475
rect 12804 26455 12806 26475
rect 12828 26455 12830 26475
rect 12852 26455 12854 26475
rect 12900 26455 12902 26475
rect 12948 26455 12950 26475
rect 13044 26455 13046 26475
rect 13068 26455 13070 26475
rect 13116 26455 13118 26475
rect 13284 26455 13286 26475
rect 13332 26455 13334 26475
rect 13428 26455 13430 26475
rect 13524 26455 13526 26475
rect 13572 26455 13574 26475
rect 13644 26455 13646 26475
rect 13668 26455 13670 26475
rect 13764 26455 13766 26475
rect 13812 26455 13814 26475
rect 13860 26455 13862 26475
rect 13908 26455 13910 26475
rect 13956 26455 13958 26475
rect 14004 26455 14006 26475
rect 14100 26455 14102 26475
rect 14196 26455 14198 26475
rect 14244 26455 14246 26475
rect 14292 26455 14294 26475
rect 15132 26455 15134 26475
rect 15228 26455 15230 26475
rect 15252 26455 15254 26475
rect 15300 26455 15302 26475
rect 15324 26455 15326 26475
rect 15396 26455 15398 26475
rect 15420 26455 15422 26475
rect 15492 26455 15494 26475
rect 15540 26455 15542 26475
rect 15636 26455 15638 26475
rect 15660 26455 15662 26475
rect 15708 26455 15710 26475
rect 15732 26455 15734 26475
rect 15756 26455 15758 26475
rect 15804 26455 15806 26475
rect 15828 26455 15830 26475
rect 15852 26455 15854 26475
rect 15900 26455 15902 26475
rect 15948 26455 15950 26475
rect 15996 26455 15998 26475
rect 16044 26455 16046 26475
rect 16092 26455 16094 26475
rect 16140 26455 16142 26475
rect 16236 26455 16238 26475
rect 16260 26455 16262 26475
rect 16308 26455 16310 26475
rect 16332 26455 16334 26475
rect 16356 26455 16358 26475
rect 16404 26455 16406 26475
rect 16452 26455 16454 26475
rect 16548 26455 16550 26475
rect 16572 26455 16574 26475
rect 16620 26455 16622 26475
rect 16668 26455 16670 26475
rect 16716 26455 16718 26475
rect 16764 26455 16766 26475
rect 16836 26455 16838 26475
rect 16884 26455 16886 26475
rect 16980 26455 16982 26475
rect 16993 26470 16996 26475
rect 17004 26470 17006 26475
rect 17003 26456 17006 26470
rect 17052 26455 17054 26475
rect 17100 26472 17102 26475
rect 17100 26455 17103 26472
rect 17196 26455 17198 26475
rect 17220 26455 17222 26475
rect 17292 26455 17294 26475
rect 17316 26455 17318 26475
rect 18084 26455 18086 26475
rect 18132 26455 18134 26475
rect 18396 26455 18398 26475
rect 18492 26455 18494 26475
rect 18516 26455 18518 26475
rect 18564 26455 18566 26475
rect 18612 26455 18614 26475
rect 18660 26455 18662 26475
rect 18708 26455 18710 26475
rect 18756 26455 18758 26475
rect 18804 26455 18806 26475
rect 18852 26455 18854 26475
rect 18900 26455 18902 26475
rect 18996 26455 18998 26475
rect 19020 26455 19022 26475
rect 19092 26455 19094 26475
rect 19116 26455 19118 26475
rect 19140 26455 19142 26475
rect 19188 26455 19190 26475
rect 19236 26455 19238 26475
rect 19332 26455 19334 26475
rect 19476 26455 19478 26475
rect 19620 26455 19622 26475
rect 19716 26455 19718 26475
rect 19788 26455 19790 26475
rect 19836 26455 19838 26475
rect 19860 26455 19862 26475
rect 19884 26455 19886 26475
rect 19932 26455 19934 26475
rect 19956 26455 19958 26475
rect 19980 26455 19982 26475
rect 20028 26455 20030 26475
rect 20052 26455 20054 26475
rect 20076 26455 20078 26475
rect 20148 26455 20150 26475
rect 20172 26455 20174 26475
rect 20196 26455 20198 26475
rect 20268 26455 20270 26475
rect 20292 26455 20294 26475
rect 20388 26455 20390 26475
rect 20412 26455 20414 26475
rect 20508 26455 20510 26475
rect 20556 26455 20558 26475
rect 20604 26455 20606 26475
rect 20916 26455 20918 26475
rect 20964 26455 20966 26475
rect 21012 26455 21014 26475
rect 21060 26455 21062 26475
rect 21084 26455 21086 26475
rect 21108 26455 21110 26475
rect 21204 26455 21206 26475
rect 21300 26455 21302 26475
rect 21324 26455 21326 26475
rect 21444 26455 21446 26475
rect 21468 26455 21470 26475
rect 21564 26455 21566 26475
rect 21612 26455 21614 26475
rect 21684 26455 21686 26475
rect 21708 26455 21710 26475
rect 21804 26455 21806 26475
rect 21828 26455 21830 26475
rect 21924 26455 21926 26475
rect 21948 26455 21950 26475
rect 22044 26455 22046 26475
rect 22068 26455 22070 26475
rect 22188 26455 22190 26475
rect 22212 26455 22214 26475
rect 23004 26455 23006 26475
rect 23052 26455 23054 26475
rect 23076 26455 23078 26475
rect 23100 26455 23102 26475
rect 23148 26455 23150 26475
rect 23220 26455 23222 26475
rect 23244 26455 23246 26475
rect 23316 26455 23318 26475
rect 23340 26455 23342 26475
rect 23412 26455 23414 26475
rect 23556 26455 23558 26475
rect 23628 26455 23630 26475
rect 23652 26455 23654 26475
rect 23676 26455 23678 26475
rect 23724 26455 23726 26475
rect 23772 26455 23774 26475
rect 23820 26455 23822 26475
rect 23823 26472 23837 26475
rect 23868 26455 23870 26475
rect 23881 26470 23884 26475
rect 23892 26470 23894 26475
rect 23891 26456 23894 26470
rect 23916 26455 23918 26475
rect 23988 26472 23990 26475
rect 23988 26455 23991 26472
rect 24012 26455 24014 26475
rect 24084 26455 24086 26475
rect 24372 26455 24374 26475
rect 24396 26455 24398 26475
rect 24492 26455 24494 26475
rect 24516 26455 24518 26475
rect 24588 26455 24590 26475
rect 24612 26455 24614 26475
rect 24708 26455 24710 26475
rect 24732 26455 24734 26475
rect 24756 26455 24758 26475
rect 24852 26455 24854 26475
rect 24876 26455 24878 26475
rect 24972 26455 24974 26475
rect 24996 26455 24998 26475
rect 25092 26455 25094 26475
rect 25260 26455 25262 26475
rect 25356 26455 25358 26475
rect 25380 26455 25382 26475
rect 25452 26455 25454 26475
rect 25476 26455 25478 26475
rect 25500 26455 25502 26475
rect 25572 26455 25574 26475
rect 25596 26455 25598 26475
rect 27060 26455 27062 26475
rect 27108 26455 27110 26475
rect 27180 26455 27182 26475
rect 27324 26455 27326 26475
rect 27396 26455 27398 26475
rect 27420 26455 27422 26475
rect 27540 26455 27542 26475
rect 27564 26455 27566 26475
rect 30636 26455 30638 26475
rect 30660 26455 30662 26475
rect 30780 26455 30782 26475
rect 30804 26455 30806 26475
rect 30924 26455 30926 26475
rect 30948 26455 30950 26475
rect 31068 26455 31070 26475
rect 31092 26455 31094 26475
rect 31188 26456 31190 26475
rect 31153 26455 31211 26456
rect 31236 26455 31238 26475
rect 31908 26455 31910 26475
rect 31983 26472 31997 26475
rect 32004 26475 32099 26479
rect 32004 26472 32021 26475
rect 32004 26456 32006 26472
rect 32065 26470 32068 26475
rect 32076 26470 32078 26475
rect 32075 26456 32078 26470
rect 31993 26455 32027 26456
rect -17519 26451 -17179 26455
rect -18527 26427 -18187 26431
rect -18527 26424 -18523 26427
rect -18516 26424 -18513 26427
rect -18201 26424 -18187 26427
rect -18177 26427 -17467 26431
rect -18177 26424 -18163 26427
rect -18407 26407 -18373 26408
rect -18167 26407 -18109 26408
rect -18108 26407 -18106 26427
rect -18036 26407 -18034 26427
rect -17951 26422 -17948 26427
rect -17820 26424 -17818 26427
rect -17941 26408 -17938 26422
rect -17940 26407 -17938 26408
rect -17820 26407 -17817 26424
rect -17615 26407 -17557 26408
rect -17532 26407 -17530 26427
rect -17481 26424 -17467 26427
rect -17460 26424 -17457 26448
rect -17460 26407 -17458 26424
rect -17436 26407 -17434 26451
rect -17412 26448 -17410 26451
rect -17412 26431 -17409 26448
rect -17375 26446 -17372 26451
rect -17364 26446 -17362 26451
rect -17365 26432 -17362 26446
rect -17316 26431 -17314 26451
rect -17268 26448 -17266 26451
rect -17292 26431 -17289 26448
rect -17268 26431 -17265 26448
rect -17196 26431 -17194 26451
rect -17193 26448 -17179 26451
rect -17169 26451 5981 26455
rect -17169 26448 -17155 26451
rect -17087 26431 -17053 26432
rect -17028 26431 -17026 26451
rect -16860 26431 -16858 26451
rect -16812 26431 -16810 26451
rect -16764 26431 -16762 26451
rect -16716 26431 -16714 26451
rect -16668 26431 -16666 26451
rect -16596 26431 -16594 26451
rect -16500 26431 -16498 26451
rect -16404 26431 -16402 26451
rect -16380 26431 -16378 26451
rect -16308 26431 -16306 26451
rect -16284 26431 -16282 26451
rect -16236 26431 -16234 26451
rect -16212 26431 -16210 26451
rect -16188 26431 -16186 26451
rect -15372 26431 -15370 26451
rect -15300 26431 -15298 26451
rect -15177 26448 -15163 26451
rect -15084 26431 -15082 26451
rect -15036 26431 -15034 26451
rect -14868 26431 -14866 26451
rect -14783 26431 -14725 26432
rect -14724 26431 -14722 26451
rect -14652 26431 -14650 26451
rect -14508 26431 -14506 26451
rect -14436 26431 -14434 26451
rect -14388 26431 -14386 26451
rect -14268 26431 -14266 26451
rect -14172 26431 -14170 26451
rect -14076 26431 -14074 26451
rect -14028 26431 -14026 26451
rect -13980 26431 -13978 26451
rect -13956 26431 -13954 26451
rect -13932 26431 -13930 26451
rect -13860 26431 -13858 26451
rect -13764 26431 -13762 26451
rect -13716 26431 -13714 26451
rect -13644 26431 -13642 26451
rect -13596 26431 -13594 26451
rect -13500 26431 -13498 26451
rect -13404 26431 -13402 26451
rect -13356 26431 -13354 26451
rect -13284 26431 -13282 26451
rect -13079 26431 -13021 26432
rect -12828 26431 -12826 26451
rect -12780 26431 -12778 26451
rect -12695 26446 -12692 26451
rect -12684 26446 -12682 26451
rect -12685 26432 -12682 26446
rect -12660 26431 -12658 26451
rect -12588 26448 -12586 26451
rect -12588 26431 -12585 26448
rect -12564 26431 -12562 26451
rect -12492 26431 -12490 26451
rect -12396 26431 -12394 26451
rect -12348 26431 -12346 26451
rect -12276 26431 -12274 26451
rect -12252 26431 -12250 26451
rect -12156 26431 -12154 26451
rect -12060 26431 -12058 26451
rect -12012 26431 -12010 26451
rect -11916 26431 -11914 26451
rect -11892 26431 -11890 26451
rect -11844 26431 -11842 26451
rect -11796 26431 -11794 26451
rect -11676 26431 -11674 26451
rect -11580 26431 -11578 26451
rect -11556 26431 -11554 26451
rect -11484 26431 -11482 26451
rect -11460 26431 -11458 26451
rect -11436 26431 -11434 26451
rect -11388 26431 -11386 26451
rect -11364 26431 -11362 26451
rect -11340 26431 -11338 26451
rect -11268 26431 -11266 26451
rect -11172 26431 -11170 26451
rect -11124 26431 -11122 26451
rect -11076 26431 -11074 26451
rect -11028 26431 -11026 26451
rect -10788 26431 -10786 26451
rect -10668 26431 -10666 26451
rect -9876 26431 -9874 26451
rect -9828 26431 -9826 26451
rect -9732 26431 -9730 26451
rect -9708 26431 -9706 26451
rect -9612 26431 -9610 26451
rect -9516 26431 -9514 26451
rect -9468 26431 -9466 26451
rect -9420 26431 -9418 26451
rect -9396 26431 -9394 26451
rect -9372 26431 -9370 26451
rect -9300 26431 -9298 26451
rect -9252 26431 -9250 26451
rect -9132 26431 -9130 26451
rect -9084 26431 -9082 26451
rect -9036 26431 -9034 26451
rect -8988 26431 -8986 26451
rect -8940 26431 -8938 26451
rect -8892 26431 -8890 26451
rect -8844 26431 -8842 26451
rect -8796 26431 -8794 26451
rect -8700 26431 -8698 26451
rect -8604 26431 -8602 26451
rect -8508 26431 -8506 26451
rect -8484 26431 -8482 26451
rect -8388 26431 -8386 26451
rect -8364 26431 -8362 26451
rect -8351 26431 -8293 26432
rect -8292 26431 -8290 26451
rect -8268 26431 -8266 26451
rect -8196 26431 -8194 26451
rect -8100 26431 -8098 26451
rect -8052 26431 -8050 26451
rect -7932 26431 -7930 26451
rect -7836 26431 -7834 26451
rect -7740 26431 -7738 26451
rect -7692 26431 -7690 26451
rect -7620 26431 -7618 26451
rect -7415 26446 -7412 26451
rect -7405 26432 -7402 26446
rect -7404 26431 -7402 26432
rect -7356 26431 -7354 26451
rect -7284 26448 -7282 26451
rect -7308 26431 -7305 26448
rect -7284 26431 -7281 26448
rect -7212 26431 -7210 26451
rect -7188 26431 -7186 26451
rect -7116 26431 -7114 26451
rect -7068 26431 -7066 26451
rect -6972 26431 -6970 26451
rect -6948 26431 -6946 26451
rect -6876 26431 -6874 26451
rect -6852 26431 -6850 26451
rect -6804 26431 -6802 26451
rect -6780 26431 -6778 26451
rect -6756 26431 -6754 26451
rect -6708 26431 -6706 26451
rect -6684 26431 -6682 26451
rect -6660 26431 -6658 26451
rect -6612 26431 -6610 26451
rect -6588 26431 -6586 26451
rect -6564 26431 -6562 26451
rect -6516 26431 -6514 26451
rect -6492 26431 -6490 26451
rect -6468 26431 -6466 26451
rect -6420 26431 -6418 26451
rect -6396 26431 -6394 26451
rect -6372 26431 -6370 26451
rect -6324 26431 -6322 26451
rect -6300 26431 -6298 26451
rect -6276 26431 -6274 26451
rect -6228 26431 -6226 26451
rect -6180 26431 -6178 26451
rect -6060 26431 -6058 26451
rect -5964 26431 -5962 26451
rect -5940 26431 -5938 26451
rect -5868 26431 -5866 26451
rect -5652 26431 -5650 26451
rect -5316 26431 -5314 26451
rect -5268 26431 -5266 26451
rect -5196 26431 -5194 26451
rect -5172 26431 -5170 26451
rect -5100 26431 -5098 26451
rect -5076 26431 -5074 26451
rect -4980 26431 -4978 26451
rect -4956 26431 -4954 26451
rect -4884 26431 -4882 26451
rect -4860 26431 -4858 26451
rect -4788 26431 -4786 26451
rect -4692 26431 -4690 26451
rect -4644 26431 -4642 26451
rect -4596 26431 -4594 26451
rect -4548 26431 -4546 26451
rect -4428 26431 -4426 26451
rect -4332 26431 -4330 26451
rect -4308 26431 -4306 26451
rect -4260 26431 -4258 26451
rect -4212 26431 -4210 26451
rect -4116 26431 -4114 26451
rect -4092 26431 -4090 26451
rect -4020 26431 -4018 26451
rect -3876 26431 -3874 26451
rect -3732 26431 -3730 26451
rect -3588 26431 -3586 26451
rect -3564 26431 -3562 26451
rect -3516 26431 -3514 26451
rect -3492 26431 -3490 26451
rect -3468 26431 -3466 26451
rect -3420 26431 -3418 26451
rect -3335 26446 -3332 26451
rect -3325 26432 -3322 26446
rect -3324 26431 -3322 26432
rect -3252 26431 -3250 26451
rect -3228 26431 -3225 26448
rect -3156 26431 -3154 26451
rect -3132 26431 -3130 26451
rect -3060 26431 -3058 26451
rect -3012 26431 -3010 26451
rect -2964 26431 -2962 26451
rect -2916 26431 -2914 26451
rect -2892 26431 -2890 26451
rect -2820 26431 -2818 26451
rect -2796 26431 -2794 26451
rect -2748 26431 -2746 26451
rect -2700 26431 -2698 26451
rect -2604 26431 -2602 26451
rect -2580 26431 -2578 26451
rect -2364 26431 -2362 26451
rect -2292 26431 -2290 26451
rect -2268 26431 -2266 26451
rect -2244 26431 -2242 26451
rect -2172 26431 -2170 26451
rect -2148 26431 -2146 26451
rect -2076 26431 -2074 26451
rect -2052 26431 -2050 26451
rect -1980 26431 -1978 26451
rect -1884 26431 -1882 26451
rect -1836 26431 -1834 26451
rect -1716 26431 -1714 26451
rect -1596 26431 -1594 26451
rect -1476 26431 -1474 26451
rect -1380 26431 -1378 26451
rect -1356 26431 -1354 26451
rect -1308 26431 -1306 26451
rect -1260 26431 -1258 26451
rect -1140 26431 -1138 26451
rect -852 26431 -850 26451
rect -804 26431 -802 26451
rect -756 26431 -754 26451
rect -708 26431 -706 26451
rect -612 26431 -610 26451
rect -588 26431 -586 26451
rect -540 26431 -538 26451
rect -516 26431 -514 26451
rect -492 26431 -490 26451
rect -444 26431 -442 26451
rect -396 26431 -394 26451
rect -300 26431 -298 26451
rect -276 26431 -274 26451
rect -204 26431 -202 26451
rect -108 26431 -106 26451
rect 12 26431 14 26451
rect 108 26431 110 26451
rect 156 26431 158 26451
rect 204 26431 206 26451
rect 228 26431 230 26451
rect 252 26431 254 26451
rect 348 26431 350 26451
rect 468 26431 470 26451
rect 492 26431 495 26448
rect 564 26431 566 26451
rect 588 26431 590 26451
rect 636 26431 638 26451
rect 660 26431 662 26451
rect 684 26431 686 26451
rect 732 26431 734 26451
rect 756 26431 758 26451
rect 780 26431 782 26451
rect 876 26431 878 26451
rect 972 26431 974 26451
rect 1020 26431 1022 26451
rect 1068 26431 1070 26451
rect 1092 26431 1094 26451
rect 1116 26431 1118 26451
rect 1164 26431 1166 26451
rect 1212 26431 1214 26451
rect 1308 26431 1310 26451
rect 1332 26431 1334 26451
rect 1380 26431 1382 26451
rect 1428 26431 1430 26451
rect 1524 26431 1526 26451
rect 1548 26431 1550 26451
rect 1596 26431 1598 26451
rect 1620 26431 1622 26451
rect 1644 26431 1646 26451
rect 1692 26431 1694 26451
rect 1716 26431 1718 26451
rect 1740 26431 1742 26451
rect 1788 26431 1790 26451
rect 1836 26431 1838 26451
rect 1884 26431 1886 26451
rect 1932 26431 1934 26451
rect 1980 26431 1982 26451
rect 2028 26431 2030 26451
rect 2076 26431 2078 26451
rect 2100 26431 2102 26451
rect 2124 26431 2126 26451
rect 2172 26431 2174 26451
rect 2196 26431 2198 26451
rect 2220 26431 2222 26451
rect 2268 26431 2270 26451
rect 2292 26431 2294 26451
rect 2316 26431 2318 26451
rect 2364 26431 2366 26451
rect 2412 26431 2414 26451
rect 2460 26431 2462 26451
rect 2508 26431 2510 26451
rect 2556 26431 2558 26451
rect 2580 26431 2582 26451
rect 2604 26431 2606 26451
rect 2652 26431 2654 26451
rect 2676 26431 2678 26451
rect 2700 26431 2702 26451
rect 2748 26431 2750 26451
rect 2772 26431 2774 26451
rect 2796 26431 2798 26451
rect 2844 26431 2846 26451
rect 2868 26431 2870 26451
rect 2892 26431 2894 26451
rect 2940 26431 2942 26451
rect 3012 26431 3014 26451
rect 3108 26431 3110 26451
rect 3156 26431 3158 26451
rect 3252 26431 3254 26451
rect 3348 26431 3350 26451
rect 3396 26431 3398 26451
rect 3468 26431 3470 26451
rect 3492 26431 3494 26451
rect 3588 26431 3590 26451
rect 3612 26431 3614 26451
rect 3636 26431 3638 26451
rect 3708 26431 3710 26451
rect 3732 26431 3734 26451
rect 3804 26431 3806 26451
rect 3828 26431 3830 26451
rect 3924 26431 3926 26451
rect 4020 26431 4022 26451
rect 4044 26431 4046 26451
rect 4092 26431 4094 26451
rect 4116 26431 4118 26451
rect 4140 26431 4142 26451
rect 4188 26431 4190 26451
rect 4212 26431 4214 26451
rect 4236 26431 4238 26451
rect 4308 26431 4310 26451
rect 4332 26431 4334 26451
rect 4404 26431 4406 26451
rect 4500 26431 4502 26451
rect 4596 26431 4598 26451
rect 4860 26431 4862 26451
rect 4956 26431 4958 26451
rect 4980 26431 4982 26451
rect 5004 26431 5006 26451
rect 5076 26431 5078 26451
rect 5100 26431 5102 26451
rect 5124 26431 5126 26451
rect 5172 26431 5174 26451
rect 5196 26431 5198 26451
rect 5220 26431 5222 26451
rect 5268 26431 5270 26451
rect 5292 26431 5294 26451
rect 5388 26431 5390 26451
rect 5484 26431 5486 26451
rect 5508 26431 5510 26451
rect 5532 26431 5534 26451
rect 5580 26431 5582 26451
rect 5628 26431 5630 26451
rect 5724 26431 5726 26451
rect 5748 26431 5750 26451
rect 5796 26431 5798 26451
rect 5820 26431 5822 26451
rect 5844 26431 5846 26451
rect 5892 26431 5894 26451
rect 5967 26448 5981 26451
rect 5991 26451 12365 26455
rect 5991 26448 6005 26451
rect 6132 26431 6134 26451
rect 6180 26431 6182 26451
rect 6228 26431 6230 26451
rect 6252 26431 6254 26451
rect 6276 26431 6278 26451
rect 6324 26431 6326 26451
rect 6372 26431 6374 26451
rect 6492 26431 6494 26451
rect 6588 26431 6590 26451
rect 6612 26431 6614 26451
rect 6660 26431 6662 26451
rect 6684 26431 6686 26451
rect 6708 26431 6710 26451
rect 6780 26431 6782 26451
rect 6804 26431 6806 26451
rect 6828 26431 6830 26451
rect 6900 26431 6902 26451
rect 6924 26431 6926 26451
rect 7020 26431 7022 26451
rect 7140 26431 7142 26451
rect 7236 26431 7238 26451
rect 7332 26431 7334 26451
rect 7380 26431 7382 26451
rect 7428 26431 7430 26451
rect 7452 26431 7454 26451
rect 7476 26431 7478 26451
rect 7524 26431 7526 26451
rect 7548 26431 7550 26451
rect 7572 26431 7574 26451
rect 7620 26431 7622 26451
rect 7644 26431 7646 26451
rect 7668 26431 7670 26451
rect 7716 26431 7718 26451
rect 7740 26431 7742 26451
rect 7836 26431 7838 26451
rect 7884 26431 7886 26451
rect 7932 26431 7934 26451
rect 7956 26431 7958 26451
rect 7980 26431 7982 26451
rect 8052 26431 8054 26451
rect 8148 26431 8150 26451
rect 8196 26431 8198 26451
rect 8244 26431 8246 26451
rect 8268 26431 8270 26451
rect 8292 26431 8294 26451
rect 8340 26431 8342 26451
rect 8364 26431 8366 26451
rect 8388 26431 8390 26451
rect 8436 26431 8438 26451
rect 8460 26431 8462 26451
rect 8556 26431 8558 26451
rect 8604 26431 8606 26451
rect 8641 26446 8644 26451
rect 8665 26446 8668 26451
rect 8676 26446 8678 26451
rect 8651 26432 8654 26446
rect 8675 26432 8678 26446
rect 8652 26431 8654 26432
rect 8700 26431 8702 26451
rect 8724 26431 8726 26451
rect 8772 26448 8774 26451
rect 8748 26431 8751 26448
rect 8772 26431 8775 26448
rect 8820 26431 8822 26451
rect 8844 26431 8846 26451
rect 8868 26431 8870 26451
rect 9516 26431 9518 26451
rect 9612 26431 9614 26451
rect 9660 26431 9662 26451
rect 9684 26431 9686 26451
rect 9708 26431 9710 26451
rect 9756 26431 9758 26451
rect 9780 26431 9782 26451
rect 9804 26431 9806 26451
rect 9852 26431 9854 26451
rect 9876 26431 9878 26451
rect 9900 26431 9902 26451
rect 9948 26431 9950 26451
rect 9972 26431 9974 26451
rect 9996 26431 9998 26451
rect 10068 26431 10070 26451
rect 10092 26431 10094 26451
rect 10116 26431 10118 26451
rect 10164 26431 10166 26451
rect 10188 26431 10190 26451
rect 10212 26431 10214 26451
rect 10260 26431 10262 26451
rect 10284 26431 10286 26451
rect 10308 26431 10310 26451
rect 10380 26431 10382 26451
rect 10404 26431 10406 26451
rect 10428 26431 10430 26451
rect 10476 26431 10478 26451
rect 10500 26431 10502 26451
rect 10524 26431 10526 26451
rect 10572 26431 10574 26451
rect 10596 26431 10598 26451
rect 10620 26431 10622 26451
rect 10668 26431 10670 26451
rect 10692 26431 10694 26451
rect 10716 26431 10718 26451
rect 10788 26431 10790 26451
rect 10836 26431 10838 26451
rect 10956 26431 10958 26451
rect 11052 26431 11054 26451
rect 11076 26431 11078 26451
rect 11124 26431 11126 26451
rect 11172 26431 11174 26451
rect 11220 26431 11222 26451
rect 11340 26431 11342 26451
rect 11436 26431 11438 26451
rect 11532 26431 11534 26451
rect 11580 26431 11582 26451
rect 11628 26431 11630 26451
rect 11676 26431 11678 26451
rect 11772 26431 11774 26451
rect 11796 26431 11798 26451
rect 11844 26431 11846 26451
rect 11892 26431 11894 26451
rect 11988 26431 11990 26451
rect 12049 26446 12052 26451
rect 12073 26446 12076 26451
rect 12084 26446 12086 26451
rect 12059 26432 12062 26446
rect 12083 26432 12086 26446
rect 12060 26431 12062 26432
rect 12132 26431 12134 26451
rect 12228 26431 12230 26451
rect 12231 26448 12245 26451
rect 12324 26431 12326 26451
rect 12327 26448 12341 26451
rect 12348 26448 12365 26451
rect 12375 26451 32027 26455
rect 12375 26448 12389 26451
rect 12396 26448 12399 26451
rect 12420 26431 12422 26451
rect 12444 26431 12446 26451
rect 12492 26431 12494 26451
rect 12516 26431 12518 26451
rect 12540 26431 12542 26451
rect 12588 26431 12590 26451
rect 12636 26431 12638 26451
rect 12732 26431 12734 26451
rect 12756 26431 12758 26451
rect 12804 26431 12806 26451
rect 12828 26431 12830 26451
rect 12852 26431 12854 26451
rect 12900 26431 12902 26451
rect 12948 26431 12950 26451
rect 13044 26431 13046 26451
rect 13068 26431 13070 26451
rect 13116 26431 13118 26451
rect 13284 26431 13286 26451
rect 13332 26431 13334 26451
rect 13428 26431 13430 26451
rect 13524 26431 13526 26451
rect 13572 26431 13574 26451
rect 13644 26431 13646 26451
rect 13668 26431 13670 26451
rect 13764 26431 13766 26451
rect 13812 26431 13814 26451
rect 13860 26431 13862 26451
rect 13908 26431 13910 26451
rect 13956 26431 13958 26451
rect 14004 26431 14006 26451
rect 14100 26431 14102 26451
rect 14196 26431 14198 26451
rect 14244 26431 14246 26451
rect 14292 26431 14294 26451
rect 15132 26431 15134 26451
rect 15228 26431 15230 26451
rect 15252 26431 15254 26451
rect 15300 26431 15302 26451
rect 15324 26431 15326 26451
rect 15396 26431 15398 26451
rect 15420 26431 15422 26451
rect 15492 26431 15494 26451
rect 15540 26431 15542 26451
rect 15636 26431 15638 26451
rect 15660 26431 15662 26451
rect 15708 26431 15710 26451
rect 15732 26431 15734 26451
rect 15756 26431 15758 26451
rect 15804 26431 15806 26451
rect 15828 26431 15830 26451
rect 15852 26431 15854 26451
rect 15900 26431 15902 26451
rect 15948 26431 15950 26451
rect 15996 26431 15998 26451
rect 16044 26431 16046 26451
rect 16092 26431 16094 26451
rect 16140 26431 16142 26451
rect 16236 26431 16238 26451
rect 16260 26431 16262 26451
rect 16308 26431 16310 26451
rect 16332 26431 16334 26451
rect 16356 26431 16358 26451
rect 16404 26431 16406 26451
rect 16452 26431 16454 26451
rect 16548 26431 16550 26451
rect 16572 26431 16574 26451
rect 16620 26431 16622 26451
rect 16668 26431 16670 26451
rect 16716 26431 16718 26451
rect 16764 26431 16766 26451
rect 16836 26431 16838 26451
rect 16884 26431 16886 26451
rect 16980 26431 16982 26451
rect 17052 26431 17054 26451
rect 17079 26448 17093 26451
rect 17100 26448 17103 26451
rect 17196 26431 17198 26451
rect 17220 26431 17222 26451
rect 17292 26431 17294 26451
rect 17316 26431 17318 26451
rect 18084 26431 18086 26451
rect 18132 26431 18134 26451
rect 18396 26431 18398 26451
rect 18492 26431 18494 26451
rect 18516 26431 18518 26451
rect 18564 26431 18566 26451
rect 18612 26431 18614 26451
rect 18660 26431 18662 26451
rect 18708 26431 18710 26451
rect 18756 26431 18758 26451
rect 18804 26431 18806 26451
rect 18852 26431 18854 26451
rect 18900 26431 18902 26451
rect 18996 26431 18998 26451
rect 19020 26431 19022 26451
rect 19092 26431 19094 26451
rect 19116 26431 19118 26451
rect 19140 26431 19142 26451
rect 19188 26431 19190 26451
rect 19236 26431 19238 26451
rect 19332 26431 19334 26451
rect 19476 26431 19478 26451
rect 19620 26431 19622 26451
rect 19716 26431 19718 26451
rect 19788 26431 19790 26451
rect 19836 26431 19838 26451
rect 19860 26431 19862 26451
rect 19884 26431 19886 26451
rect 19932 26431 19934 26451
rect 19956 26431 19958 26451
rect 19980 26431 19982 26451
rect 20028 26431 20030 26451
rect 20052 26431 20054 26451
rect 20076 26431 20078 26451
rect 20148 26431 20150 26451
rect 20172 26431 20174 26451
rect 20196 26431 20198 26451
rect 20268 26431 20270 26451
rect 20292 26431 20294 26451
rect 20388 26431 20390 26451
rect 20412 26431 20414 26451
rect 20508 26431 20510 26451
rect 20556 26431 20558 26451
rect 20604 26431 20606 26451
rect 20916 26431 20918 26451
rect 20964 26431 20966 26451
rect 21012 26431 21014 26451
rect 21060 26431 21062 26451
rect 21084 26431 21086 26451
rect 21108 26431 21110 26451
rect 21204 26431 21206 26451
rect 21300 26431 21302 26451
rect 21324 26431 21326 26451
rect 21444 26431 21446 26451
rect 21468 26431 21470 26451
rect 21564 26431 21566 26451
rect 21612 26431 21614 26451
rect 21684 26431 21686 26451
rect 21708 26431 21710 26451
rect 21804 26431 21806 26451
rect 21828 26431 21830 26451
rect 21924 26431 21926 26451
rect 21948 26431 21950 26451
rect 22044 26431 22046 26451
rect 22068 26431 22070 26451
rect 22188 26431 22190 26451
rect 22212 26431 22214 26451
rect 23004 26431 23006 26451
rect 23052 26431 23054 26451
rect 23076 26431 23078 26451
rect 23100 26431 23102 26451
rect 23148 26431 23150 26451
rect 23220 26431 23222 26451
rect 23244 26431 23246 26451
rect 23316 26431 23318 26451
rect 23340 26431 23342 26451
rect 23412 26431 23414 26451
rect 23556 26431 23558 26451
rect 23628 26431 23630 26451
rect 23652 26431 23654 26451
rect 23676 26431 23678 26451
rect 23724 26431 23726 26451
rect 23772 26431 23774 26451
rect 23820 26431 23822 26451
rect 23868 26431 23870 26451
rect 23916 26431 23918 26451
rect 23967 26448 23981 26451
rect 23988 26448 23991 26451
rect 24012 26431 24014 26451
rect 24084 26431 24086 26451
rect 24372 26431 24374 26451
rect 24396 26431 24398 26451
rect 24492 26431 24494 26451
rect 24516 26431 24518 26451
rect 24588 26431 24590 26451
rect 24612 26431 24614 26451
rect 24708 26431 24710 26451
rect 24732 26431 24734 26451
rect 24756 26431 24758 26451
rect 24852 26431 24854 26451
rect 24876 26431 24878 26451
rect 24972 26431 24974 26451
rect 24996 26431 24998 26451
rect 25092 26431 25094 26451
rect 25260 26431 25262 26451
rect 25356 26431 25358 26451
rect 25380 26431 25382 26451
rect 25452 26431 25454 26451
rect 25476 26431 25478 26451
rect 25500 26431 25502 26451
rect 25572 26431 25574 26451
rect 25596 26431 25598 26451
rect 27060 26431 27062 26451
rect 27108 26431 27110 26451
rect 27180 26431 27182 26451
rect 27324 26431 27326 26451
rect 27396 26431 27398 26451
rect 27420 26431 27422 26451
rect 27540 26431 27542 26451
rect 27564 26431 27566 26451
rect 30457 26431 30515 26432
rect 30636 26431 30638 26451
rect 30660 26431 30662 26451
rect 30780 26431 30782 26451
rect 30804 26431 30806 26451
rect 30924 26431 30926 26451
rect 30948 26431 30950 26451
rect 31068 26431 31070 26451
rect 31092 26431 31094 26451
rect 31153 26446 31156 26451
rect 31177 26446 31180 26451
rect 31188 26446 31190 26451
rect 31163 26432 31166 26446
rect 31187 26432 31190 26446
rect 31164 26431 31166 26432
rect 31236 26431 31238 26451
rect 31908 26432 31910 26451
rect 31993 26446 31996 26451
rect 32004 26446 32006 26451
rect 32003 26432 32006 26446
rect 31801 26431 31835 26432
rect -17433 26427 -17299 26431
rect -17433 26424 -17419 26427
rect -17412 26424 -17409 26427
rect -17316 26407 -17314 26427
rect -17313 26424 -17299 26427
rect -17292 26427 -7315 26431
rect -17292 26424 -17275 26427
rect -17268 26424 -17265 26427
rect -17292 26407 -17290 26424
rect -17196 26407 -17194 26427
rect -17028 26407 -17026 26427
rect -16860 26407 -16858 26427
rect -16812 26407 -16810 26427
rect -16764 26407 -16762 26427
rect -16716 26407 -16714 26427
rect -16668 26407 -16666 26427
rect -16596 26407 -16594 26427
rect -16500 26407 -16498 26427
rect -16404 26407 -16402 26427
rect -16380 26407 -16378 26427
rect -16367 26407 -16333 26408
rect -18407 26403 -18259 26407
rect -18273 26400 -18259 26403
rect -18249 26403 -17851 26407
rect -18249 26400 -18235 26403
rect -18108 26383 -18106 26403
rect -18036 26400 -18034 26403
rect -18036 26383 -18033 26400
rect -17999 26383 -17941 26384
rect -17940 26383 -17938 26403
rect -17865 26400 -17851 26403
rect -17841 26403 -16333 26407
rect -17841 26400 -17827 26403
rect -17820 26400 -17817 26403
rect -17615 26398 -17612 26403
rect -17605 26384 -17602 26398
rect -17903 26383 -17869 26384
rect -17604 26383 -17602 26384
rect -17532 26383 -17530 26403
rect -17460 26383 -17458 26403
rect -17436 26383 -17434 26403
rect -17316 26384 -17314 26403
rect -17327 26383 -17293 26384
rect -17292 26383 -17290 26403
rect -17196 26383 -17194 26403
rect -17028 26383 -17026 26403
rect -17001 26400 -16987 26403
rect -16860 26383 -16858 26403
rect -16812 26383 -16810 26403
rect -16764 26383 -16762 26403
rect -16751 26383 -16717 26384
rect -18321 26379 -18067 26383
rect -18321 26376 -18307 26379
rect -18273 26359 -18253 26360
rect -18215 26359 -18181 26360
rect -18108 26359 -18106 26379
rect -18081 26376 -18067 26379
rect -18057 26379 -17515 26383
rect -18057 26376 -18043 26379
rect -18036 26376 -18033 26379
rect -17940 26359 -17938 26379
rect -17892 26374 -17889 26376
rect -17893 26366 -17889 26374
rect -17879 26366 -17875 26374
rect -17893 26360 -17879 26366
rect -17735 26359 -17677 26360
rect -17604 26359 -17602 26379
rect -17532 26359 -17530 26379
rect -17529 26376 -17515 26379
rect -17505 26379 -16717 26383
rect -17505 26376 -17491 26379
rect -17460 26359 -17458 26379
rect -17436 26359 -17434 26379
rect -17327 26374 -17324 26379
rect -17316 26374 -17314 26379
rect -17317 26360 -17314 26374
rect -17292 26359 -17290 26379
rect -17196 26359 -17194 26379
rect -17028 26359 -17026 26379
rect -16860 26359 -16858 26379
rect -16812 26360 -16810 26379
rect -16847 26359 -16789 26360
rect -16764 26359 -16762 26379
rect -16716 26359 -16714 26403
rect -16703 26383 -16669 26384
rect -16668 26383 -16666 26403
rect -16596 26383 -16594 26403
rect -16500 26383 -16498 26403
rect -16404 26384 -16402 26403
rect -16415 26383 -16381 26384
rect -16380 26383 -16378 26403
rect -16367 26398 -16364 26403
rect -16357 26384 -16354 26398
rect -16356 26383 -16354 26384
rect -16308 26383 -16306 26427
rect -16284 26408 -16282 26427
rect -16295 26407 -16261 26408
rect -16236 26407 -16234 26427
rect -16212 26407 -16210 26427
rect -16188 26407 -16186 26427
rect -15372 26408 -15370 26427
rect -15383 26407 -15349 26408
rect -15300 26407 -15298 26427
rect -15084 26407 -15082 26427
rect -15036 26407 -15034 26427
rect -14868 26407 -14866 26427
rect -14783 26422 -14780 26427
rect -14773 26408 -14770 26422
rect -14772 26407 -14770 26408
rect -14724 26407 -14722 26427
rect -14652 26424 -14650 26427
rect -14652 26407 -14649 26424
rect -14508 26407 -14506 26427
rect -14436 26407 -14434 26427
rect -14388 26407 -14386 26427
rect -14375 26407 -14341 26408
rect -14268 26407 -14266 26427
rect -14172 26407 -14170 26427
rect -14076 26407 -14074 26427
rect -14063 26407 -14029 26408
rect -14028 26407 -14026 26427
rect -13980 26407 -13978 26427
rect -13956 26407 -13954 26427
rect -13932 26407 -13930 26427
rect -13860 26407 -13858 26427
rect -13764 26407 -13762 26427
rect -13716 26407 -13714 26427
rect -13644 26407 -13642 26427
rect -13596 26407 -13594 26427
rect -13500 26407 -13498 26427
rect -13404 26407 -13402 26427
rect -13356 26407 -13354 26427
rect -13284 26407 -13282 26427
rect -13079 26422 -13076 26427
rect -13069 26408 -13066 26422
rect -13068 26407 -13066 26408
rect -12828 26407 -12826 26427
rect -12780 26407 -12778 26427
rect -12660 26407 -12658 26427
rect -12609 26424 -12595 26427
rect -12588 26424 -12585 26427
rect -12564 26407 -12562 26427
rect -12492 26407 -12490 26427
rect -12396 26407 -12394 26427
rect -12348 26407 -12346 26427
rect -12276 26407 -12274 26427
rect -12252 26407 -12250 26427
rect -12156 26407 -12154 26427
rect -12060 26407 -12058 26427
rect -12012 26407 -12010 26427
rect -11916 26407 -11914 26427
rect -11892 26407 -11890 26427
rect -11844 26407 -11842 26427
rect -11796 26407 -11794 26427
rect -11676 26407 -11674 26427
rect -11580 26407 -11578 26427
rect -11556 26407 -11554 26427
rect -11484 26407 -11482 26427
rect -11460 26407 -11458 26427
rect -11436 26407 -11434 26427
rect -11388 26407 -11386 26427
rect -11364 26407 -11362 26427
rect -11340 26407 -11338 26427
rect -11268 26407 -11266 26427
rect -11172 26407 -11170 26427
rect -11124 26407 -11122 26427
rect -11076 26407 -11074 26427
rect -11028 26407 -11026 26427
rect -10788 26407 -10786 26427
rect -10668 26407 -10666 26427
rect -9876 26407 -9874 26427
rect -9828 26407 -9826 26427
rect -9732 26407 -9730 26427
rect -9708 26407 -9706 26427
rect -9612 26407 -9610 26427
rect -9516 26407 -9514 26427
rect -9468 26407 -9466 26427
rect -9420 26407 -9418 26427
rect -9396 26407 -9394 26427
rect -9372 26407 -9370 26427
rect -9300 26407 -9298 26427
rect -9252 26407 -9250 26427
rect -9132 26407 -9130 26427
rect -9084 26407 -9082 26427
rect -9036 26407 -9034 26427
rect -8988 26407 -8986 26427
rect -8940 26407 -8938 26427
rect -8892 26407 -8890 26427
rect -8844 26407 -8842 26427
rect -8796 26407 -8794 26427
rect -8700 26407 -8698 26427
rect -8604 26407 -8602 26427
rect -8508 26407 -8506 26427
rect -8484 26407 -8482 26427
rect -8388 26407 -8386 26427
rect -8364 26407 -8362 26427
rect -8351 26422 -8348 26427
rect -8341 26408 -8338 26422
rect -8340 26407 -8338 26408
rect -8292 26407 -8290 26427
rect -8268 26407 -8266 26427
rect -8196 26407 -8194 26427
rect -8100 26407 -8098 26427
rect -8052 26407 -8050 26427
rect -7932 26407 -7930 26427
rect -7836 26407 -7834 26427
rect -7740 26407 -7738 26427
rect -7692 26407 -7690 26427
rect -7620 26407 -7618 26427
rect -7404 26407 -7402 26427
rect -7356 26407 -7354 26427
rect -7329 26424 -7315 26427
rect -7308 26427 -3235 26431
rect -7308 26424 -7291 26427
rect -7284 26424 -7281 26427
rect -7308 26407 -7306 26424
rect -7212 26407 -7210 26427
rect -7188 26407 -7186 26427
rect -7116 26407 -7114 26427
rect -7068 26407 -7066 26427
rect -6972 26407 -6970 26427
rect -6948 26407 -6946 26427
rect -6876 26407 -6874 26427
rect -6852 26407 -6850 26427
rect -6804 26407 -6802 26427
rect -6780 26407 -6778 26427
rect -6756 26407 -6754 26427
rect -6708 26407 -6706 26427
rect -6684 26407 -6682 26427
rect -6660 26407 -6658 26427
rect -6612 26407 -6610 26427
rect -6588 26407 -6586 26427
rect -6564 26407 -6562 26427
rect -6516 26407 -6514 26427
rect -6492 26407 -6490 26427
rect -6468 26407 -6466 26427
rect -6420 26407 -6418 26427
rect -6396 26407 -6394 26427
rect -6372 26407 -6370 26427
rect -6324 26407 -6322 26427
rect -6300 26407 -6298 26427
rect -6276 26407 -6274 26427
rect -6228 26407 -6226 26427
rect -6180 26407 -6178 26427
rect -6060 26407 -6058 26427
rect -5964 26407 -5962 26427
rect -5940 26407 -5938 26427
rect -5868 26407 -5866 26427
rect -5652 26407 -5650 26427
rect -5316 26407 -5314 26427
rect -5268 26407 -5266 26427
rect -5196 26407 -5194 26427
rect -5172 26407 -5170 26427
rect -5100 26407 -5098 26427
rect -5076 26407 -5074 26427
rect -4980 26407 -4978 26427
rect -4956 26407 -4954 26427
rect -4884 26407 -4882 26427
rect -4860 26407 -4858 26427
rect -4788 26407 -4786 26427
rect -4692 26407 -4690 26427
rect -4644 26407 -4642 26427
rect -4596 26407 -4594 26427
rect -4548 26407 -4546 26427
rect -4428 26407 -4426 26427
rect -4332 26407 -4330 26427
rect -4308 26407 -4306 26427
rect -4260 26407 -4258 26427
rect -4212 26407 -4210 26427
rect -4116 26407 -4114 26427
rect -4092 26407 -4090 26427
rect -4020 26407 -4018 26427
rect -3876 26407 -3874 26427
rect -3732 26407 -3730 26427
rect -3588 26407 -3586 26427
rect -3564 26407 -3562 26427
rect -3516 26407 -3514 26427
rect -3492 26407 -3490 26427
rect -3468 26407 -3466 26427
rect -3420 26407 -3418 26427
rect -3324 26407 -3322 26427
rect -3252 26407 -3250 26427
rect -3249 26424 -3235 26427
rect -3228 26427 485 26431
rect -3228 26424 -3211 26427
rect -3228 26407 -3226 26424
rect -3156 26407 -3154 26427
rect -3132 26407 -3130 26427
rect -3060 26407 -3058 26427
rect -3012 26407 -3010 26427
rect -2964 26407 -2962 26427
rect -2916 26407 -2914 26427
rect -2892 26407 -2890 26427
rect -2820 26407 -2818 26427
rect -2796 26407 -2794 26427
rect -2748 26407 -2746 26427
rect -2700 26407 -2698 26427
rect -2604 26407 -2602 26427
rect -2580 26407 -2578 26427
rect -2364 26407 -2362 26427
rect -2292 26407 -2290 26427
rect -2268 26407 -2266 26427
rect -2244 26407 -2242 26427
rect -2172 26407 -2170 26427
rect -2148 26407 -2146 26427
rect -2076 26407 -2074 26427
rect -2052 26407 -2050 26427
rect -1980 26407 -1978 26427
rect -1884 26407 -1882 26427
rect -1836 26407 -1834 26427
rect -1716 26407 -1714 26427
rect -1596 26407 -1594 26427
rect -1476 26407 -1474 26427
rect -1380 26407 -1378 26427
rect -1356 26407 -1354 26427
rect -1308 26407 -1306 26427
rect -1260 26407 -1258 26427
rect -1140 26407 -1138 26427
rect -852 26407 -850 26427
rect -804 26407 -802 26427
rect -756 26407 -754 26427
rect -708 26407 -706 26427
rect -612 26407 -610 26427
rect -588 26407 -586 26427
rect -540 26407 -538 26427
rect -516 26407 -514 26427
rect -492 26407 -490 26427
rect -444 26407 -442 26427
rect -396 26407 -394 26427
rect -300 26407 -298 26427
rect -276 26407 -274 26427
rect -204 26407 -202 26427
rect -108 26407 -106 26427
rect 12 26407 14 26427
rect 108 26407 110 26427
rect 156 26407 158 26427
rect 204 26407 206 26427
rect 228 26407 230 26427
rect 252 26407 254 26427
rect 348 26407 350 26427
rect 468 26407 470 26427
rect 471 26424 485 26427
rect 492 26427 8741 26431
rect 492 26424 509 26427
rect 492 26407 494 26424
rect 564 26407 566 26427
rect 588 26407 590 26427
rect 636 26407 638 26427
rect 660 26407 662 26427
rect 684 26407 686 26427
rect 732 26407 734 26427
rect 756 26407 758 26427
rect 780 26407 782 26427
rect 876 26407 878 26427
rect 972 26407 974 26427
rect 1020 26407 1022 26427
rect 1068 26407 1070 26427
rect 1092 26407 1094 26427
rect 1116 26407 1118 26427
rect 1164 26407 1166 26427
rect 1212 26407 1214 26427
rect 1308 26407 1310 26427
rect 1332 26407 1334 26427
rect 1380 26407 1382 26427
rect 1428 26407 1430 26427
rect 1524 26407 1526 26427
rect 1548 26407 1550 26427
rect 1596 26407 1598 26427
rect 1620 26407 1622 26427
rect 1644 26407 1646 26427
rect 1692 26407 1694 26427
rect 1716 26407 1718 26427
rect 1740 26407 1742 26427
rect 1788 26407 1790 26427
rect 1836 26407 1838 26427
rect 1884 26407 1886 26427
rect 1932 26407 1934 26427
rect 1980 26407 1982 26427
rect 2028 26407 2030 26427
rect 2076 26407 2078 26427
rect 2100 26407 2102 26427
rect 2124 26407 2126 26427
rect 2172 26407 2174 26427
rect 2196 26407 2198 26427
rect 2220 26407 2222 26427
rect 2268 26407 2270 26427
rect 2292 26407 2294 26427
rect 2316 26407 2318 26427
rect 2364 26407 2366 26427
rect 2412 26407 2414 26427
rect 2460 26407 2462 26427
rect 2508 26407 2510 26427
rect 2556 26407 2558 26427
rect 2580 26407 2582 26427
rect 2604 26407 2606 26427
rect 2652 26407 2654 26427
rect 2676 26407 2678 26427
rect 2700 26407 2702 26427
rect 2748 26407 2750 26427
rect 2772 26407 2774 26427
rect 2796 26407 2798 26427
rect 2844 26407 2846 26427
rect 2868 26407 2870 26427
rect 2892 26407 2894 26427
rect 2940 26407 2942 26427
rect 3012 26407 3014 26427
rect 3108 26407 3110 26427
rect 3156 26407 3158 26427
rect 3252 26407 3254 26427
rect 3348 26407 3350 26427
rect 3396 26407 3398 26427
rect 3468 26407 3470 26427
rect 3492 26407 3494 26427
rect 3588 26407 3590 26427
rect 3612 26407 3614 26427
rect 3636 26407 3638 26427
rect 3708 26407 3710 26427
rect 3732 26407 3734 26427
rect 3804 26407 3806 26427
rect 3828 26407 3830 26427
rect 3924 26407 3926 26427
rect 4020 26407 4022 26427
rect 4044 26407 4046 26427
rect 4092 26407 4094 26427
rect 4116 26407 4118 26427
rect 4140 26407 4142 26427
rect 4188 26407 4190 26427
rect 4212 26407 4214 26427
rect 4236 26407 4238 26427
rect 4308 26407 4310 26427
rect 4332 26407 4334 26427
rect 4404 26407 4406 26427
rect 4500 26407 4502 26427
rect 4596 26407 4598 26427
rect 4860 26407 4862 26427
rect 4956 26407 4958 26427
rect 4980 26407 4982 26427
rect 5004 26407 5006 26427
rect 5076 26407 5078 26427
rect 5100 26407 5102 26427
rect 5124 26407 5126 26427
rect 5172 26407 5174 26427
rect 5196 26407 5198 26427
rect 5220 26407 5222 26427
rect 5268 26407 5270 26427
rect 5292 26407 5294 26427
rect 5388 26407 5390 26427
rect 5484 26407 5486 26427
rect 5508 26407 5510 26427
rect 5532 26407 5534 26427
rect 5580 26407 5582 26427
rect 5628 26407 5630 26427
rect 5724 26407 5726 26427
rect 5748 26407 5750 26427
rect 5796 26407 5798 26427
rect 5820 26407 5822 26427
rect 5844 26407 5846 26427
rect 5892 26407 5894 26427
rect 6132 26407 6134 26427
rect 6180 26407 6182 26427
rect 6228 26407 6230 26427
rect 6252 26407 6254 26427
rect 6276 26407 6278 26427
rect 6324 26407 6326 26427
rect 6372 26407 6374 26427
rect 6492 26407 6494 26427
rect 6588 26407 6590 26427
rect 6612 26407 6614 26427
rect 6660 26407 6662 26427
rect 6684 26407 6686 26427
rect 6708 26407 6710 26427
rect 6780 26407 6782 26427
rect 6804 26407 6806 26427
rect 6828 26407 6830 26427
rect 6900 26407 6902 26427
rect 6924 26407 6926 26427
rect 7020 26407 7022 26427
rect 7140 26407 7142 26427
rect 7236 26407 7238 26427
rect 7332 26407 7334 26427
rect 7380 26407 7382 26427
rect 7428 26407 7430 26427
rect 7452 26407 7454 26427
rect 7476 26407 7478 26427
rect 7524 26407 7526 26427
rect 7548 26407 7550 26427
rect 7572 26407 7574 26427
rect 7620 26407 7622 26427
rect 7644 26407 7646 26427
rect 7668 26407 7670 26427
rect 7716 26407 7718 26427
rect 7740 26407 7742 26427
rect 7836 26407 7838 26427
rect 7884 26407 7886 26427
rect 7932 26407 7934 26427
rect 7956 26407 7958 26427
rect 7980 26407 7982 26427
rect 8052 26407 8054 26427
rect 8148 26407 8150 26427
rect 8196 26407 8198 26427
rect 8244 26407 8246 26427
rect 8268 26407 8270 26427
rect 8292 26407 8294 26427
rect 8340 26407 8342 26427
rect 8364 26407 8366 26427
rect 8388 26407 8390 26427
rect 8436 26407 8438 26427
rect 8460 26407 8462 26427
rect 8556 26407 8558 26427
rect 8604 26407 8606 26427
rect 8652 26407 8654 26427
rect 8700 26407 8702 26427
rect 8724 26407 8726 26427
rect 8727 26424 8741 26427
rect 8748 26427 12149 26431
rect 8748 26424 8765 26427
rect 8772 26424 8775 26427
rect 8748 26407 8750 26424
rect 8820 26407 8822 26427
rect 8844 26407 8846 26427
rect 8868 26407 8870 26427
rect 9516 26407 9518 26427
rect 9612 26407 9614 26427
rect 9660 26407 9662 26427
rect 9684 26407 9686 26427
rect 9708 26407 9710 26427
rect 9756 26407 9758 26427
rect 9780 26407 9782 26427
rect 9804 26407 9806 26427
rect 9852 26407 9854 26427
rect 9876 26407 9878 26427
rect 9900 26407 9902 26427
rect 9948 26407 9950 26427
rect 9972 26407 9974 26427
rect 9996 26407 9998 26427
rect 10068 26407 10070 26427
rect 10092 26407 10094 26427
rect 10116 26407 10118 26427
rect 10164 26407 10166 26427
rect 10188 26407 10190 26427
rect 10212 26407 10214 26427
rect 10260 26407 10262 26427
rect 10284 26407 10286 26427
rect 10308 26407 10310 26427
rect 10380 26407 10382 26427
rect 10404 26407 10406 26427
rect 10428 26407 10430 26427
rect 10476 26407 10478 26427
rect 10500 26407 10502 26427
rect 10524 26407 10526 26427
rect 10572 26407 10574 26427
rect 10596 26407 10598 26427
rect 10620 26407 10622 26427
rect 10668 26407 10670 26427
rect 10692 26407 10694 26427
rect 10716 26407 10718 26427
rect 10788 26407 10790 26427
rect 10836 26407 10838 26427
rect 10956 26407 10958 26427
rect 11052 26407 11054 26427
rect 11076 26407 11078 26427
rect 11124 26407 11126 26427
rect 11172 26407 11174 26427
rect 11220 26407 11222 26427
rect 11340 26407 11342 26427
rect 11436 26407 11438 26427
rect 11532 26407 11534 26427
rect 11580 26407 11582 26427
rect 11628 26407 11630 26427
rect 11676 26407 11678 26427
rect 11772 26407 11774 26427
rect 11796 26407 11798 26427
rect 11844 26407 11846 26427
rect 11892 26407 11894 26427
rect 11988 26407 11990 26427
rect 12060 26407 12062 26427
rect 12132 26407 12134 26427
rect 12135 26424 12149 26427
rect 12159 26427 31253 26431
rect 12159 26424 12173 26427
rect 12228 26407 12230 26427
rect 12324 26407 12326 26427
rect 12420 26407 12422 26427
rect 12444 26407 12446 26427
rect 12492 26407 12494 26427
rect 12516 26407 12518 26427
rect 12540 26407 12542 26427
rect 12588 26407 12590 26427
rect 12636 26407 12638 26427
rect 12732 26407 12734 26427
rect 12756 26407 12758 26427
rect 12804 26407 12806 26427
rect 12828 26407 12830 26427
rect 12852 26407 12854 26427
rect 12900 26407 12902 26427
rect 12948 26407 12950 26427
rect 13044 26407 13046 26427
rect 13068 26407 13070 26427
rect 13116 26407 13118 26427
rect 13284 26407 13286 26427
rect 13332 26407 13334 26427
rect 13428 26407 13430 26427
rect 13524 26407 13526 26427
rect 13572 26407 13574 26427
rect 13644 26407 13646 26427
rect 13668 26407 13670 26427
rect 13764 26407 13766 26427
rect 13812 26407 13814 26427
rect 13860 26407 13862 26427
rect 13908 26407 13910 26427
rect 13956 26407 13958 26427
rect 14004 26407 14006 26427
rect 14100 26407 14102 26427
rect 14196 26407 14198 26427
rect 14244 26407 14246 26427
rect 14292 26407 14294 26427
rect 15132 26407 15134 26427
rect 15228 26407 15230 26427
rect 15252 26407 15254 26427
rect 15300 26407 15302 26427
rect 15324 26407 15326 26427
rect 15396 26407 15398 26427
rect 15420 26407 15422 26427
rect 15492 26407 15494 26427
rect 15540 26407 15542 26427
rect 15636 26407 15638 26427
rect 15660 26407 15662 26427
rect 15708 26407 15710 26427
rect 15732 26407 15734 26427
rect 15756 26407 15758 26427
rect 15804 26407 15806 26427
rect 15828 26407 15830 26427
rect 15852 26407 15854 26427
rect 15900 26407 15902 26427
rect 15948 26407 15950 26427
rect 15996 26407 15998 26427
rect 16044 26407 16046 26427
rect 16092 26407 16094 26427
rect 16140 26407 16142 26427
rect 16236 26407 16238 26427
rect 16260 26407 16262 26427
rect 16308 26407 16310 26427
rect 16332 26407 16334 26427
rect 16356 26407 16358 26427
rect 16404 26407 16406 26427
rect 16452 26407 16454 26427
rect 16548 26407 16550 26427
rect 16572 26407 16574 26427
rect 16620 26407 16622 26427
rect 16668 26407 16670 26427
rect 16716 26407 16718 26427
rect 16764 26407 16766 26427
rect 16836 26407 16838 26427
rect 16884 26407 16886 26427
rect 16980 26407 16982 26427
rect 17052 26407 17054 26427
rect 17196 26407 17198 26427
rect 17220 26407 17222 26427
rect 17292 26407 17294 26427
rect 17316 26407 17318 26427
rect 18084 26407 18086 26427
rect 18132 26407 18134 26427
rect 18396 26407 18398 26427
rect 18492 26407 18494 26427
rect 18516 26407 18518 26427
rect 18564 26407 18566 26427
rect 18612 26407 18614 26427
rect 18660 26407 18662 26427
rect 18708 26407 18710 26427
rect 18756 26407 18758 26427
rect 18804 26407 18806 26427
rect 18852 26407 18854 26427
rect 18900 26407 18902 26427
rect 18996 26407 18998 26427
rect 19020 26407 19022 26427
rect 19092 26407 19094 26427
rect 19116 26407 19118 26427
rect 19140 26407 19142 26427
rect 19188 26407 19190 26427
rect 19236 26407 19238 26427
rect 19332 26407 19334 26427
rect 19476 26407 19478 26427
rect 19620 26407 19622 26427
rect 19716 26407 19718 26427
rect 19788 26407 19790 26427
rect 19836 26407 19838 26427
rect 19860 26407 19862 26427
rect 19884 26407 19886 26427
rect 19932 26407 19934 26427
rect 19956 26407 19958 26427
rect 19980 26407 19982 26427
rect 20028 26407 20030 26427
rect 20052 26407 20054 26427
rect 20076 26407 20078 26427
rect 20148 26407 20150 26427
rect 20172 26407 20174 26427
rect 20196 26407 20198 26427
rect 20268 26407 20270 26427
rect 20292 26407 20294 26427
rect 20388 26407 20390 26427
rect 20412 26407 20414 26427
rect 20508 26407 20510 26427
rect 20556 26407 20558 26427
rect 20604 26407 20606 26427
rect 20916 26407 20918 26427
rect 20964 26407 20966 26427
rect 21012 26407 21014 26427
rect 21060 26407 21062 26427
rect 21084 26407 21086 26427
rect 21108 26407 21110 26427
rect 21204 26407 21206 26427
rect 21300 26407 21302 26427
rect 21324 26407 21326 26427
rect 21444 26407 21446 26427
rect 21468 26407 21470 26427
rect 21564 26407 21566 26427
rect 21612 26407 21614 26427
rect 21684 26407 21686 26427
rect 21708 26407 21710 26427
rect 21804 26407 21806 26427
rect 21828 26407 21830 26427
rect 21924 26407 21926 26427
rect 21948 26407 21950 26427
rect 22044 26407 22046 26427
rect 22068 26407 22070 26427
rect 22188 26407 22190 26427
rect 22212 26407 22214 26427
rect 23004 26407 23006 26427
rect 23052 26407 23054 26427
rect 23076 26407 23078 26427
rect 23100 26407 23102 26427
rect 23148 26407 23150 26427
rect 23220 26407 23222 26427
rect 23244 26407 23246 26427
rect 23316 26407 23318 26427
rect 23340 26407 23342 26427
rect 23412 26407 23414 26427
rect 23556 26407 23558 26427
rect 23628 26407 23630 26427
rect 23652 26407 23654 26427
rect 23676 26407 23678 26427
rect 23724 26407 23726 26427
rect 23772 26407 23774 26427
rect 23820 26407 23822 26427
rect 23868 26407 23870 26427
rect 23916 26407 23918 26427
rect 24012 26407 24014 26427
rect 24084 26407 24086 26427
rect 24372 26407 24374 26427
rect 24396 26407 24398 26427
rect 24492 26407 24494 26427
rect 24516 26407 24518 26427
rect 24588 26407 24590 26427
rect 24612 26407 24614 26427
rect 24708 26407 24710 26427
rect 24732 26407 24734 26427
rect 24756 26407 24758 26427
rect 24852 26407 24854 26427
rect 24876 26407 24878 26427
rect 24972 26407 24974 26427
rect 24996 26407 24998 26427
rect 25092 26407 25094 26427
rect 25260 26407 25262 26427
rect 25356 26407 25358 26427
rect 25380 26407 25382 26427
rect 25452 26407 25454 26427
rect 25476 26407 25478 26427
rect 25500 26407 25502 26427
rect 25572 26407 25574 26427
rect 25596 26407 25598 26427
rect 27060 26407 27062 26427
rect 27108 26407 27110 26427
rect 27180 26407 27182 26427
rect 27324 26407 27326 26427
rect 27396 26407 27398 26427
rect 27420 26407 27422 26427
rect 27540 26407 27542 26427
rect 27564 26407 27566 26427
rect 30564 26407 30567 26424
rect 30636 26407 30638 26427
rect 30660 26407 30662 26427
rect 30780 26407 30782 26427
rect 30804 26407 30806 26427
rect 30924 26407 30926 26427
rect 30948 26407 30950 26427
rect 31068 26407 31070 26427
rect 31092 26407 31094 26427
rect 31164 26407 31166 26427
rect 31236 26407 31238 26427
rect 31239 26424 31253 26427
rect 31263 26427 31835 26431
rect 31897 26431 31931 26432
rect 31969 26431 32003 26432
rect 31897 26427 32003 26431
rect 31263 26424 31277 26427
rect 31897 26422 31900 26427
rect 31908 26424 31910 26427
rect 31908 26422 31911 26424
rect 31907 26408 31911 26422
rect 31993 26414 31997 26422
rect 31983 26408 31993 26414
rect 31441 26407 31475 26408
rect -16295 26403 -14683 26407
rect -16295 26398 -16292 26403
rect -16284 26398 -16282 26403
rect -16285 26384 -16282 26398
rect -16271 26390 -16267 26398
rect -16281 26384 -16271 26390
rect -16271 26383 -16267 26384
rect -16703 26379 -16267 26383
rect -16668 26359 -16666 26379
rect -16596 26376 -16594 26379
rect -16596 26359 -16593 26376
rect -16500 26359 -16498 26379
rect -16415 26374 -16412 26379
rect -16404 26374 -16402 26379
rect -16405 26360 -16402 26374
rect -16380 26359 -16378 26379
rect -16356 26359 -16354 26379
rect -16308 26376 -16306 26379
rect -16281 26376 -16267 26379
rect -16308 26359 -16305 26376
rect -16271 26374 -16268 26376
rect -16261 26360 -16258 26374
rect -16260 26359 -16258 26360
rect -16236 26359 -16234 26403
rect -16212 26359 -16210 26403
rect -16188 26400 -16186 26403
rect -16188 26384 -16185 26400
rect -15383 26398 -15380 26403
rect -15372 26398 -15370 26403
rect -15373 26384 -15370 26398
rect -16199 26383 -16165 26384
rect -15300 26383 -15298 26403
rect -15084 26383 -15082 26403
rect -15036 26383 -15034 26403
rect -14868 26383 -14866 26403
rect -14772 26383 -14770 26403
rect -14724 26383 -14722 26403
rect -14697 26400 -14683 26403
rect -14673 26403 -12979 26407
rect -14673 26400 -14659 26403
rect -14652 26400 -14649 26403
rect -14508 26383 -14506 26403
rect -14436 26383 -14434 26403
rect -14388 26383 -14386 26403
rect -14268 26400 -14266 26403
rect -14268 26383 -14265 26400
rect -14172 26383 -14170 26403
rect -14076 26383 -14074 26403
rect -14028 26383 -14026 26403
rect -13980 26383 -13978 26403
rect -13956 26400 -13954 26403
rect -13956 26384 -13953 26400
rect -13967 26383 -13933 26384
rect -13932 26383 -13930 26403
rect -13860 26383 -13858 26403
rect -13764 26383 -13762 26403
rect -13716 26383 -13714 26403
rect -13644 26383 -13642 26403
rect -13596 26383 -13594 26403
rect -13500 26383 -13498 26403
rect -13404 26383 -13402 26403
rect -13356 26383 -13354 26403
rect -13284 26383 -13282 26403
rect -13068 26383 -13066 26403
rect -12993 26400 -12979 26403
rect -12969 26403 -8251 26407
rect -12969 26400 -12955 26403
rect -12828 26383 -12826 26403
rect -12780 26383 -12778 26403
rect -12660 26383 -12658 26403
rect -12564 26383 -12562 26403
rect -12492 26383 -12490 26403
rect -12396 26383 -12394 26403
rect -12348 26383 -12346 26403
rect -12276 26383 -12274 26403
rect -12252 26383 -12250 26403
rect -12156 26383 -12154 26403
rect -12060 26383 -12058 26403
rect -12012 26384 -12010 26403
rect -12023 26383 -11989 26384
rect -11916 26383 -11914 26403
rect -11892 26383 -11890 26403
rect -11844 26383 -11842 26403
rect -11796 26383 -11794 26403
rect -11676 26383 -11674 26403
rect -11580 26383 -11578 26403
rect -11556 26383 -11554 26403
rect -11484 26383 -11482 26403
rect -11460 26383 -11458 26403
rect -11436 26383 -11434 26403
rect -11388 26383 -11386 26403
rect -11364 26383 -11362 26403
rect -11340 26383 -11338 26403
rect -11268 26383 -11266 26403
rect -11172 26383 -11170 26403
rect -11124 26383 -11122 26403
rect -11076 26383 -11074 26403
rect -11028 26383 -11026 26403
rect -10788 26383 -10786 26403
rect -10668 26383 -10666 26403
rect -9876 26383 -9874 26403
rect -9828 26383 -9826 26403
rect -9732 26383 -9730 26403
rect -9708 26383 -9706 26403
rect -9612 26383 -9610 26403
rect -9516 26383 -9514 26403
rect -9468 26383 -9466 26403
rect -9420 26383 -9418 26403
rect -9396 26383 -9394 26403
rect -9372 26383 -9370 26403
rect -9300 26383 -9298 26403
rect -9252 26383 -9250 26403
rect -9132 26383 -9130 26403
rect -9084 26383 -9082 26403
rect -9036 26383 -9034 26403
rect -8988 26383 -8986 26403
rect -8940 26383 -8938 26403
rect -8892 26383 -8890 26403
rect -8844 26383 -8842 26403
rect -8796 26384 -8794 26403
rect -8807 26383 -8773 26384
rect -8700 26383 -8698 26403
rect -8604 26383 -8602 26403
rect -8508 26383 -8506 26403
rect -8484 26383 -8482 26403
rect -8388 26383 -8386 26403
rect -8364 26383 -8362 26403
rect -8340 26383 -8338 26403
rect -8292 26383 -8290 26403
rect -8268 26383 -8266 26403
rect -8265 26400 -8251 26403
rect -8241 26403 30557 26407
rect -8241 26400 -8227 26403
rect -8196 26383 -8194 26403
rect -8100 26383 -8098 26403
rect -8052 26383 -8050 26403
rect -7932 26383 -7930 26403
rect -7836 26383 -7834 26403
rect -7740 26383 -7738 26403
rect -7692 26383 -7690 26403
rect -7620 26383 -7618 26403
rect -7404 26383 -7402 26403
rect -7356 26383 -7354 26403
rect -7308 26383 -7306 26403
rect -7212 26383 -7210 26403
rect -7188 26383 -7186 26403
rect -7116 26383 -7114 26403
rect -7068 26383 -7066 26403
rect -6972 26383 -6970 26403
rect -6948 26383 -6946 26403
rect -6876 26383 -6874 26403
rect -6852 26383 -6850 26403
rect -6804 26383 -6802 26403
rect -6780 26383 -6778 26403
rect -6756 26383 -6754 26403
rect -6708 26383 -6706 26403
rect -6684 26383 -6682 26403
rect -6660 26383 -6658 26403
rect -6612 26383 -6610 26403
rect -6588 26383 -6586 26403
rect -6564 26383 -6562 26403
rect -6516 26383 -6514 26403
rect -6492 26383 -6490 26403
rect -6468 26383 -6466 26403
rect -6420 26383 -6418 26403
rect -6396 26383 -6394 26403
rect -6372 26383 -6370 26403
rect -6324 26383 -6322 26403
rect -6300 26383 -6298 26403
rect -6276 26383 -6274 26403
rect -6228 26383 -6226 26403
rect -6180 26383 -6178 26403
rect -6060 26383 -6058 26403
rect -5964 26383 -5962 26403
rect -5940 26383 -5938 26403
rect -5868 26383 -5866 26403
rect -5652 26383 -5650 26403
rect -5316 26383 -5314 26403
rect -5268 26383 -5266 26403
rect -5196 26383 -5194 26403
rect -5172 26383 -5170 26403
rect -5100 26383 -5098 26403
rect -5076 26383 -5074 26403
rect -4980 26383 -4978 26403
rect -4956 26383 -4954 26403
rect -4884 26383 -4882 26403
rect -4860 26383 -4858 26403
rect -4788 26383 -4786 26403
rect -4692 26383 -4690 26403
rect -4644 26383 -4642 26403
rect -4596 26383 -4594 26403
rect -4548 26383 -4546 26403
rect -4428 26383 -4426 26403
rect -4332 26383 -4330 26403
rect -4308 26383 -4306 26403
rect -4260 26383 -4258 26403
rect -4212 26383 -4210 26403
rect -4116 26383 -4114 26403
rect -4092 26383 -4090 26403
rect -4020 26383 -4018 26403
rect -3876 26383 -3874 26403
rect -3732 26383 -3730 26403
rect -3588 26383 -3586 26403
rect -3564 26383 -3562 26403
rect -3516 26383 -3514 26403
rect -3492 26383 -3490 26403
rect -3468 26383 -3466 26403
rect -3420 26383 -3418 26403
rect -3324 26383 -3322 26403
rect -3252 26383 -3250 26403
rect -3228 26383 -3226 26403
rect -3156 26383 -3154 26403
rect -3132 26383 -3130 26403
rect -3060 26383 -3058 26403
rect -3012 26383 -3010 26403
rect -2964 26383 -2962 26403
rect -2916 26383 -2914 26403
rect -2892 26383 -2890 26403
rect -2820 26383 -2818 26403
rect -2796 26383 -2794 26403
rect -2748 26383 -2746 26403
rect -2700 26383 -2698 26403
rect -2604 26383 -2602 26403
rect -2580 26383 -2578 26403
rect -2364 26383 -2362 26403
rect -2292 26383 -2290 26403
rect -2268 26383 -2266 26403
rect -2244 26383 -2242 26403
rect -2172 26383 -2170 26403
rect -2148 26383 -2146 26403
rect -2076 26383 -2074 26403
rect -2052 26383 -2050 26403
rect -1980 26383 -1978 26403
rect -1884 26383 -1882 26403
rect -1836 26383 -1834 26403
rect -1716 26383 -1714 26403
rect -1596 26383 -1594 26403
rect -1476 26383 -1474 26403
rect -1380 26383 -1378 26403
rect -1356 26383 -1354 26403
rect -1308 26383 -1306 26403
rect -1260 26383 -1258 26403
rect -1140 26383 -1138 26403
rect -852 26383 -850 26403
rect -804 26383 -802 26403
rect -756 26383 -754 26403
rect -708 26383 -706 26403
rect -612 26383 -610 26403
rect -588 26383 -586 26403
rect -540 26383 -538 26403
rect -516 26383 -514 26403
rect -492 26383 -490 26403
rect -444 26383 -442 26403
rect -396 26383 -394 26403
rect -300 26383 -298 26403
rect -276 26383 -274 26403
rect -204 26383 -202 26403
rect -108 26383 -106 26403
rect 12 26383 14 26403
rect 108 26383 110 26403
rect 156 26383 158 26403
rect 204 26383 206 26403
rect 228 26383 230 26403
rect 252 26383 254 26403
rect 348 26383 350 26403
rect 468 26383 470 26403
rect 492 26383 494 26403
rect 564 26383 566 26403
rect 588 26383 590 26403
rect 636 26383 638 26403
rect 660 26383 662 26403
rect 684 26383 686 26403
rect 732 26383 734 26403
rect 756 26383 758 26403
rect 780 26383 782 26403
rect 876 26383 878 26403
rect 972 26383 974 26403
rect 1020 26383 1022 26403
rect 1068 26383 1070 26403
rect 1092 26383 1094 26403
rect 1116 26383 1118 26403
rect 1164 26383 1166 26403
rect 1212 26383 1214 26403
rect 1308 26383 1310 26403
rect 1332 26383 1334 26403
rect 1380 26383 1382 26403
rect 1428 26383 1430 26403
rect 1524 26383 1526 26403
rect 1548 26383 1550 26403
rect 1596 26383 1598 26403
rect 1620 26383 1622 26403
rect 1644 26383 1646 26403
rect 1692 26383 1694 26403
rect 1716 26383 1718 26403
rect 1740 26383 1742 26403
rect 1788 26383 1790 26403
rect 1836 26383 1838 26403
rect 1884 26383 1886 26403
rect 1932 26383 1934 26403
rect 1980 26383 1982 26403
rect 2028 26383 2030 26403
rect 2076 26383 2078 26403
rect 2100 26383 2102 26403
rect 2124 26383 2126 26403
rect 2172 26383 2174 26403
rect 2196 26383 2198 26403
rect 2220 26383 2222 26403
rect 2268 26383 2270 26403
rect 2292 26383 2294 26403
rect 2316 26383 2318 26403
rect 2364 26383 2366 26403
rect 2412 26383 2414 26403
rect 2460 26383 2462 26403
rect 2508 26383 2510 26403
rect 2556 26383 2558 26403
rect 2580 26383 2582 26403
rect 2604 26383 2606 26403
rect 2652 26383 2654 26403
rect 2676 26383 2678 26403
rect 2700 26383 2702 26403
rect 2748 26383 2750 26403
rect 2772 26383 2774 26403
rect 2796 26383 2798 26403
rect 2844 26383 2846 26403
rect 2868 26383 2870 26403
rect 2892 26383 2894 26403
rect 2940 26383 2942 26403
rect 3012 26383 3014 26403
rect 3108 26383 3110 26403
rect 3156 26383 3158 26403
rect 3252 26383 3254 26403
rect 3348 26383 3350 26403
rect 3396 26383 3398 26403
rect 3468 26383 3470 26403
rect 3492 26383 3494 26403
rect 3588 26383 3590 26403
rect 3612 26383 3614 26403
rect 3636 26383 3638 26403
rect 3708 26383 3710 26403
rect 3732 26383 3734 26403
rect 3804 26383 3806 26403
rect 3828 26383 3830 26403
rect 3924 26383 3926 26403
rect 4020 26383 4022 26403
rect 4044 26383 4046 26403
rect 4092 26383 4094 26403
rect 4116 26383 4118 26403
rect 4140 26383 4142 26403
rect 4188 26383 4190 26403
rect 4212 26383 4214 26403
rect 4236 26383 4238 26403
rect 4308 26383 4310 26403
rect 4332 26383 4334 26403
rect 4404 26383 4406 26403
rect 4500 26383 4502 26403
rect 4596 26383 4598 26403
rect 4860 26383 4862 26403
rect 4956 26383 4958 26403
rect 4980 26383 4982 26403
rect 5004 26383 5006 26403
rect 5076 26383 5078 26403
rect 5100 26383 5102 26403
rect 5124 26383 5126 26403
rect 5172 26383 5174 26403
rect 5196 26383 5198 26403
rect 5220 26383 5222 26403
rect 5268 26383 5270 26403
rect 5292 26383 5294 26403
rect 5388 26383 5390 26403
rect 5484 26383 5486 26403
rect 5508 26383 5510 26403
rect 5532 26383 5534 26403
rect 5580 26383 5582 26403
rect 5628 26383 5630 26403
rect 5724 26384 5726 26403
rect 5713 26383 5747 26384
rect 5748 26383 5750 26403
rect 5796 26383 5798 26403
rect 5820 26383 5822 26403
rect 5844 26383 5846 26403
rect 5892 26383 5894 26403
rect 6132 26383 6134 26403
rect 6180 26383 6182 26403
rect 6228 26383 6230 26403
rect 6252 26383 6254 26403
rect 6276 26383 6278 26403
rect 6324 26383 6326 26403
rect 6372 26383 6374 26403
rect 6492 26383 6494 26403
rect 6588 26383 6590 26403
rect 6612 26383 6614 26403
rect 6660 26383 6662 26403
rect 6684 26383 6686 26403
rect 6708 26383 6710 26403
rect 6780 26383 6782 26403
rect 6804 26383 6806 26403
rect 6828 26383 6830 26403
rect 6900 26383 6902 26403
rect 6924 26383 6926 26403
rect 7020 26383 7022 26403
rect 7140 26383 7142 26403
rect 7236 26383 7238 26403
rect 7332 26383 7334 26403
rect 7380 26383 7382 26403
rect 7428 26383 7430 26403
rect 7452 26383 7454 26403
rect 7476 26383 7478 26403
rect 7524 26383 7526 26403
rect 7548 26383 7550 26403
rect 7572 26383 7574 26403
rect 7620 26383 7622 26403
rect 7644 26383 7646 26403
rect 7668 26383 7670 26403
rect 7716 26383 7718 26403
rect 7740 26383 7742 26403
rect 7836 26383 7838 26403
rect 7884 26383 7886 26403
rect 7932 26383 7934 26403
rect 7956 26383 7958 26403
rect 7980 26383 7982 26403
rect 8052 26383 8054 26403
rect 8148 26383 8150 26403
rect 8196 26383 8198 26403
rect 8244 26383 8246 26403
rect 8268 26383 8270 26403
rect 8292 26383 8294 26403
rect 8340 26383 8342 26403
rect 8364 26383 8366 26403
rect 8388 26383 8390 26403
rect 8436 26383 8438 26403
rect 8460 26383 8462 26403
rect 8556 26383 8558 26403
rect 8604 26383 8606 26403
rect 8652 26383 8654 26403
rect 8700 26383 8702 26403
rect 8724 26383 8726 26403
rect 8748 26383 8750 26403
rect 8820 26383 8822 26403
rect 8844 26383 8846 26403
rect 8868 26383 8870 26403
rect 9516 26383 9518 26403
rect 9612 26383 9614 26403
rect 9660 26383 9662 26403
rect 9684 26383 9686 26403
rect 9708 26383 9710 26403
rect 9756 26383 9758 26403
rect 9780 26383 9782 26403
rect 9804 26383 9806 26403
rect 9852 26383 9854 26403
rect 9876 26383 9878 26403
rect 9900 26383 9902 26403
rect 9948 26383 9950 26403
rect 9972 26383 9974 26403
rect 9996 26383 9998 26403
rect 10068 26383 10070 26403
rect 10092 26383 10094 26403
rect 10116 26383 10118 26403
rect 10164 26383 10166 26403
rect 10188 26383 10190 26403
rect 10212 26383 10214 26403
rect 10260 26383 10262 26403
rect 10284 26383 10286 26403
rect 10308 26383 10310 26403
rect 10380 26383 10382 26403
rect 10404 26383 10406 26403
rect 10428 26383 10430 26403
rect 10476 26383 10478 26403
rect 10500 26383 10502 26403
rect 10524 26383 10526 26403
rect 10572 26383 10574 26403
rect 10596 26383 10598 26403
rect 10620 26383 10622 26403
rect 10668 26383 10670 26403
rect 10692 26383 10694 26403
rect 10716 26383 10718 26403
rect 10788 26383 10790 26403
rect 10836 26383 10838 26403
rect 10956 26383 10958 26403
rect 11052 26383 11054 26403
rect 11076 26383 11078 26403
rect 11124 26383 11126 26403
rect 11172 26383 11174 26403
rect 11220 26383 11222 26403
rect 11340 26383 11342 26403
rect 11436 26383 11438 26403
rect 11532 26383 11534 26403
rect 11580 26383 11582 26403
rect 11628 26383 11630 26403
rect 11676 26383 11678 26403
rect 11772 26383 11774 26403
rect 11796 26383 11798 26403
rect 11844 26383 11846 26403
rect 11892 26383 11894 26403
rect 11988 26383 11990 26403
rect 12060 26383 12062 26403
rect 12132 26383 12134 26403
rect 12228 26383 12230 26403
rect 12324 26383 12326 26403
rect 12420 26383 12422 26403
rect 12444 26383 12446 26403
rect 12492 26383 12494 26403
rect 12516 26383 12518 26403
rect 12540 26383 12542 26403
rect 12588 26383 12590 26403
rect 12636 26383 12638 26403
rect 12732 26383 12734 26403
rect 12756 26383 12758 26403
rect 12804 26383 12806 26403
rect 12828 26383 12830 26403
rect 12852 26383 12854 26403
rect 12900 26383 12902 26403
rect 12948 26383 12950 26403
rect 13044 26383 13046 26403
rect 13068 26383 13070 26403
rect 13116 26383 13118 26403
rect 13284 26383 13286 26403
rect 13332 26383 13334 26403
rect 13428 26383 13430 26403
rect 13524 26383 13526 26403
rect 13572 26383 13574 26403
rect 13644 26383 13646 26403
rect 13668 26383 13670 26403
rect 13764 26383 13766 26403
rect 13812 26383 13814 26403
rect 13860 26383 13862 26403
rect 13908 26383 13910 26403
rect 13956 26383 13958 26403
rect 14004 26383 14006 26403
rect 14100 26383 14102 26403
rect 14196 26383 14198 26403
rect 14244 26383 14246 26403
rect 14292 26383 14294 26403
rect 15132 26383 15134 26403
rect 15228 26383 15230 26403
rect 15252 26383 15254 26403
rect 15300 26383 15302 26403
rect 15324 26383 15326 26403
rect 15396 26383 15398 26403
rect 15420 26383 15422 26403
rect 15492 26383 15494 26403
rect 15540 26383 15542 26403
rect 15636 26383 15638 26403
rect 15660 26383 15662 26403
rect 15708 26383 15710 26403
rect 15732 26383 15734 26403
rect 15756 26383 15758 26403
rect 15804 26383 15806 26403
rect 15828 26383 15830 26403
rect 15852 26383 15854 26403
rect 15900 26383 15902 26403
rect 15948 26383 15950 26403
rect 15996 26383 15998 26403
rect 16044 26383 16046 26403
rect 16092 26383 16094 26403
rect 16140 26383 16142 26403
rect 16236 26383 16238 26403
rect 16260 26383 16262 26403
rect 16308 26383 16310 26403
rect 16332 26383 16334 26403
rect 16356 26383 16358 26403
rect 16404 26383 16406 26403
rect 16452 26383 16454 26403
rect 16548 26383 16550 26403
rect 16572 26383 16574 26403
rect 16620 26383 16622 26403
rect 16668 26383 16670 26403
rect 16716 26383 16718 26403
rect 16764 26383 16766 26403
rect 16836 26383 16838 26403
rect 16884 26383 16886 26403
rect 16980 26383 16982 26403
rect 17052 26383 17054 26403
rect 17196 26383 17198 26403
rect 17220 26383 17222 26403
rect 17292 26383 17294 26403
rect 17316 26383 17318 26403
rect 18084 26383 18086 26403
rect 18132 26383 18134 26403
rect 18396 26383 18398 26403
rect 18492 26383 18494 26403
rect 18516 26383 18518 26403
rect 18564 26383 18566 26403
rect 18612 26383 18614 26403
rect 18660 26383 18662 26403
rect 18708 26383 18710 26403
rect 18756 26383 18758 26403
rect 18804 26383 18806 26403
rect 18852 26383 18854 26403
rect 18900 26383 18902 26403
rect 18996 26383 18998 26403
rect 19020 26383 19022 26403
rect 19092 26383 19094 26403
rect 19116 26383 19118 26403
rect 19140 26383 19142 26403
rect 19188 26383 19190 26403
rect 19236 26383 19238 26403
rect 19332 26383 19334 26403
rect 19476 26383 19478 26403
rect 19620 26383 19622 26403
rect 19716 26383 19718 26403
rect 19788 26383 19790 26403
rect 19836 26383 19838 26403
rect 19860 26383 19862 26403
rect 19884 26383 19886 26403
rect 19932 26383 19934 26403
rect 19956 26383 19958 26403
rect 19980 26383 19982 26403
rect 20028 26383 20030 26403
rect 20052 26383 20054 26403
rect 20076 26383 20078 26403
rect 20148 26383 20150 26403
rect 20172 26383 20174 26403
rect 20196 26383 20198 26403
rect 20268 26383 20270 26403
rect 20292 26383 20294 26403
rect 20388 26383 20390 26403
rect 20412 26383 20414 26403
rect 20508 26383 20510 26403
rect 20556 26383 20558 26403
rect 20604 26383 20606 26403
rect 20916 26383 20918 26403
rect 20964 26383 20966 26403
rect 21012 26383 21014 26403
rect 21060 26383 21062 26403
rect 21084 26383 21086 26403
rect 21108 26383 21110 26403
rect 21204 26383 21206 26403
rect 21300 26383 21302 26403
rect 21324 26383 21326 26403
rect 21444 26383 21446 26403
rect 21468 26383 21470 26403
rect 21564 26383 21566 26403
rect 21612 26383 21614 26403
rect 21684 26383 21686 26403
rect 21708 26383 21710 26403
rect 21804 26383 21806 26403
rect 21828 26383 21830 26403
rect 21924 26383 21926 26403
rect 21948 26383 21950 26403
rect 22044 26383 22046 26403
rect 22068 26383 22070 26403
rect 22188 26383 22190 26403
rect 22212 26383 22214 26403
rect 23004 26383 23006 26403
rect 23052 26383 23054 26403
rect 23076 26383 23078 26403
rect 23100 26383 23102 26403
rect 23148 26383 23150 26403
rect 23220 26383 23222 26403
rect 23244 26383 23246 26403
rect 23316 26383 23318 26403
rect 23340 26383 23342 26403
rect 23412 26383 23414 26403
rect 23556 26383 23558 26403
rect 23628 26383 23630 26403
rect 23652 26383 23654 26403
rect 23676 26383 23678 26403
rect 23724 26383 23726 26403
rect 23772 26383 23774 26403
rect 23820 26383 23822 26403
rect 23868 26383 23870 26403
rect 23916 26383 23918 26403
rect 24012 26383 24014 26403
rect 24084 26383 24086 26403
rect 24372 26383 24374 26403
rect 24396 26383 24398 26403
rect 24492 26383 24494 26403
rect 24516 26383 24518 26403
rect 24588 26383 24590 26403
rect 24612 26383 24614 26403
rect 24708 26383 24710 26403
rect 24732 26383 24734 26403
rect 24756 26383 24758 26403
rect 24852 26383 24854 26403
rect 24876 26383 24878 26403
rect 24972 26383 24974 26403
rect 24996 26383 24998 26403
rect 25092 26383 25094 26403
rect 25260 26383 25262 26403
rect 25356 26383 25358 26403
rect 25380 26383 25382 26403
rect 25452 26383 25454 26403
rect 25476 26384 25478 26403
rect 25465 26383 25499 26384
rect 25500 26383 25502 26403
rect 25572 26383 25574 26403
rect 25596 26383 25598 26403
rect 27060 26383 27062 26403
rect 27108 26383 27110 26403
rect 27180 26383 27182 26403
rect 27324 26383 27326 26403
rect 27396 26383 27398 26403
rect 27420 26383 27422 26403
rect 27540 26383 27542 26403
rect 27564 26383 27566 26403
rect 30543 26400 30557 26403
rect 30564 26403 31475 26407
rect 30564 26400 30581 26403
rect 30564 26383 30566 26400
rect 30636 26383 30638 26403
rect 30660 26383 30662 26403
rect 30780 26383 30782 26403
rect 30804 26383 30806 26403
rect 30924 26383 30926 26403
rect 30948 26383 30950 26403
rect 31068 26383 31070 26403
rect 31092 26383 31094 26403
rect 31164 26383 31166 26403
rect 31236 26383 31238 26403
rect 31393 26383 31427 26384
rect -16199 26379 31427 26383
rect -16199 26376 -16195 26379
rect -16188 26376 -16185 26379
rect -16175 26366 -16171 26374
rect -16185 26360 -16175 26366
rect -15300 26359 -15298 26379
rect -15297 26376 -15283 26379
rect -15084 26359 -15082 26379
rect -15036 26359 -15034 26379
rect -14868 26359 -14866 26379
rect -14772 26359 -14770 26379
rect -14724 26359 -14722 26379
rect -14508 26359 -14506 26379
rect -14436 26359 -14434 26379
rect -14388 26359 -14386 26379
rect -14289 26376 -14275 26379
rect -14268 26376 -14265 26379
rect -14172 26359 -14170 26379
rect -14135 26359 -14101 26360
rect -14076 26359 -14074 26379
rect -14028 26359 -14026 26379
rect -13980 26359 -13978 26379
rect -13977 26376 -13963 26379
rect -13956 26376 -13953 26379
rect -13932 26359 -13930 26379
rect -13860 26376 -13858 26379
rect -13860 26359 -13857 26376
rect -13764 26359 -13762 26379
rect -13716 26359 -13714 26379
rect -13644 26359 -13642 26379
rect -13596 26359 -13594 26379
rect -13500 26359 -13498 26379
rect -13404 26359 -13402 26379
rect -13356 26359 -13354 26379
rect -13284 26359 -13282 26379
rect -13068 26359 -13066 26379
rect -12828 26359 -12826 26379
rect -12780 26359 -12778 26379
rect -12660 26359 -12658 26379
rect -12564 26359 -12562 26379
rect -12492 26359 -12490 26379
rect -12396 26359 -12394 26379
rect -12348 26359 -12346 26379
rect -12276 26359 -12274 26379
rect -12252 26359 -12250 26379
rect -12156 26359 -12154 26379
rect -12060 26359 -12058 26379
rect -12023 26374 -12020 26379
rect -12012 26374 -12010 26379
rect -12013 26360 -12010 26374
rect -11916 26376 -11914 26379
rect -11916 26359 -11913 26376
rect -11892 26359 -11890 26379
rect -11844 26359 -11842 26379
rect -11796 26359 -11794 26379
rect -11676 26359 -11674 26379
rect -11580 26359 -11578 26379
rect -11556 26359 -11554 26379
rect -11484 26360 -11482 26379
rect -11519 26359 -11461 26360
rect -11460 26359 -11458 26379
rect -11436 26359 -11434 26379
rect -11388 26359 -11386 26379
rect -11364 26359 -11362 26379
rect -11340 26359 -11338 26379
rect -11268 26359 -11266 26379
rect -11172 26359 -11170 26379
rect -11124 26359 -11122 26379
rect -11076 26359 -11074 26379
rect -11028 26359 -11026 26379
rect -10788 26359 -10786 26379
rect -10668 26359 -10666 26379
rect -9876 26359 -9874 26379
rect -9828 26359 -9826 26379
rect -9732 26359 -9730 26379
rect -9708 26359 -9706 26379
rect -9612 26359 -9610 26379
rect -9516 26359 -9514 26379
rect -9468 26359 -9466 26379
rect -9420 26359 -9418 26379
rect -9396 26359 -9394 26379
rect -9372 26359 -9370 26379
rect -9300 26359 -9298 26379
rect -9252 26359 -9250 26379
rect -9132 26359 -9130 26379
rect -9084 26359 -9082 26379
rect -9036 26359 -9034 26379
rect -8988 26359 -8986 26379
rect -8940 26359 -8938 26379
rect -8892 26359 -8890 26379
rect -8844 26359 -8842 26379
rect -8807 26374 -8804 26379
rect -8796 26374 -8794 26379
rect -8797 26360 -8794 26374
rect -8700 26376 -8698 26379
rect -8700 26359 -8697 26376
rect -8604 26359 -8602 26379
rect -8508 26359 -8506 26379
rect -8484 26359 -8482 26379
rect -8388 26359 -8386 26379
rect -8364 26359 -8362 26379
rect -8340 26359 -8338 26379
rect -8292 26359 -8290 26379
rect -8268 26359 -8266 26379
rect -8196 26359 -8194 26379
rect -8100 26359 -8098 26379
rect -8052 26359 -8050 26379
rect -7932 26359 -7930 26379
rect -7836 26359 -7834 26379
rect -7740 26359 -7738 26379
rect -7692 26359 -7690 26379
rect -7620 26359 -7618 26379
rect -7404 26359 -7402 26379
rect -7356 26359 -7354 26379
rect -7308 26359 -7306 26379
rect -7212 26359 -7210 26379
rect -7188 26359 -7186 26379
rect -7116 26359 -7114 26379
rect -7068 26359 -7066 26379
rect -6972 26359 -6970 26379
rect -6948 26359 -6946 26379
rect -6876 26359 -6874 26379
rect -6852 26359 -6850 26379
rect -6804 26359 -6802 26379
rect -6780 26359 -6778 26379
rect -6756 26359 -6754 26379
rect -6708 26359 -6706 26379
rect -6684 26359 -6682 26379
rect -6660 26359 -6658 26379
rect -6612 26359 -6610 26379
rect -6588 26359 -6586 26379
rect -6564 26359 -6562 26379
rect -6516 26359 -6514 26379
rect -6492 26359 -6490 26379
rect -6468 26359 -6466 26379
rect -6420 26359 -6418 26379
rect -6396 26359 -6394 26379
rect -6372 26359 -6370 26379
rect -6324 26359 -6322 26379
rect -6300 26359 -6298 26379
rect -6276 26359 -6274 26379
rect -6228 26359 -6226 26379
rect -6180 26359 -6178 26379
rect -6060 26359 -6058 26379
rect -5964 26359 -5962 26379
rect -5940 26359 -5938 26379
rect -5868 26359 -5866 26379
rect -5652 26359 -5650 26379
rect -5316 26359 -5314 26379
rect -5268 26359 -5266 26379
rect -5196 26359 -5194 26379
rect -5172 26359 -5170 26379
rect -5100 26359 -5098 26379
rect -5076 26359 -5074 26379
rect -4980 26359 -4978 26379
rect -4956 26359 -4954 26379
rect -4884 26359 -4882 26379
rect -4860 26359 -4858 26379
rect -4788 26359 -4786 26379
rect -4692 26359 -4690 26379
rect -4644 26359 -4642 26379
rect -4596 26359 -4594 26379
rect -4548 26359 -4546 26379
rect -4428 26359 -4426 26379
rect -4332 26359 -4330 26379
rect -4308 26359 -4306 26379
rect -4260 26359 -4258 26379
rect -4212 26359 -4210 26379
rect -4116 26359 -4114 26379
rect -4092 26359 -4090 26379
rect -4020 26359 -4018 26379
rect -3876 26359 -3874 26379
rect -3732 26359 -3730 26379
rect -3588 26359 -3586 26379
rect -3564 26359 -3562 26379
rect -3516 26359 -3514 26379
rect -3492 26359 -3490 26379
rect -3468 26359 -3466 26379
rect -3420 26359 -3418 26379
rect -3324 26359 -3322 26379
rect -3252 26359 -3250 26379
rect -3228 26359 -3226 26379
rect -3156 26359 -3154 26379
rect -3132 26359 -3130 26379
rect -3060 26359 -3058 26379
rect -3012 26359 -3010 26379
rect -2964 26359 -2962 26379
rect -2916 26359 -2914 26379
rect -2892 26359 -2890 26379
rect -2820 26359 -2818 26379
rect -2796 26359 -2794 26379
rect -2748 26359 -2746 26379
rect -2700 26359 -2698 26379
rect -2604 26359 -2602 26379
rect -2580 26359 -2578 26379
rect -2364 26359 -2362 26379
rect -2292 26359 -2290 26379
rect -2268 26359 -2266 26379
rect -2244 26359 -2242 26379
rect -2172 26359 -2170 26379
rect -2148 26359 -2146 26379
rect -2076 26359 -2074 26379
rect -2052 26359 -2050 26379
rect -1980 26359 -1978 26379
rect -1884 26359 -1882 26379
rect -1836 26359 -1834 26379
rect -1716 26359 -1714 26379
rect -1596 26359 -1594 26379
rect -1476 26359 -1474 26379
rect -1380 26359 -1378 26379
rect -1356 26359 -1354 26379
rect -1308 26359 -1306 26379
rect -1260 26359 -1258 26379
rect -1140 26359 -1138 26379
rect -852 26359 -850 26379
rect -804 26359 -802 26379
rect -756 26359 -754 26379
rect -708 26359 -706 26379
rect -612 26359 -610 26379
rect -588 26359 -586 26379
rect -540 26359 -538 26379
rect -516 26359 -514 26379
rect -492 26359 -490 26379
rect -444 26359 -442 26379
rect -396 26359 -394 26379
rect -300 26359 -298 26379
rect -276 26359 -274 26379
rect -204 26359 -202 26379
rect -108 26359 -106 26379
rect 12 26359 14 26379
rect 108 26359 110 26379
rect 156 26359 158 26379
rect 204 26359 206 26379
rect 228 26359 230 26379
rect 252 26359 254 26379
rect 348 26359 350 26379
rect 468 26359 470 26379
rect 492 26359 494 26379
rect 564 26359 566 26379
rect 588 26359 590 26379
rect 636 26359 638 26379
rect 660 26359 662 26379
rect 684 26359 686 26379
rect 732 26359 734 26379
rect 756 26359 758 26379
rect 780 26359 782 26379
rect 876 26359 878 26379
rect 972 26359 974 26379
rect 1020 26359 1022 26379
rect 1068 26359 1070 26379
rect 1092 26359 1094 26379
rect 1116 26359 1118 26379
rect 1164 26359 1166 26379
rect 1212 26359 1214 26379
rect 1308 26359 1310 26379
rect 1332 26359 1334 26379
rect 1380 26359 1382 26379
rect 1428 26359 1430 26379
rect 1524 26359 1526 26379
rect 1548 26359 1550 26379
rect 1596 26359 1598 26379
rect 1620 26359 1622 26379
rect 1644 26359 1646 26379
rect 1692 26359 1694 26379
rect 1716 26359 1718 26379
rect 1740 26359 1742 26379
rect 1788 26359 1790 26379
rect 1836 26359 1838 26379
rect 1884 26359 1886 26379
rect 1932 26359 1934 26379
rect 1980 26359 1982 26379
rect 2028 26359 2030 26379
rect 2076 26359 2078 26379
rect 2100 26359 2102 26379
rect 2124 26359 2126 26379
rect 2172 26359 2174 26379
rect 2196 26359 2198 26379
rect 2220 26359 2222 26379
rect 2268 26359 2270 26379
rect 2292 26359 2294 26379
rect 2316 26359 2318 26379
rect 2364 26359 2366 26379
rect 2412 26359 2414 26379
rect 2460 26359 2462 26379
rect 2508 26359 2510 26379
rect 2556 26359 2558 26379
rect 2580 26359 2582 26379
rect 2604 26359 2606 26379
rect 2652 26359 2654 26379
rect 2676 26359 2678 26379
rect 2700 26359 2702 26379
rect 2748 26359 2750 26379
rect 2772 26359 2774 26379
rect 2796 26359 2798 26379
rect 2844 26359 2846 26379
rect 2868 26359 2870 26379
rect 2892 26359 2894 26379
rect 2940 26359 2942 26379
rect 3012 26359 3014 26379
rect 3108 26359 3110 26379
rect 3156 26359 3158 26379
rect 3252 26359 3254 26379
rect 3348 26359 3350 26379
rect 3396 26359 3398 26379
rect 3468 26359 3470 26379
rect 3492 26359 3494 26379
rect 3588 26359 3590 26379
rect 3612 26359 3614 26379
rect 3636 26359 3638 26379
rect 3708 26359 3710 26379
rect 3732 26359 3734 26379
rect 3804 26359 3806 26379
rect 3828 26359 3830 26379
rect 3924 26359 3926 26379
rect 4020 26359 4022 26379
rect 4044 26359 4046 26379
rect 4092 26359 4094 26379
rect 4116 26359 4118 26379
rect 4140 26359 4142 26379
rect 4188 26359 4190 26379
rect 4212 26359 4214 26379
rect 4236 26359 4238 26379
rect 4308 26359 4310 26379
rect 4332 26359 4334 26379
rect 4404 26359 4406 26379
rect 4500 26359 4502 26379
rect 4596 26359 4598 26379
rect 4860 26359 4862 26379
rect 4956 26359 4958 26379
rect 4980 26359 4982 26379
rect 5004 26359 5006 26379
rect 5076 26359 5078 26379
rect 5100 26359 5102 26379
rect 5124 26359 5126 26379
rect 5172 26359 5174 26379
rect 5196 26359 5198 26379
rect 5220 26359 5222 26379
rect 5268 26359 5270 26379
rect 5292 26359 5294 26379
rect 5388 26359 5390 26379
rect 5484 26359 5486 26379
rect 5508 26359 5510 26379
rect 5532 26359 5534 26379
rect 5580 26359 5582 26379
rect 5628 26359 5630 26379
rect 5713 26374 5716 26379
rect 5724 26374 5726 26379
rect 5723 26360 5726 26374
rect 5748 26359 5750 26379
rect 5796 26359 5798 26379
rect 5820 26376 5822 26379
rect 5820 26359 5823 26376
rect 5844 26359 5846 26379
rect 5892 26359 5894 26379
rect 6132 26359 6134 26379
rect 6180 26359 6182 26379
rect 6228 26359 6230 26379
rect 6252 26359 6254 26379
rect 6276 26359 6278 26379
rect 6324 26359 6326 26379
rect 6372 26359 6374 26379
rect 6492 26359 6494 26379
rect 6588 26359 6590 26379
rect 6612 26359 6614 26379
rect 6660 26359 6662 26379
rect 6684 26359 6686 26379
rect 6708 26359 6710 26379
rect 6780 26359 6782 26379
rect 6804 26359 6806 26379
rect 6828 26359 6830 26379
rect 6900 26359 6902 26379
rect 6924 26359 6926 26379
rect 7020 26359 7022 26379
rect 7140 26359 7142 26379
rect 7236 26359 7238 26379
rect 7332 26359 7334 26379
rect 7380 26359 7382 26379
rect 7428 26359 7430 26379
rect 7452 26359 7454 26379
rect 7476 26359 7478 26379
rect 7524 26359 7526 26379
rect 7548 26359 7550 26379
rect 7572 26359 7574 26379
rect 7620 26359 7622 26379
rect 7644 26359 7646 26379
rect 7668 26359 7670 26379
rect 7716 26359 7718 26379
rect 7740 26359 7742 26379
rect 7836 26359 7838 26379
rect 7884 26359 7886 26379
rect 7932 26359 7934 26379
rect 7956 26359 7958 26379
rect 7980 26359 7982 26379
rect 8052 26359 8054 26379
rect 8148 26359 8150 26379
rect 8196 26359 8198 26379
rect 8244 26359 8246 26379
rect 8268 26359 8270 26379
rect 8292 26359 8294 26379
rect 8340 26359 8342 26379
rect 8364 26359 8366 26379
rect 8388 26359 8390 26379
rect 8436 26359 8438 26379
rect 8460 26359 8462 26379
rect 8556 26359 8558 26379
rect 8604 26359 8606 26379
rect 8652 26359 8654 26379
rect 8700 26359 8702 26379
rect 8724 26359 8726 26379
rect 8748 26359 8750 26379
rect 8820 26359 8822 26379
rect 8844 26359 8846 26379
rect 8868 26359 8870 26379
rect 9516 26359 9518 26379
rect 9612 26359 9614 26379
rect 9660 26359 9662 26379
rect 9684 26359 9686 26379
rect 9708 26359 9710 26379
rect 9756 26359 9758 26379
rect 9780 26359 9782 26379
rect 9804 26359 9806 26379
rect 9852 26359 9854 26379
rect 9876 26359 9878 26379
rect 9900 26359 9902 26379
rect 9948 26359 9950 26379
rect 9972 26359 9974 26379
rect 9996 26359 9998 26379
rect 10068 26359 10070 26379
rect 10092 26359 10094 26379
rect 10116 26359 10118 26379
rect 10164 26359 10166 26379
rect 10188 26359 10190 26379
rect 10212 26359 10214 26379
rect 10260 26359 10262 26379
rect 10284 26359 10286 26379
rect 10308 26359 10310 26379
rect 10380 26359 10382 26379
rect 10404 26359 10406 26379
rect 10428 26359 10430 26379
rect 10476 26359 10478 26379
rect 10500 26359 10502 26379
rect 10524 26359 10526 26379
rect 10572 26359 10574 26379
rect 10596 26359 10598 26379
rect 10620 26359 10622 26379
rect 10668 26359 10670 26379
rect 10692 26359 10694 26379
rect 10716 26359 10718 26379
rect 10788 26359 10790 26379
rect 10836 26359 10838 26379
rect 10956 26359 10958 26379
rect 11052 26359 11054 26379
rect 11076 26359 11078 26379
rect 11124 26359 11126 26379
rect 11172 26359 11174 26379
rect 11220 26359 11222 26379
rect 11340 26359 11342 26379
rect 11436 26359 11438 26379
rect 11532 26359 11534 26379
rect 11580 26359 11582 26379
rect 11628 26359 11630 26379
rect 11676 26359 11678 26379
rect 11772 26359 11774 26379
rect 11796 26359 11798 26379
rect 11844 26359 11846 26379
rect 11892 26359 11894 26379
rect 11988 26359 11990 26379
rect 12060 26359 12062 26379
rect 12132 26359 12134 26379
rect 12169 26359 12227 26360
rect 12228 26359 12230 26379
rect 12324 26359 12326 26379
rect 12420 26359 12422 26379
rect 12444 26359 12446 26379
rect 12492 26359 12494 26379
rect 12516 26359 12518 26379
rect 12540 26359 12542 26379
rect 12588 26359 12590 26379
rect 12636 26359 12638 26379
rect 12732 26359 12734 26379
rect 12756 26359 12758 26379
rect 12804 26359 12806 26379
rect 12828 26359 12830 26379
rect 12852 26359 12854 26379
rect 12900 26359 12902 26379
rect 12948 26359 12950 26379
rect 13044 26359 13046 26379
rect 13068 26359 13070 26379
rect 13116 26359 13118 26379
rect 13284 26359 13286 26379
rect 13332 26359 13334 26379
rect 13428 26359 13430 26379
rect 13524 26359 13526 26379
rect 13572 26359 13574 26379
rect 13644 26359 13646 26379
rect 13668 26359 13670 26379
rect 13764 26359 13766 26379
rect 13812 26359 13814 26379
rect 13860 26359 13862 26379
rect 13908 26359 13910 26379
rect 13956 26359 13958 26379
rect 14004 26359 14006 26379
rect 14100 26359 14102 26379
rect 14196 26359 14198 26379
rect 14244 26359 14246 26379
rect 14292 26359 14294 26379
rect 15132 26359 15134 26379
rect 15228 26359 15230 26379
rect 15252 26359 15254 26379
rect 15300 26359 15302 26379
rect 15324 26359 15326 26379
rect 15396 26359 15398 26379
rect 15420 26359 15422 26379
rect 15492 26359 15494 26379
rect 15540 26359 15542 26379
rect 15636 26359 15638 26379
rect 15660 26359 15662 26379
rect 15708 26359 15710 26379
rect 15732 26359 15734 26379
rect 15756 26359 15758 26379
rect 15804 26359 15806 26379
rect 15828 26359 15830 26379
rect 15852 26359 15854 26379
rect 15900 26359 15902 26379
rect 15948 26359 15950 26379
rect 15996 26359 15998 26379
rect 16044 26359 16046 26379
rect 16092 26359 16094 26379
rect 16140 26359 16142 26379
rect 16236 26359 16238 26379
rect 16260 26359 16262 26379
rect 16308 26359 16310 26379
rect 16332 26359 16334 26379
rect 16356 26359 16358 26379
rect 16404 26359 16406 26379
rect 16452 26359 16454 26379
rect 16548 26359 16550 26379
rect 16572 26359 16574 26379
rect 16620 26359 16622 26379
rect 16668 26359 16670 26379
rect 16716 26359 16718 26379
rect 16764 26359 16766 26379
rect 16836 26359 16838 26379
rect 16884 26359 16886 26379
rect 16980 26359 16982 26379
rect 17052 26359 17054 26379
rect 17196 26359 17198 26379
rect 17220 26359 17222 26379
rect 17292 26359 17294 26379
rect 17316 26359 17318 26379
rect 18084 26359 18086 26379
rect 18132 26359 18134 26379
rect 18396 26359 18398 26379
rect 18492 26359 18494 26379
rect 18516 26359 18518 26379
rect 18564 26359 18566 26379
rect 18612 26359 18614 26379
rect 18660 26359 18662 26379
rect 18708 26359 18710 26379
rect 18756 26359 18758 26379
rect 18804 26359 18806 26379
rect 18852 26359 18854 26379
rect 18900 26359 18902 26379
rect 18996 26359 18998 26379
rect 19020 26359 19022 26379
rect 19092 26359 19094 26379
rect 19116 26359 19118 26379
rect 19140 26359 19142 26379
rect 19188 26359 19190 26379
rect 19236 26359 19238 26379
rect 19332 26359 19334 26379
rect 19476 26359 19478 26379
rect 19620 26359 19622 26379
rect 19716 26359 19718 26379
rect 19788 26359 19790 26379
rect 19836 26359 19838 26379
rect 19860 26359 19862 26379
rect 19884 26359 19886 26379
rect 19932 26359 19934 26379
rect 19956 26359 19958 26379
rect 19980 26359 19982 26379
rect 20028 26359 20030 26379
rect 20052 26359 20054 26379
rect 20076 26359 20078 26379
rect 20148 26359 20150 26379
rect 20172 26359 20174 26379
rect 20196 26359 20198 26379
rect 20268 26359 20270 26379
rect 20292 26359 20294 26379
rect 20388 26359 20390 26379
rect 20412 26359 20414 26379
rect 20508 26359 20510 26379
rect 20556 26359 20558 26379
rect 20604 26359 20606 26379
rect 20916 26359 20918 26379
rect 20964 26359 20966 26379
rect 21012 26359 21014 26379
rect 21060 26359 21062 26379
rect 21084 26359 21086 26379
rect 21108 26359 21110 26379
rect 21204 26359 21206 26379
rect 21300 26359 21302 26379
rect 21324 26359 21326 26379
rect 21444 26359 21446 26379
rect 21468 26359 21470 26379
rect 21564 26359 21566 26379
rect 21612 26359 21614 26379
rect 21684 26359 21686 26379
rect 21708 26359 21710 26379
rect 21804 26359 21806 26379
rect 21828 26359 21830 26379
rect 21924 26359 21926 26379
rect 21948 26359 21950 26379
rect 22044 26359 22046 26379
rect 22068 26359 22070 26379
rect 22188 26359 22190 26379
rect 22212 26359 22214 26379
rect 23004 26359 23006 26379
rect 23052 26359 23054 26379
rect 23076 26359 23078 26379
rect 23100 26359 23102 26379
rect 23148 26359 23150 26379
rect 23220 26359 23222 26379
rect 23244 26359 23246 26379
rect 23316 26359 23318 26379
rect 23340 26359 23342 26379
rect 23412 26359 23414 26379
rect 23556 26359 23558 26379
rect 23628 26359 23630 26379
rect 23652 26359 23654 26379
rect 23676 26359 23678 26379
rect 23724 26359 23726 26379
rect 23772 26359 23774 26379
rect 23820 26359 23822 26379
rect 23868 26359 23870 26379
rect 23916 26359 23918 26379
rect 24012 26359 24014 26379
rect 24084 26359 24086 26379
rect 24372 26359 24374 26379
rect 24396 26359 24398 26379
rect 24492 26359 24494 26379
rect 24516 26359 24518 26379
rect 24588 26359 24590 26379
rect 24612 26359 24614 26379
rect 24708 26359 24710 26379
rect 24732 26359 24734 26379
rect 24756 26359 24758 26379
rect 24852 26359 24854 26379
rect 24876 26359 24878 26379
rect 24972 26359 24974 26379
rect 24996 26359 24998 26379
rect 25092 26359 25094 26379
rect 25260 26359 25262 26379
rect 25356 26359 25358 26379
rect 25380 26359 25382 26379
rect 25452 26359 25454 26379
rect 25465 26374 25468 26379
rect 25476 26374 25478 26379
rect 25475 26360 25478 26374
rect 25500 26359 25502 26379
rect 25572 26376 25574 26379
rect 25572 26359 25575 26376
rect 25596 26359 25598 26379
rect 27060 26359 27062 26379
rect 27108 26359 27110 26379
rect 27180 26359 27182 26379
rect 27324 26359 27326 26379
rect 27396 26359 27398 26379
rect 27420 26359 27422 26379
rect 27540 26359 27542 26379
rect 27564 26359 27566 26379
rect 30564 26359 30566 26379
rect 30636 26359 30638 26379
rect 30660 26359 30662 26379
rect 30780 26359 30782 26379
rect 30804 26359 30806 26379
rect 30924 26359 30926 26379
rect 30948 26359 30950 26379
rect 31068 26359 31070 26379
rect 31092 26359 31094 26379
rect 31164 26360 31166 26379
rect 31236 26360 31238 26379
rect 31129 26359 31187 26360
rect 31225 26359 31259 26360
rect -18273 26355 -17899 26359
rect -18273 26352 -18259 26355
rect -18108 26352 -18106 26355
rect -18191 26342 -18187 26350
rect -18201 26336 -18191 26342
rect -18108 26335 -18105 26352
rect -17940 26335 -17938 26355
rect -17913 26352 -17899 26355
rect -17889 26355 -16651 26359
rect -17889 26352 -17875 26355
rect -17817 26352 -17803 26355
rect -17735 26350 -17732 26355
rect -17604 26352 -17602 26355
rect -17725 26336 -17722 26350
rect -17855 26335 -17797 26336
rect -17724 26335 -17722 26336
rect -17628 26335 -17625 26352
rect -17604 26335 -17601 26352
rect -17532 26335 -17530 26355
rect -17460 26335 -17458 26355
rect -17436 26335 -17434 26355
rect -17292 26335 -17290 26355
rect -17241 26352 -17227 26355
rect -17196 26335 -17194 26355
rect -17028 26335 -17026 26355
rect -16860 26335 -16858 26355
rect -16823 26350 -16820 26355
rect -16812 26350 -16810 26355
rect -16813 26336 -16810 26350
rect -16764 26335 -16762 26355
rect -16716 26352 -16714 26355
rect -16740 26335 -16737 26352
rect -16716 26335 -16713 26352
rect -16668 26335 -16666 26355
rect -16665 26352 -16651 26355
rect -16617 26355 -16171 26359
rect -16617 26352 -16603 26355
rect -16596 26352 -16593 26355
rect -16500 26335 -16498 26355
rect -16380 26335 -16378 26355
rect -16356 26335 -16354 26355
rect -16329 26352 -16315 26355
rect -16308 26352 -16305 26355
rect -16260 26335 -16258 26355
rect -16236 26335 -16234 26355
rect -16212 26335 -16210 26355
rect -16185 26352 -16171 26355
rect -16113 26355 31259 26359
rect -16113 26352 -16099 26355
rect -15300 26335 -15298 26355
rect -15084 26335 -15082 26355
rect -15036 26335 -15034 26355
rect -14868 26335 -14866 26355
rect -14772 26335 -14770 26355
rect -14724 26335 -14722 26355
rect -14508 26335 -14506 26355
rect -14436 26335 -14434 26355
rect -14388 26335 -14386 26355
rect -14172 26335 -14170 26355
rect -14076 26335 -14074 26355
rect -14028 26352 -14026 26355
rect -14028 26335 -14025 26352
rect -13980 26335 -13978 26355
rect -13932 26335 -13930 26355
rect -13881 26352 -13867 26355
rect -13860 26352 -13857 26355
rect -13895 26335 -13837 26336
rect -13764 26335 -13762 26355
rect -13716 26335 -13714 26355
rect -13644 26335 -13642 26355
rect -13596 26335 -13594 26355
rect -13500 26335 -13498 26355
rect -13404 26335 -13402 26355
rect -13356 26335 -13354 26355
rect -13284 26335 -13282 26355
rect -13068 26335 -13066 26355
rect -12828 26335 -12826 26355
rect -12780 26335 -12778 26355
rect -12660 26335 -12658 26355
rect -12564 26335 -12562 26355
rect -12492 26335 -12490 26355
rect -12396 26335 -12394 26355
rect -12348 26335 -12346 26355
rect -12276 26335 -12274 26355
rect -12252 26335 -12250 26355
rect -12156 26335 -12154 26355
rect -12060 26335 -12058 26355
rect -11937 26352 -11923 26355
rect -11916 26352 -11913 26355
rect -11892 26335 -11890 26355
rect -11844 26335 -11842 26355
rect -11796 26335 -11794 26355
rect -11676 26335 -11674 26355
rect -11580 26335 -11578 26355
rect -11556 26335 -11554 26355
rect -11519 26350 -11516 26355
rect -11495 26350 -11492 26355
rect -11484 26350 -11482 26355
rect -11509 26336 -11506 26350
rect -11485 26336 -11482 26350
rect -11508 26335 -11506 26336
rect -11460 26335 -11458 26355
rect -11436 26335 -11434 26355
rect -11388 26352 -11386 26355
rect -11388 26335 -11385 26352
rect -11364 26335 -11362 26355
rect -11340 26335 -11338 26355
rect -11268 26335 -11266 26355
rect -11172 26335 -11170 26355
rect -11124 26335 -11122 26355
rect -11076 26335 -11074 26355
rect -11028 26335 -11026 26355
rect -10788 26335 -10786 26355
rect -10668 26335 -10666 26355
rect -9876 26335 -9874 26355
rect -9828 26335 -9826 26355
rect -9732 26335 -9730 26355
rect -9708 26335 -9706 26355
rect -9612 26335 -9610 26355
rect -9516 26335 -9514 26355
rect -9468 26335 -9466 26355
rect -9420 26335 -9418 26355
rect -9396 26335 -9394 26355
rect -9372 26335 -9370 26355
rect -9300 26335 -9298 26355
rect -9252 26335 -9250 26355
rect -9132 26335 -9130 26355
rect -9084 26335 -9082 26355
rect -9036 26335 -9034 26355
rect -8988 26335 -8986 26355
rect -8940 26335 -8938 26355
rect -8892 26335 -8890 26355
rect -8844 26335 -8842 26355
rect -8721 26352 -8707 26355
rect -8700 26352 -8697 26355
rect -8604 26335 -8602 26355
rect -8508 26335 -8506 26355
rect -8484 26335 -8482 26355
rect -8388 26335 -8386 26355
rect -8364 26335 -8362 26355
rect -8340 26335 -8338 26355
rect -8292 26335 -8290 26355
rect -8268 26335 -8266 26355
rect -8196 26335 -8194 26355
rect -8100 26335 -8098 26355
rect -8052 26335 -8050 26355
rect -7932 26335 -7930 26355
rect -7836 26335 -7834 26355
rect -7740 26335 -7738 26355
rect -7692 26335 -7690 26355
rect -7620 26335 -7618 26355
rect -7404 26335 -7402 26355
rect -7356 26335 -7354 26355
rect -7308 26335 -7306 26355
rect -7212 26335 -7210 26355
rect -7188 26335 -7186 26355
rect -7116 26335 -7114 26355
rect -7068 26335 -7066 26355
rect -6972 26335 -6970 26355
rect -6948 26335 -6946 26355
rect -6876 26335 -6874 26355
rect -6852 26335 -6850 26355
rect -6804 26335 -6802 26355
rect -6780 26335 -6778 26355
rect -6756 26335 -6754 26355
rect -6708 26335 -6706 26355
rect -6684 26335 -6682 26355
rect -6660 26335 -6658 26355
rect -6612 26335 -6610 26355
rect -6588 26335 -6586 26355
rect -6564 26335 -6562 26355
rect -6516 26335 -6514 26355
rect -6492 26335 -6490 26355
rect -6468 26335 -6466 26355
rect -6420 26335 -6418 26355
rect -6396 26335 -6394 26355
rect -6372 26335 -6370 26355
rect -6324 26335 -6322 26355
rect -6300 26335 -6298 26355
rect -6276 26335 -6274 26355
rect -6228 26335 -6226 26355
rect -6180 26335 -6178 26355
rect -6060 26335 -6058 26355
rect -5964 26336 -5962 26355
rect -5999 26335 -5941 26336
rect -5940 26335 -5938 26355
rect -5868 26335 -5866 26355
rect -5652 26335 -5650 26355
rect -5316 26335 -5314 26355
rect -5268 26335 -5266 26355
rect -5196 26335 -5194 26355
rect -5172 26335 -5170 26355
rect -5100 26335 -5098 26355
rect -5076 26335 -5074 26355
rect -4980 26335 -4978 26355
rect -4956 26335 -4954 26355
rect -4884 26335 -4882 26355
rect -4860 26335 -4858 26355
rect -4788 26335 -4786 26355
rect -4692 26335 -4690 26355
rect -4644 26335 -4642 26355
rect -4596 26335 -4594 26355
rect -4548 26335 -4546 26355
rect -4428 26335 -4426 26355
rect -4332 26335 -4330 26355
rect -4308 26335 -4306 26355
rect -4260 26335 -4258 26355
rect -4212 26335 -4210 26355
rect -4116 26335 -4114 26355
rect -4092 26335 -4090 26355
rect -4020 26335 -4018 26355
rect -3876 26335 -3874 26355
rect -3732 26335 -3730 26355
rect -3588 26335 -3586 26355
rect -3564 26335 -3562 26355
rect -3516 26335 -3514 26355
rect -3492 26335 -3490 26355
rect -3468 26335 -3466 26355
rect -3420 26335 -3418 26355
rect -3324 26335 -3322 26355
rect -3252 26335 -3250 26355
rect -3228 26335 -3226 26355
rect -3156 26335 -3154 26355
rect -3132 26335 -3130 26355
rect -3060 26335 -3058 26355
rect -3012 26335 -3010 26355
rect -2964 26335 -2962 26355
rect -2916 26335 -2914 26355
rect -2892 26335 -2890 26355
rect -2820 26335 -2818 26355
rect -2796 26335 -2794 26355
rect -2748 26335 -2746 26355
rect -2700 26335 -2698 26355
rect -2604 26335 -2602 26355
rect -2580 26335 -2578 26355
rect -2364 26335 -2362 26355
rect -2292 26335 -2290 26355
rect -2268 26335 -2266 26355
rect -2244 26335 -2242 26355
rect -2172 26335 -2170 26355
rect -2148 26335 -2146 26355
rect -2076 26335 -2074 26355
rect -2052 26335 -2050 26355
rect -1980 26335 -1978 26355
rect -1884 26335 -1882 26355
rect -1836 26335 -1834 26355
rect -1716 26335 -1714 26355
rect -1679 26335 -1621 26336
rect -1596 26335 -1594 26355
rect -1476 26335 -1474 26355
rect -1380 26335 -1378 26355
rect -1356 26335 -1354 26355
rect -1308 26335 -1306 26355
rect -1260 26335 -1258 26355
rect -1140 26335 -1138 26355
rect -852 26335 -850 26355
rect -804 26335 -802 26355
rect -756 26335 -754 26355
rect -708 26335 -706 26355
rect -612 26335 -610 26355
rect -588 26335 -586 26355
rect -540 26335 -538 26355
rect -516 26335 -514 26355
rect -492 26335 -490 26355
rect -444 26335 -442 26355
rect -396 26335 -394 26355
rect -300 26335 -298 26355
rect -276 26335 -274 26355
rect -204 26335 -202 26355
rect -108 26335 -106 26355
rect 12 26335 14 26355
rect 108 26335 110 26355
rect 156 26335 158 26355
rect 204 26335 206 26355
rect 228 26335 230 26355
rect 252 26335 254 26355
rect 348 26335 350 26355
rect 468 26335 470 26355
rect 492 26335 494 26355
rect 564 26335 566 26355
rect 588 26335 590 26355
rect 636 26335 638 26355
rect 660 26335 662 26355
rect 684 26336 686 26355
rect 673 26335 707 26336
rect 732 26335 734 26355
rect 756 26335 758 26355
rect 780 26335 782 26355
rect 876 26335 878 26355
rect 972 26335 974 26355
rect 1020 26335 1022 26355
rect 1068 26335 1070 26355
rect 1092 26335 1094 26355
rect 1116 26335 1118 26355
rect 1164 26335 1166 26355
rect 1212 26335 1214 26355
rect 1308 26335 1310 26355
rect 1332 26335 1334 26355
rect 1380 26335 1382 26355
rect 1428 26335 1430 26355
rect 1524 26335 1526 26355
rect 1548 26335 1550 26355
rect 1596 26335 1598 26355
rect 1620 26335 1622 26355
rect 1644 26335 1646 26355
rect 1692 26335 1694 26355
rect 1716 26335 1718 26355
rect 1740 26335 1742 26355
rect 1788 26335 1790 26355
rect 1836 26336 1838 26355
rect 1825 26335 1859 26336
rect 1884 26335 1886 26355
rect 1932 26335 1934 26355
rect 1980 26335 1982 26355
rect 2028 26335 2030 26355
rect 2076 26335 2078 26355
rect 2100 26335 2102 26355
rect 2124 26335 2126 26355
rect 2172 26335 2174 26355
rect 2196 26335 2198 26355
rect 2220 26335 2222 26355
rect 2268 26335 2270 26355
rect 2292 26335 2294 26355
rect 2316 26335 2318 26355
rect 2364 26335 2366 26355
rect 2412 26335 2414 26355
rect 2460 26335 2462 26355
rect 2508 26335 2510 26355
rect 2556 26335 2558 26355
rect 2580 26335 2582 26355
rect 2604 26335 2606 26355
rect 2652 26335 2654 26355
rect 2676 26335 2678 26355
rect 2700 26335 2702 26355
rect 2748 26335 2750 26355
rect 2772 26335 2774 26355
rect 2796 26335 2798 26355
rect 2844 26335 2846 26355
rect 2868 26335 2870 26355
rect 2892 26335 2894 26355
rect 2940 26335 2942 26355
rect 3012 26335 3014 26355
rect 3108 26335 3110 26355
rect 3156 26335 3158 26355
rect 3252 26335 3254 26355
rect 3348 26335 3350 26355
rect 3396 26335 3398 26355
rect 3468 26335 3470 26355
rect 3492 26335 3494 26355
rect 3588 26335 3590 26355
rect 3612 26335 3614 26355
rect 3636 26335 3638 26355
rect 3708 26335 3710 26355
rect 3732 26335 3734 26355
rect 3804 26335 3806 26355
rect 3828 26335 3830 26355
rect 3924 26335 3926 26355
rect 4020 26335 4022 26355
rect 4044 26335 4046 26355
rect 4092 26335 4094 26355
rect 4116 26335 4118 26355
rect 4140 26335 4142 26355
rect 4188 26335 4190 26355
rect 4212 26335 4214 26355
rect 4236 26335 4238 26355
rect 4308 26335 4310 26355
rect 4332 26335 4334 26355
rect 4404 26335 4406 26355
rect 4500 26335 4502 26355
rect 4596 26335 4598 26355
rect 4860 26335 4862 26355
rect 4956 26335 4958 26355
rect 4980 26335 4982 26355
rect 5004 26335 5006 26355
rect 5076 26335 5078 26355
rect 5100 26335 5102 26355
rect 5124 26335 5126 26355
rect 5172 26335 5174 26355
rect 5196 26335 5198 26355
rect 5220 26335 5222 26355
rect 5268 26335 5270 26355
rect 5292 26335 5294 26355
rect 5388 26335 5390 26355
rect 5484 26335 5486 26355
rect 5508 26335 5510 26355
rect 5532 26335 5534 26355
rect 5580 26336 5582 26355
rect 5545 26335 5603 26336
rect 5628 26335 5630 26355
rect 5748 26335 5750 26355
rect 5796 26335 5798 26355
rect 5799 26352 5813 26355
rect 5820 26352 5823 26355
rect 5844 26335 5846 26355
rect 5892 26335 5894 26355
rect 6132 26335 6134 26355
rect 6180 26335 6182 26355
rect 6228 26335 6230 26355
rect 6252 26335 6254 26355
rect 6276 26335 6278 26355
rect 6324 26335 6326 26355
rect 6372 26335 6374 26355
rect 6492 26335 6494 26355
rect 6588 26335 6590 26355
rect 6612 26335 6614 26355
rect 6660 26335 6662 26355
rect 6684 26335 6686 26355
rect 6708 26335 6710 26355
rect 6780 26335 6782 26355
rect 6804 26335 6806 26355
rect 6828 26335 6830 26355
rect 6900 26335 6902 26355
rect 6924 26335 6926 26355
rect 7020 26335 7022 26355
rect 7140 26335 7142 26355
rect 7236 26335 7238 26355
rect 7332 26335 7334 26355
rect 7380 26335 7382 26355
rect 7428 26335 7430 26355
rect 7452 26335 7454 26355
rect 7476 26335 7478 26355
rect 7524 26335 7526 26355
rect 7548 26335 7550 26355
rect 7572 26335 7574 26355
rect 7620 26335 7622 26355
rect 7644 26335 7646 26355
rect 7668 26335 7670 26355
rect 7716 26335 7718 26355
rect 7740 26335 7742 26355
rect 7836 26335 7838 26355
rect 7884 26335 7886 26355
rect 7932 26335 7934 26355
rect 7956 26335 7958 26355
rect 7980 26335 7982 26355
rect 8052 26336 8054 26355
rect 8017 26335 8075 26336
rect 8148 26335 8150 26355
rect 8196 26335 8198 26355
rect 8244 26335 8246 26355
rect 8268 26335 8270 26355
rect 8292 26335 8294 26355
rect 8340 26335 8342 26355
rect 8364 26335 8366 26355
rect 8388 26335 8390 26355
rect 8436 26335 8438 26355
rect 8460 26335 8462 26355
rect 8556 26335 8558 26355
rect 8604 26335 8606 26355
rect 8652 26335 8654 26355
rect 8700 26335 8702 26355
rect 8724 26335 8726 26355
rect 8748 26335 8750 26355
rect 8820 26335 8822 26355
rect 8844 26335 8846 26355
rect 8868 26335 8870 26355
rect 9516 26335 9518 26355
rect 9612 26335 9614 26355
rect 9660 26335 9662 26355
rect 9684 26335 9686 26355
rect 9708 26335 9710 26355
rect 9756 26335 9758 26355
rect 9780 26335 9782 26355
rect 9804 26335 9806 26355
rect 9852 26335 9854 26355
rect 9876 26335 9878 26355
rect 9900 26335 9902 26355
rect 9948 26335 9950 26355
rect 9972 26335 9974 26355
rect 9996 26335 9998 26355
rect 10068 26335 10070 26355
rect 10092 26335 10094 26355
rect 10116 26335 10118 26355
rect 10164 26335 10166 26355
rect 10188 26335 10190 26355
rect 10212 26335 10214 26355
rect 10260 26335 10262 26355
rect 10284 26335 10286 26355
rect 10308 26335 10310 26355
rect 10380 26335 10382 26355
rect 10404 26335 10406 26355
rect 10428 26335 10430 26355
rect 10476 26335 10478 26355
rect 10500 26335 10502 26355
rect 10524 26335 10526 26355
rect 10572 26335 10574 26355
rect 10596 26335 10598 26355
rect 10620 26335 10622 26355
rect 10668 26335 10670 26355
rect 10692 26335 10694 26355
rect 10716 26335 10718 26355
rect 10788 26335 10790 26355
rect 10836 26335 10838 26355
rect 10956 26335 10958 26355
rect 11052 26335 11054 26355
rect 11076 26335 11078 26355
rect 11124 26335 11126 26355
rect 11172 26335 11174 26355
rect 11220 26335 11222 26355
rect 11340 26335 11342 26355
rect 11436 26335 11438 26355
rect 11532 26335 11534 26355
rect 11580 26335 11582 26355
rect 11628 26335 11630 26355
rect 11676 26335 11678 26355
rect 11772 26335 11774 26355
rect 11796 26335 11798 26355
rect 11844 26335 11846 26355
rect 11892 26335 11894 26355
rect 11988 26335 11990 26355
rect 12060 26335 12062 26355
rect 12132 26335 12134 26355
rect 12228 26335 12230 26355
rect 12276 26335 12279 26352
rect 12324 26335 12326 26355
rect 12420 26335 12422 26355
rect 12444 26335 12446 26355
rect 12492 26335 12494 26355
rect 12516 26335 12518 26355
rect 12540 26335 12542 26355
rect 12588 26335 12590 26355
rect 12636 26335 12638 26355
rect 12732 26335 12734 26355
rect 12756 26335 12758 26355
rect 12804 26335 12806 26355
rect 12828 26335 12830 26355
rect 12852 26335 12854 26355
rect 12900 26335 12902 26355
rect 12948 26335 12950 26355
rect 13044 26335 13046 26355
rect 13068 26335 13070 26355
rect 13116 26335 13118 26355
rect 13284 26335 13286 26355
rect 13332 26335 13334 26355
rect 13428 26335 13430 26355
rect 13524 26335 13526 26355
rect 13572 26335 13574 26355
rect 13644 26335 13646 26355
rect 13668 26335 13670 26355
rect 13764 26335 13766 26355
rect 13812 26335 13814 26355
rect 13860 26335 13862 26355
rect 13908 26335 13910 26355
rect 13956 26335 13958 26355
rect 14004 26335 14006 26355
rect 14100 26335 14102 26355
rect 14196 26335 14198 26355
rect 14244 26335 14246 26355
rect 14292 26335 14294 26355
rect 15132 26335 15134 26355
rect 15169 26335 15227 26336
rect 15228 26335 15230 26355
rect 15252 26335 15254 26355
rect 15300 26335 15302 26355
rect 15324 26335 15326 26355
rect 15396 26335 15398 26355
rect 15420 26335 15422 26355
rect 15492 26335 15494 26355
rect 15540 26335 15542 26355
rect 15636 26335 15638 26355
rect 15660 26335 15662 26355
rect 15708 26335 15710 26355
rect 15732 26335 15734 26355
rect 15756 26335 15758 26355
rect 15804 26335 15806 26355
rect 15828 26335 15830 26355
rect 15852 26335 15854 26355
rect 15900 26335 15902 26355
rect 15948 26335 15950 26355
rect 15996 26335 15998 26355
rect 16044 26335 16046 26355
rect 16092 26335 16094 26355
rect 16140 26335 16142 26355
rect 16236 26335 16238 26355
rect 16260 26335 16262 26355
rect 16308 26335 16310 26355
rect 16332 26335 16334 26355
rect 16356 26335 16358 26355
rect 16404 26335 16406 26355
rect 16452 26335 16454 26355
rect 16548 26335 16550 26355
rect 16572 26335 16574 26355
rect 16620 26335 16622 26355
rect 16668 26335 16670 26355
rect 16716 26335 16718 26355
rect 16764 26335 16766 26355
rect 16836 26335 16838 26355
rect 16884 26335 16886 26355
rect 16980 26335 16982 26355
rect 17052 26335 17054 26355
rect 17196 26335 17198 26355
rect 17220 26335 17222 26355
rect 17292 26335 17294 26355
rect 17316 26335 17318 26355
rect 18084 26335 18086 26355
rect 18132 26335 18134 26355
rect 18396 26335 18398 26355
rect 18492 26335 18494 26355
rect 18516 26335 18518 26355
rect 18564 26335 18566 26355
rect 18612 26335 18614 26355
rect 18660 26335 18662 26355
rect 18708 26335 18710 26355
rect 18756 26335 18758 26355
rect 18804 26335 18806 26355
rect 18852 26335 18854 26355
rect 18900 26335 18902 26355
rect 18996 26335 18998 26355
rect 19020 26335 19022 26355
rect 19092 26335 19094 26355
rect 19116 26335 19118 26355
rect 19140 26335 19142 26355
rect 19188 26335 19190 26355
rect 19236 26335 19238 26355
rect 19332 26335 19334 26355
rect 19476 26335 19478 26355
rect 19620 26335 19622 26355
rect 19716 26335 19718 26355
rect 19788 26335 19790 26355
rect 19836 26335 19838 26355
rect 19860 26335 19862 26355
rect 19884 26335 19886 26355
rect 19932 26335 19934 26355
rect 19956 26335 19958 26355
rect 19980 26335 19982 26355
rect 20028 26335 20030 26355
rect 20052 26335 20054 26355
rect 20076 26335 20078 26355
rect 20148 26335 20150 26355
rect 20172 26335 20174 26355
rect 20196 26335 20198 26355
rect 20268 26335 20270 26355
rect 20292 26335 20294 26355
rect 20388 26335 20390 26355
rect 20412 26335 20414 26355
rect 20508 26335 20510 26355
rect 20556 26335 20558 26355
rect 20604 26335 20606 26355
rect 20916 26335 20918 26355
rect 20964 26335 20966 26355
rect 21012 26335 21014 26355
rect 21060 26335 21062 26355
rect 21084 26335 21086 26355
rect 21108 26335 21110 26355
rect 21204 26335 21206 26355
rect 21300 26335 21302 26355
rect 21324 26335 21326 26355
rect 21444 26335 21446 26355
rect 21468 26335 21470 26355
rect 21564 26335 21566 26355
rect 21612 26335 21614 26355
rect 21684 26335 21686 26355
rect 21708 26335 21710 26355
rect 21804 26335 21806 26355
rect 21828 26335 21830 26355
rect 21924 26335 21926 26355
rect 21948 26335 21950 26355
rect 22044 26335 22046 26355
rect 22068 26335 22070 26355
rect 22188 26335 22190 26355
rect 22212 26335 22214 26355
rect 23004 26335 23006 26355
rect 23052 26335 23054 26355
rect 23076 26335 23078 26355
rect 23100 26335 23102 26355
rect 23148 26335 23150 26355
rect 23220 26335 23222 26355
rect 23244 26335 23246 26355
rect 23316 26335 23318 26355
rect 23340 26335 23342 26355
rect 23412 26335 23414 26355
rect 23556 26335 23558 26355
rect 23628 26335 23630 26355
rect 23652 26335 23654 26355
rect 23676 26335 23678 26355
rect 23724 26335 23726 26355
rect 23772 26335 23774 26355
rect 23820 26335 23822 26355
rect 23868 26335 23870 26355
rect 23916 26335 23918 26355
rect 24012 26335 24014 26355
rect 24084 26335 24086 26355
rect 24372 26335 24374 26355
rect 24396 26335 24398 26355
rect 24492 26335 24494 26355
rect 24516 26335 24518 26355
rect 24588 26335 24590 26355
rect 24612 26335 24614 26355
rect 24708 26335 24710 26355
rect 24732 26335 24734 26355
rect 24756 26335 24758 26355
rect 24852 26335 24854 26355
rect 24876 26335 24878 26355
rect 24972 26335 24974 26355
rect 24996 26335 24998 26355
rect 25092 26335 25094 26355
rect 25260 26335 25262 26355
rect 25356 26335 25358 26355
rect 25380 26335 25382 26355
rect 25452 26335 25454 26355
rect 25500 26335 25502 26355
rect 25551 26352 25565 26355
rect 25572 26352 25575 26355
rect 25596 26335 25598 26355
rect 27060 26335 27062 26355
rect 27108 26335 27110 26355
rect 27180 26335 27182 26355
rect 27324 26335 27326 26355
rect 27396 26335 27398 26355
rect 27420 26335 27422 26355
rect 27540 26335 27542 26355
rect 27564 26335 27566 26355
rect 30564 26335 30566 26355
rect 30636 26335 30638 26355
rect 30660 26335 30662 26355
rect 30780 26335 30782 26355
rect 30804 26335 30806 26355
rect 30924 26335 30926 26355
rect 30948 26335 30950 26355
rect 31068 26335 31070 26355
rect 31092 26335 31094 26355
rect 31153 26350 31156 26355
rect 31164 26350 31166 26355
rect 31225 26350 31228 26355
rect 31236 26352 31238 26355
rect 31236 26350 31239 26352
rect 31163 26336 31166 26350
rect 31235 26342 31239 26350
rect 31249 26342 31253 26350
rect 31235 26336 31249 26342
rect 31105 26335 31139 26336
rect -18201 26331 -18150 26335
rect -18129 26331 -17635 26335
rect -18201 26328 -18187 26331
rect -18129 26328 -18115 26331
rect -18108 26328 -18105 26331
rect -18150 26311 -18133 26312
rect -17940 26311 -17938 26331
rect -17855 26326 -17852 26331
rect -17724 26328 -17722 26331
rect -17649 26328 -17635 26331
rect -17628 26331 -16747 26335
rect -17628 26328 -17611 26331
rect -17604 26328 -17601 26331
rect -17845 26312 -17842 26326
rect -17844 26311 -17842 26312
rect -17724 26311 -17721 26328
rect -17628 26311 -17626 26328
rect -17532 26311 -17530 26331
rect -17460 26311 -17458 26331
rect -17436 26311 -17434 26331
rect -17292 26311 -17290 26331
rect -17196 26311 -17194 26331
rect -17028 26311 -17026 26331
rect -16943 26311 -16885 26312
rect -16860 26311 -16858 26331
rect -16764 26311 -16762 26331
rect -16761 26328 -16747 26331
rect -16740 26331 -11419 26335
rect -16740 26328 -16723 26331
rect -16716 26328 -16713 26331
rect -16740 26311 -16738 26328
rect -16668 26311 -16666 26331
rect -16500 26311 -16498 26331
rect -16380 26311 -16378 26331
rect -16356 26311 -16354 26331
rect -16260 26311 -16258 26331
rect -16236 26311 -16234 26331
rect -16212 26311 -16210 26331
rect -15300 26311 -15298 26331
rect -15084 26311 -15082 26331
rect -15036 26311 -15034 26331
rect -14868 26311 -14866 26331
rect -14772 26311 -14770 26331
rect -14724 26311 -14722 26331
rect -14508 26311 -14506 26331
rect -14436 26311 -14434 26331
rect -14388 26311 -14386 26331
rect -14172 26311 -14170 26331
rect -14076 26311 -14074 26331
rect -14049 26328 -14035 26331
rect -14028 26328 -14025 26331
rect -13980 26311 -13978 26331
rect -13932 26311 -13930 26331
rect -13895 26326 -13892 26331
rect -13764 26328 -13762 26331
rect -13885 26312 -13882 26326
rect -13884 26311 -13882 26312
rect -13764 26311 -13761 26328
rect -13716 26311 -13714 26331
rect -13644 26311 -13642 26331
rect -13596 26311 -13594 26331
rect -13500 26311 -13498 26331
rect -13404 26311 -13402 26331
rect -13356 26311 -13354 26331
rect -13284 26311 -13282 26331
rect -13127 26311 -13093 26312
rect -13068 26311 -13066 26331
rect -12828 26311 -12826 26331
rect -12780 26311 -12778 26331
rect -12660 26311 -12658 26331
rect -12564 26311 -12562 26331
rect -12492 26311 -12490 26331
rect -12396 26311 -12394 26331
rect -12348 26311 -12346 26331
rect -12276 26311 -12274 26331
rect -12252 26311 -12250 26331
rect -12156 26311 -12154 26331
rect -12060 26311 -12058 26331
rect -11892 26311 -11890 26331
rect -11844 26311 -11842 26331
rect -11796 26311 -11794 26331
rect -11676 26311 -11674 26331
rect -11580 26311 -11578 26331
rect -11556 26311 -11554 26331
rect -11508 26311 -11506 26331
rect -11460 26311 -11458 26331
rect -11436 26311 -11434 26331
rect -11433 26328 -11419 26331
rect -11409 26331 12269 26335
rect -11409 26328 -11395 26331
rect -11388 26328 -11385 26331
rect -11364 26311 -11362 26331
rect -11340 26311 -11338 26331
rect -11268 26311 -11266 26331
rect -11172 26311 -11170 26331
rect -11124 26311 -11122 26331
rect -11076 26311 -11074 26331
rect -11028 26311 -11026 26331
rect -10788 26311 -10786 26331
rect -10668 26311 -10666 26331
rect -9876 26311 -9874 26331
rect -9828 26312 -9826 26331
rect -9839 26311 -9805 26312
rect -9732 26311 -9730 26331
rect -9708 26311 -9706 26331
rect -9612 26311 -9610 26331
rect -9516 26311 -9514 26331
rect -9468 26311 -9466 26331
rect -9420 26311 -9418 26331
rect -9396 26311 -9394 26331
rect -9372 26311 -9370 26331
rect -9300 26311 -9298 26331
rect -9252 26311 -9250 26331
rect -9132 26311 -9130 26331
rect -9084 26311 -9082 26331
rect -9036 26311 -9034 26331
rect -8988 26311 -8986 26331
rect -8940 26311 -8938 26331
rect -8892 26311 -8890 26331
rect -8844 26311 -8842 26331
rect -8604 26311 -8602 26331
rect -8508 26311 -8506 26331
rect -8484 26311 -8482 26331
rect -8388 26311 -8386 26331
rect -8364 26311 -8362 26331
rect -8340 26311 -8338 26331
rect -8292 26311 -8290 26331
rect -8268 26311 -8266 26331
rect -8196 26311 -8194 26331
rect -8100 26311 -8098 26331
rect -8052 26311 -8050 26331
rect -7932 26311 -7930 26331
rect -7836 26312 -7834 26331
rect -7871 26311 -7813 26312
rect -7740 26311 -7738 26331
rect -7692 26311 -7690 26331
rect -7620 26311 -7618 26331
rect -7404 26311 -7402 26331
rect -7356 26311 -7354 26331
rect -7308 26311 -7306 26331
rect -7212 26311 -7210 26331
rect -7188 26311 -7186 26331
rect -7116 26311 -7114 26331
rect -7068 26311 -7066 26331
rect -6972 26311 -6970 26331
rect -6948 26311 -6946 26331
rect -6876 26311 -6874 26331
rect -6852 26311 -6850 26331
rect -6804 26311 -6802 26331
rect -6780 26311 -6778 26331
rect -6756 26311 -6754 26331
rect -6708 26311 -6706 26331
rect -6684 26311 -6682 26331
rect -6660 26311 -6658 26331
rect -6612 26311 -6610 26331
rect -6588 26311 -6586 26331
rect -6564 26311 -6562 26331
rect -6516 26311 -6514 26331
rect -6492 26311 -6490 26331
rect -6468 26311 -6466 26331
rect -6420 26311 -6418 26331
rect -6396 26311 -6394 26331
rect -6372 26311 -6370 26331
rect -6324 26311 -6322 26331
rect -6300 26311 -6298 26331
rect -6276 26311 -6274 26331
rect -6228 26311 -6226 26331
rect -6180 26311 -6178 26331
rect -6060 26311 -6058 26331
rect -5975 26326 -5972 26331
rect -5964 26326 -5962 26331
rect -5965 26312 -5962 26326
rect -5940 26311 -5938 26331
rect -5868 26328 -5866 26331
rect -5892 26311 -5889 26328
rect -5868 26311 -5865 26328
rect -5652 26311 -5650 26331
rect -5316 26311 -5314 26331
rect -5268 26311 -5266 26331
rect -5196 26311 -5194 26331
rect -5172 26311 -5170 26331
rect -5100 26311 -5098 26331
rect -5076 26311 -5074 26331
rect -4980 26311 -4978 26331
rect -4956 26311 -4954 26331
rect -4884 26311 -4882 26331
rect -4860 26311 -4858 26331
rect -4788 26311 -4786 26331
rect -4692 26311 -4690 26331
rect -4644 26311 -4642 26331
rect -4596 26311 -4594 26331
rect -4548 26311 -4546 26331
rect -4428 26311 -4426 26331
rect -4332 26311 -4330 26331
rect -4308 26311 -4306 26331
rect -4260 26311 -4258 26331
rect -4212 26311 -4210 26331
rect -4116 26311 -4114 26331
rect -4092 26311 -4090 26331
rect -4020 26311 -4018 26331
rect -3876 26311 -3874 26331
rect -3732 26311 -3730 26331
rect -3588 26311 -3586 26331
rect -3564 26311 -3562 26331
rect -3516 26311 -3514 26331
rect -3492 26311 -3490 26331
rect -3468 26311 -3466 26331
rect -3420 26311 -3418 26331
rect -3324 26311 -3322 26331
rect -3252 26311 -3250 26331
rect -3228 26311 -3226 26331
rect -3156 26311 -3154 26331
rect -3132 26311 -3130 26331
rect -3060 26311 -3058 26331
rect -3012 26311 -3010 26331
rect -2964 26311 -2962 26331
rect -2916 26311 -2914 26331
rect -2892 26311 -2890 26331
rect -2820 26311 -2818 26331
rect -2796 26311 -2794 26331
rect -2748 26311 -2746 26331
rect -2700 26311 -2698 26331
rect -2604 26311 -2602 26331
rect -2580 26311 -2578 26331
rect -2364 26311 -2362 26331
rect -2292 26311 -2290 26331
rect -2268 26311 -2266 26331
rect -2244 26311 -2242 26331
rect -2172 26311 -2170 26331
rect -2148 26311 -2146 26331
rect -2076 26311 -2074 26331
rect -2052 26311 -2050 26331
rect -1980 26311 -1978 26331
rect -1884 26311 -1882 26331
rect -1836 26311 -1834 26331
rect -1716 26311 -1714 26331
rect -1596 26311 -1594 26331
rect -1572 26311 -1569 26328
rect -1476 26311 -1474 26331
rect -1380 26311 -1378 26331
rect -1356 26311 -1354 26331
rect -1308 26311 -1306 26331
rect -1260 26311 -1258 26331
rect -1140 26311 -1138 26331
rect -852 26311 -850 26331
rect -804 26311 -802 26331
rect -756 26311 -754 26331
rect -708 26311 -706 26331
rect -612 26311 -610 26331
rect -588 26311 -586 26331
rect -540 26311 -538 26331
rect -516 26311 -514 26331
rect -492 26311 -490 26331
rect -444 26311 -442 26331
rect -396 26311 -394 26331
rect -300 26311 -298 26331
rect -276 26311 -274 26331
rect -204 26311 -202 26331
rect -108 26311 -106 26331
rect 12 26311 14 26331
rect 108 26311 110 26331
rect 156 26311 158 26331
rect 204 26311 206 26331
rect 228 26311 230 26331
rect 252 26311 254 26331
rect 348 26311 350 26331
rect 468 26311 470 26331
rect 492 26311 494 26331
rect 564 26311 566 26331
rect 588 26311 590 26331
rect 636 26311 638 26331
rect 660 26311 662 26331
rect 673 26326 676 26331
rect 684 26326 686 26331
rect 683 26312 686 26326
rect 732 26311 734 26331
rect 756 26311 758 26331
rect 780 26328 782 26331
rect 780 26311 783 26328
rect 876 26311 878 26331
rect 972 26311 974 26331
rect 1020 26311 1022 26331
rect 1068 26311 1070 26331
rect 1092 26311 1094 26331
rect 1116 26311 1118 26331
rect 1164 26311 1166 26331
rect 1212 26311 1214 26331
rect 1308 26311 1310 26331
rect 1332 26311 1334 26331
rect 1380 26311 1382 26331
rect 1428 26311 1430 26331
rect 1524 26311 1526 26331
rect 1548 26311 1550 26331
rect 1596 26311 1598 26331
rect 1620 26311 1622 26331
rect 1644 26311 1646 26331
rect 1692 26311 1694 26331
rect 1716 26311 1718 26331
rect 1740 26311 1742 26331
rect 1788 26311 1790 26331
rect 1825 26326 1828 26331
rect 1836 26326 1838 26331
rect 1835 26312 1838 26326
rect 1884 26311 1886 26331
rect 1932 26328 1934 26331
rect 1932 26311 1935 26328
rect 1980 26311 1982 26331
rect 2028 26311 2030 26331
rect 2076 26311 2078 26331
rect 2100 26311 2102 26331
rect 2124 26311 2126 26331
rect 2172 26311 2174 26331
rect 2196 26311 2198 26331
rect 2220 26311 2222 26331
rect 2268 26311 2270 26331
rect 2292 26311 2294 26331
rect 2316 26311 2318 26331
rect 2364 26311 2366 26331
rect 2412 26311 2414 26331
rect 2460 26311 2462 26331
rect 2508 26311 2510 26331
rect 2556 26311 2558 26331
rect 2580 26311 2582 26331
rect 2604 26311 2606 26331
rect 2652 26311 2654 26331
rect 2676 26311 2678 26331
rect 2700 26311 2702 26331
rect 2748 26311 2750 26331
rect 2772 26311 2774 26331
rect 2796 26311 2798 26331
rect 2844 26311 2846 26331
rect 2868 26311 2870 26331
rect 2892 26311 2894 26331
rect 2940 26311 2942 26331
rect 3012 26311 3014 26331
rect 3108 26311 3110 26331
rect 3156 26311 3158 26331
rect 3252 26311 3254 26331
rect 3348 26311 3350 26331
rect 3396 26311 3398 26331
rect 3468 26311 3470 26331
rect 3492 26311 3494 26331
rect 3588 26311 3590 26331
rect 3612 26311 3614 26331
rect 3636 26311 3638 26331
rect 3708 26311 3710 26331
rect 3732 26311 3734 26331
rect 3804 26311 3806 26331
rect 3828 26311 3830 26331
rect 3924 26311 3926 26331
rect 4020 26311 4022 26331
rect 4044 26311 4046 26331
rect 4092 26311 4094 26331
rect 4116 26311 4118 26331
rect 4140 26311 4142 26331
rect 4188 26311 4190 26331
rect 4212 26311 4214 26331
rect 4236 26311 4238 26331
rect 4308 26311 4310 26331
rect 4332 26311 4334 26331
rect 4404 26311 4406 26331
rect 4500 26311 4502 26331
rect 4596 26311 4598 26331
rect 4860 26311 4862 26331
rect 4956 26311 4958 26331
rect 4980 26311 4982 26331
rect 5004 26311 5006 26331
rect 5076 26311 5078 26331
rect 5100 26311 5102 26331
rect 5124 26311 5126 26331
rect 5172 26311 5174 26331
rect 5196 26311 5198 26331
rect 5220 26311 5222 26331
rect 5268 26311 5270 26331
rect 5292 26311 5294 26331
rect 5388 26311 5390 26331
rect 5484 26311 5486 26331
rect 5508 26311 5510 26331
rect 5532 26311 5534 26331
rect 5569 26326 5572 26331
rect 5580 26326 5582 26331
rect 5579 26312 5582 26326
rect 5628 26311 5630 26331
rect 5652 26311 5655 26328
rect 5748 26311 5750 26331
rect 5796 26311 5798 26331
rect 5844 26311 5846 26331
rect 5892 26311 5894 26331
rect 6132 26311 6134 26331
rect 6180 26311 6182 26331
rect 6228 26311 6230 26331
rect 6252 26311 6254 26331
rect 6276 26311 6278 26331
rect 6324 26311 6326 26331
rect 6372 26311 6374 26331
rect 6492 26311 6494 26331
rect 6588 26311 6590 26331
rect 6612 26311 6614 26331
rect 6660 26311 6662 26331
rect 6684 26311 6686 26331
rect 6708 26311 6710 26331
rect 6780 26311 6782 26331
rect 6804 26311 6806 26331
rect 6828 26311 6830 26331
rect 6900 26311 6902 26331
rect 6924 26311 6926 26331
rect 7020 26311 7022 26331
rect 7140 26311 7142 26331
rect 7236 26311 7238 26331
rect 7332 26311 7334 26331
rect 7380 26311 7382 26331
rect 7428 26311 7430 26331
rect 7452 26311 7454 26331
rect 7476 26311 7478 26331
rect 7524 26311 7526 26331
rect 7548 26311 7550 26331
rect 7572 26311 7574 26331
rect 7620 26311 7622 26331
rect 7644 26311 7646 26331
rect 7668 26311 7670 26331
rect 7716 26311 7718 26331
rect 7740 26311 7742 26331
rect 7836 26311 7838 26331
rect 7884 26311 7886 26331
rect 7932 26311 7934 26331
rect 7956 26311 7958 26331
rect 7980 26311 7982 26331
rect 8017 26326 8020 26331
rect 8041 26326 8044 26331
rect 8052 26326 8054 26331
rect 8027 26312 8030 26326
rect 8051 26312 8054 26326
rect 8148 26328 8150 26331
rect 8028 26311 8030 26312
rect 8148 26311 8151 26328
rect 8196 26311 8198 26331
rect 8244 26311 8246 26331
rect 8268 26311 8270 26331
rect 8292 26311 8294 26331
rect 8340 26311 8342 26331
rect 8364 26311 8366 26331
rect 8388 26311 8390 26331
rect 8436 26311 8438 26331
rect 8460 26311 8462 26331
rect 8556 26311 8558 26331
rect 8604 26311 8606 26331
rect 8652 26311 8654 26331
rect 8700 26311 8702 26331
rect 8724 26311 8726 26331
rect 8748 26311 8750 26331
rect 8820 26311 8822 26331
rect 8844 26311 8846 26331
rect 8868 26311 8870 26331
rect 9516 26311 9518 26331
rect 9612 26311 9614 26331
rect 9660 26311 9662 26331
rect 9684 26311 9686 26331
rect 9708 26311 9710 26331
rect 9756 26311 9758 26331
rect 9780 26311 9782 26331
rect 9804 26311 9806 26331
rect 9852 26311 9854 26331
rect 9876 26311 9878 26331
rect 9900 26311 9902 26331
rect 9948 26311 9950 26331
rect 9972 26311 9974 26331
rect 9996 26311 9998 26331
rect 10068 26311 10070 26331
rect 10092 26311 10094 26331
rect 10116 26311 10118 26331
rect 10164 26311 10166 26331
rect 10188 26311 10190 26331
rect 10212 26311 10214 26331
rect 10260 26312 10262 26331
rect 10225 26311 10283 26312
rect 10284 26311 10286 26331
rect 10308 26311 10310 26331
rect 10380 26311 10382 26331
rect 10404 26311 10406 26331
rect 10428 26311 10430 26331
rect 10476 26311 10478 26331
rect 10500 26311 10502 26331
rect 10524 26311 10526 26331
rect 10572 26311 10574 26331
rect 10596 26311 10598 26331
rect 10620 26311 10622 26331
rect 10668 26311 10670 26331
rect 10692 26311 10694 26331
rect 10716 26311 10718 26331
rect 10788 26311 10790 26331
rect 10836 26311 10838 26331
rect 10956 26311 10958 26331
rect 11052 26311 11054 26331
rect 11076 26311 11078 26331
rect 11124 26311 11126 26331
rect 11172 26311 11174 26331
rect 11220 26311 11222 26331
rect 11340 26311 11342 26331
rect 11436 26311 11438 26331
rect 11532 26311 11534 26331
rect 11580 26311 11582 26331
rect 11628 26311 11630 26331
rect 11676 26311 11678 26331
rect 11772 26311 11774 26331
rect 11796 26311 11798 26331
rect 11844 26311 11846 26331
rect 11892 26311 11894 26331
rect 11988 26311 11990 26331
rect 12060 26311 12062 26331
rect 12132 26311 12134 26331
rect 12228 26311 12230 26331
rect 12255 26328 12269 26331
rect 12276 26331 31139 26335
rect 12276 26328 12293 26331
rect 12276 26311 12278 26328
rect 12324 26311 12326 26331
rect 12420 26311 12422 26331
rect 12444 26311 12446 26331
rect 12492 26311 12494 26331
rect 12516 26311 12518 26331
rect 12540 26311 12542 26331
rect 12588 26311 12590 26331
rect 12636 26311 12638 26331
rect 12732 26311 12734 26331
rect 12756 26311 12758 26331
rect 12804 26311 12806 26331
rect 12828 26311 12830 26331
rect 12852 26311 12854 26331
rect 12900 26311 12902 26331
rect 12948 26311 12950 26331
rect 13044 26311 13046 26331
rect 13068 26311 13070 26331
rect 13116 26311 13118 26331
rect 13284 26311 13286 26331
rect 13332 26311 13334 26331
rect 13428 26311 13430 26331
rect 13524 26311 13526 26331
rect 13572 26311 13574 26331
rect 13644 26311 13646 26331
rect 13668 26311 13670 26331
rect 13764 26311 13766 26331
rect 13812 26311 13814 26331
rect 13860 26311 13862 26331
rect 13908 26311 13910 26331
rect 13956 26311 13958 26331
rect 14004 26311 14006 26331
rect 14100 26311 14102 26331
rect 14196 26311 14198 26331
rect 14244 26311 14246 26331
rect 14292 26311 14294 26331
rect 15132 26311 15134 26331
rect 15169 26326 15172 26331
rect 15179 26312 15182 26326
rect 15180 26311 15182 26312
rect 15228 26311 15230 26331
rect 15252 26311 15254 26331
rect 15300 26328 15302 26331
rect 15300 26311 15303 26328
rect 15324 26311 15326 26331
rect 15396 26311 15398 26331
rect 15420 26311 15422 26331
rect 15492 26311 15494 26331
rect 15540 26311 15542 26331
rect 15636 26311 15638 26331
rect 15660 26311 15662 26331
rect 15708 26311 15710 26331
rect 15732 26311 15734 26331
rect 15756 26311 15758 26331
rect 15804 26311 15806 26331
rect 15828 26311 15830 26331
rect 15852 26311 15854 26331
rect 15900 26311 15902 26331
rect 15948 26311 15950 26331
rect 15996 26311 15998 26331
rect 16044 26311 16046 26331
rect 16092 26311 16094 26331
rect 16140 26311 16142 26331
rect 16236 26311 16238 26331
rect 16260 26311 16262 26331
rect 16308 26311 16310 26331
rect 16332 26311 16334 26331
rect 16356 26311 16358 26331
rect 16404 26311 16406 26331
rect 16452 26311 16454 26331
rect 16548 26311 16550 26331
rect 16572 26311 16574 26331
rect 16620 26311 16622 26331
rect 16668 26311 16670 26331
rect 16716 26311 16718 26331
rect 16764 26311 16766 26331
rect 16836 26311 16838 26331
rect 16884 26311 16886 26331
rect 16980 26311 16982 26331
rect 17052 26311 17054 26331
rect 17196 26311 17198 26331
rect 17220 26311 17222 26331
rect 17292 26311 17294 26331
rect 17316 26311 17318 26331
rect 18084 26311 18086 26331
rect 18132 26311 18134 26331
rect 18396 26311 18398 26331
rect 18492 26311 18494 26331
rect 18516 26311 18518 26331
rect 18564 26311 18566 26331
rect 18612 26311 18614 26331
rect 18660 26311 18662 26331
rect 18708 26311 18710 26331
rect 18756 26311 18758 26331
rect 18804 26311 18806 26331
rect 18852 26311 18854 26331
rect 18900 26311 18902 26331
rect 18996 26311 18998 26331
rect 19020 26311 19022 26331
rect 19092 26311 19094 26331
rect 19116 26311 19118 26331
rect 19140 26311 19142 26331
rect 19188 26311 19190 26331
rect 19236 26311 19238 26331
rect 19332 26311 19334 26331
rect 19476 26311 19478 26331
rect 19620 26311 19622 26331
rect 19716 26311 19718 26331
rect 19788 26311 19790 26331
rect 19836 26311 19838 26331
rect 19860 26311 19862 26331
rect 19884 26311 19886 26331
rect 19932 26311 19934 26331
rect 19956 26311 19958 26331
rect 19980 26311 19982 26331
rect 20028 26311 20030 26331
rect 20052 26311 20054 26331
rect 20076 26311 20078 26331
rect 20148 26311 20150 26331
rect 20172 26311 20174 26331
rect 20196 26311 20198 26331
rect 20268 26311 20270 26331
rect 20292 26311 20294 26331
rect 20388 26311 20390 26331
rect 20412 26311 20414 26331
rect 20508 26311 20510 26331
rect 20556 26311 20558 26331
rect 20604 26311 20606 26331
rect 20916 26311 20918 26331
rect 20964 26311 20966 26331
rect 21012 26311 21014 26331
rect 21060 26311 21062 26331
rect 21084 26311 21086 26331
rect 21108 26311 21110 26331
rect 21204 26311 21206 26331
rect 21300 26311 21302 26331
rect 21324 26311 21326 26331
rect 21444 26311 21446 26331
rect 21468 26311 21470 26331
rect 21564 26311 21566 26331
rect 21612 26311 21614 26331
rect 21684 26311 21686 26331
rect 21708 26311 21710 26331
rect 21804 26311 21806 26331
rect 21828 26311 21830 26331
rect 21924 26311 21926 26331
rect 21948 26311 21950 26331
rect 22044 26311 22046 26331
rect 22068 26311 22070 26331
rect 22188 26311 22190 26331
rect 22212 26311 22214 26331
rect 23004 26311 23006 26331
rect 23052 26311 23054 26331
rect 23076 26311 23078 26331
rect 23100 26311 23102 26331
rect 23148 26311 23150 26331
rect 23220 26311 23222 26331
rect 23244 26311 23246 26331
rect 23316 26311 23318 26331
rect 23340 26311 23342 26331
rect 23412 26311 23414 26331
rect 23556 26311 23558 26331
rect 23628 26311 23630 26331
rect 23652 26311 23654 26331
rect 23676 26311 23678 26331
rect 23724 26311 23726 26331
rect 23772 26311 23774 26331
rect 23820 26311 23822 26331
rect 23868 26311 23870 26331
rect 23916 26311 23918 26331
rect 24012 26311 24014 26331
rect 24084 26311 24086 26331
rect 24372 26311 24374 26331
rect 24396 26311 24398 26331
rect 24492 26311 24494 26331
rect 24516 26311 24518 26331
rect 24588 26311 24590 26331
rect 24612 26311 24614 26331
rect 24708 26311 24710 26331
rect 24732 26311 24734 26331
rect 24756 26311 24758 26331
rect 24852 26311 24854 26331
rect 24876 26311 24878 26331
rect 24972 26311 24974 26331
rect 24996 26311 24998 26331
rect 25092 26311 25094 26331
rect 25260 26311 25262 26331
rect 25297 26311 25355 26312
rect 25356 26311 25358 26331
rect 25380 26311 25382 26331
rect 25452 26311 25454 26331
rect 25500 26311 25502 26331
rect 25596 26311 25598 26331
rect 27060 26311 27062 26331
rect 27108 26311 27110 26331
rect 27180 26312 27182 26331
rect 27145 26311 27203 26312
rect 27324 26311 27326 26331
rect 27396 26311 27398 26331
rect 27420 26311 27422 26331
rect 27540 26311 27542 26331
rect 27564 26311 27566 26331
rect 30564 26311 30566 26331
rect 30636 26311 30638 26331
rect 30660 26311 30662 26331
rect 30780 26311 30782 26331
rect 30804 26311 30806 26331
rect 30924 26311 30926 26331
rect 30948 26311 30950 26331
rect 31068 26311 31070 26331
rect 31092 26312 31094 26331
rect 31081 26311 31115 26312
rect -18150 26307 -17755 26311
rect -17940 26287 -17938 26307
rect -17844 26287 -17842 26307
rect -17769 26304 -17755 26307
rect -17745 26307 -13795 26311
rect -17745 26304 -17731 26307
rect -17724 26304 -17721 26307
rect -17628 26288 -17626 26307
rect -17783 26287 -17749 26288
rect -17639 26287 -17605 26288
rect -17532 26287 -17530 26307
rect -17495 26287 -17461 26288
rect -18081 26283 -17461 26287
rect -18081 26280 -18067 26283
rect -18033 26263 -18013 26264
rect -17940 26263 -17938 26283
rect -17844 26263 -17842 26283
rect -17639 26278 -17636 26283
rect -17628 26278 -17626 26283
rect -17629 26264 -17626 26278
rect -17532 26280 -17530 26283
rect -17532 26264 -17529 26280
rect -17591 26263 -17557 26264
rect -18033 26259 -17557 26263
rect -17543 26263 -17509 26264
rect -17460 26263 -17458 26307
rect -17436 26263 -17434 26307
rect -17423 26287 -17389 26288
rect -17292 26287 -17290 26307
rect -17196 26287 -17194 26307
rect -17028 26287 -17026 26307
rect -16943 26302 -16940 26307
rect -16933 26288 -16930 26302
rect -16932 26287 -16930 26288
rect -16860 26287 -16858 26307
rect -16836 26287 -16833 26304
rect -16764 26287 -16762 26307
rect -16740 26287 -16738 26307
rect -16668 26287 -16666 26307
rect -16500 26287 -16498 26307
rect -16380 26287 -16378 26307
rect -16356 26287 -16354 26307
rect -16295 26287 -16261 26288
rect -17423 26283 -16843 26287
rect -17399 26270 -17395 26278
rect -17409 26264 -17399 26270
rect -17543 26259 -17395 26263
rect -18033 26256 -18019 26259
rect -17940 26256 -17938 26259
rect -17940 26239 -17937 26256
rect -17844 26239 -17842 26259
rect -17697 26256 -17683 26259
rect -17543 26256 -17539 26259
rect -17532 26256 -17529 26259
rect -17519 26239 -17491 26240
rect -17961 26235 -17491 26239
rect -17961 26232 -17947 26235
rect -17940 26232 -17937 26235
rect -17844 26215 -17842 26235
rect -17519 26230 -17516 26235
rect -17505 26232 -17491 26235
rect -17484 26232 -17481 26256
rect -17509 26216 -17506 26230
rect -17508 26215 -17506 26216
rect -17484 26215 -17482 26232
rect -17471 26230 -17468 26240
rect -17460 26230 -17458 26259
rect -17436 26256 -17434 26259
rect -17409 26256 -17395 26259
rect -17388 26256 -17385 26280
rect -17292 26263 -17290 26283
rect -17196 26263 -17194 26283
rect -17028 26263 -17026 26283
rect -16932 26263 -16930 26283
rect -16860 26263 -16858 26283
rect -16857 26280 -16843 26283
rect -16836 26283 -16261 26287
rect -16836 26280 -16819 26283
rect -16836 26263 -16834 26280
rect -16764 26263 -16762 26283
rect -16740 26263 -16738 26283
rect -16668 26263 -16666 26283
rect -16500 26263 -16498 26283
rect -16380 26263 -16378 26283
rect -16356 26263 -16354 26283
rect -16295 26278 -16292 26283
rect -16285 26264 -16282 26278
rect -16284 26263 -16282 26264
rect -16260 26263 -16258 26307
rect -16236 26263 -16234 26307
rect -16212 26288 -16210 26307
rect -16223 26287 -16189 26288
rect -15300 26287 -15298 26307
rect -15084 26287 -15082 26307
rect -15036 26287 -15034 26307
rect -14868 26287 -14866 26307
rect -14772 26287 -14770 26307
rect -14724 26287 -14722 26307
rect -14508 26287 -14506 26307
rect -14436 26287 -14434 26307
rect -14388 26287 -14386 26307
rect -14172 26287 -14170 26307
rect -14076 26287 -14074 26307
rect -13980 26287 -13978 26307
rect -13932 26287 -13930 26307
rect -13884 26287 -13882 26307
rect -13809 26304 -13795 26307
rect -13785 26307 -5899 26311
rect -13785 26304 -13771 26307
rect -13764 26304 -13761 26307
rect -13716 26287 -13714 26307
rect -13644 26287 -13642 26307
rect -13596 26287 -13594 26307
rect -13500 26287 -13498 26307
rect -13404 26287 -13402 26307
rect -13356 26287 -13354 26307
rect -13284 26287 -13282 26307
rect -13068 26287 -13066 26307
rect -12828 26287 -12826 26307
rect -12780 26287 -12778 26307
rect -12660 26287 -12658 26307
rect -12564 26287 -12562 26307
rect -12492 26287 -12490 26307
rect -12396 26287 -12394 26307
rect -12348 26287 -12346 26307
rect -12276 26287 -12274 26307
rect -12252 26287 -12250 26307
rect -12156 26287 -12154 26307
rect -12060 26287 -12058 26307
rect -11892 26287 -11890 26307
rect -11844 26287 -11842 26307
rect -11796 26287 -11794 26307
rect -11676 26287 -11674 26307
rect -11580 26287 -11578 26307
rect -11556 26287 -11554 26307
rect -11508 26287 -11506 26307
rect -11460 26287 -11458 26307
rect -11436 26287 -11434 26307
rect -11364 26287 -11362 26307
rect -11340 26287 -11338 26307
rect -11268 26287 -11266 26307
rect -11172 26287 -11170 26307
rect -11124 26287 -11122 26307
rect -11076 26287 -11074 26307
rect -11028 26287 -11026 26307
rect -10788 26287 -10786 26307
rect -10668 26287 -10666 26307
rect -9876 26287 -9874 26307
rect -9839 26302 -9836 26307
rect -9828 26302 -9826 26307
rect -9829 26288 -9826 26302
rect -9732 26304 -9730 26307
rect -9732 26287 -9729 26304
rect -9708 26287 -9706 26307
rect -9612 26287 -9610 26307
rect -9516 26287 -9514 26307
rect -9468 26287 -9466 26307
rect -9420 26287 -9418 26307
rect -9396 26287 -9394 26307
rect -9372 26287 -9370 26307
rect -9300 26287 -9298 26307
rect -9252 26287 -9250 26307
rect -9132 26287 -9130 26307
rect -9084 26287 -9082 26307
rect -9036 26287 -9034 26307
rect -8988 26287 -8986 26307
rect -8940 26287 -8938 26307
rect -8892 26287 -8890 26307
rect -8844 26287 -8842 26307
rect -8604 26287 -8602 26307
rect -8508 26287 -8506 26307
rect -8484 26287 -8482 26307
rect -8388 26287 -8386 26307
rect -8364 26287 -8362 26307
rect -8340 26287 -8338 26307
rect -8292 26288 -8290 26307
rect -8303 26287 -8269 26288
rect -8268 26287 -8266 26307
rect -8196 26287 -8194 26307
rect -8100 26287 -8098 26307
rect -8052 26287 -8050 26307
rect -7932 26287 -7930 26307
rect -7847 26302 -7844 26307
rect -7836 26302 -7834 26307
rect -7837 26288 -7834 26302
rect -7740 26304 -7738 26307
rect -7740 26287 -7737 26304
rect -7692 26287 -7690 26307
rect -7620 26287 -7618 26307
rect -7404 26287 -7402 26307
rect -7356 26287 -7354 26307
rect -7308 26287 -7306 26307
rect -7212 26287 -7210 26307
rect -7188 26287 -7186 26307
rect -7116 26287 -7114 26307
rect -7068 26287 -7066 26307
rect -6972 26287 -6970 26307
rect -6948 26287 -6946 26307
rect -6876 26287 -6874 26307
rect -6852 26287 -6850 26307
rect -6804 26287 -6802 26307
rect -6780 26287 -6778 26307
rect -6756 26287 -6754 26307
rect -6708 26287 -6706 26307
rect -6684 26288 -6682 26307
rect -6695 26287 -6661 26288
rect -6660 26287 -6658 26307
rect -6612 26287 -6610 26307
rect -6588 26287 -6586 26307
rect -6564 26287 -6562 26307
rect -6516 26287 -6514 26307
rect -6492 26287 -6490 26307
rect -6468 26287 -6466 26307
rect -6420 26287 -6418 26307
rect -6396 26287 -6394 26307
rect -6372 26287 -6370 26307
rect -6324 26287 -6322 26307
rect -6300 26287 -6298 26307
rect -6276 26287 -6274 26307
rect -6228 26287 -6226 26307
rect -6180 26287 -6178 26307
rect -6060 26287 -6058 26307
rect -5940 26287 -5938 26307
rect -5913 26304 -5899 26307
rect -5892 26307 -1579 26311
rect -5892 26304 -5875 26307
rect -5868 26304 -5865 26307
rect -5892 26287 -5890 26304
rect -5652 26287 -5650 26307
rect -5316 26287 -5314 26307
rect -5268 26287 -5266 26307
rect -5196 26287 -5194 26307
rect -5172 26287 -5170 26307
rect -5100 26287 -5098 26307
rect -5076 26287 -5074 26307
rect -4980 26287 -4978 26307
rect -4956 26287 -4954 26307
rect -4884 26287 -4882 26307
rect -4860 26287 -4858 26307
rect -4788 26287 -4786 26307
rect -4692 26287 -4690 26307
rect -4644 26287 -4642 26307
rect -4596 26287 -4594 26307
rect -4548 26287 -4546 26307
rect -4428 26288 -4426 26307
rect -4439 26287 -4405 26288
rect -4332 26287 -4330 26307
rect -4308 26287 -4306 26307
rect -4260 26287 -4258 26307
rect -4212 26287 -4210 26307
rect -4116 26287 -4114 26307
rect -4092 26287 -4090 26307
rect -4020 26287 -4018 26307
rect -3876 26287 -3874 26307
rect -3732 26287 -3730 26307
rect -3588 26287 -3586 26307
rect -3564 26287 -3562 26307
rect -3516 26287 -3514 26307
rect -3492 26287 -3490 26307
rect -3468 26287 -3466 26307
rect -3420 26287 -3418 26307
rect -3324 26287 -3322 26307
rect -3252 26287 -3250 26307
rect -3228 26287 -3226 26307
rect -3156 26287 -3154 26307
rect -3132 26287 -3130 26307
rect -3060 26287 -3058 26307
rect -3012 26287 -3010 26307
rect -2964 26287 -2962 26307
rect -2916 26287 -2914 26307
rect -2892 26287 -2890 26307
rect -2820 26287 -2818 26307
rect -2796 26287 -2794 26307
rect -2748 26287 -2746 26307
rect -2700 26287 -2698 26307
rect -2604 26287 -2602 26307
rect -2580 26287 -2578 26307
rect -2399 26287 -2365 26288
rect -2364 26287 -2362 26307
rect -2292 26287 -2290 26307
rect -2268 26287 -2266 26307
rect -2244 26287 -2242 26307
rect -2172 26287 -2170 26307
rect -2148 26287 -2146 26307
rect -2076 26287 -2074 26307
rect -2052 26287 -2050 26307
rect -1980 26287 -1978 26307
rect -1884 26287 -1882 26307
rect -1836 26287 -1834 26307
rect -1716 26287 -1714 26307
rect -1596 26287 -1594 26307
rect -1593 26304 -1579 26307
rect -1572 26307 5645 26311
rect -1572 26304 -1555 26307
rect -1572 26287 -1570 26304
rect -1476 26287 -1474 26307
rect -1380 26287 -1378 26307
rect -1356 26287 -1354 26307
rect -1308 26287 -1306 26307
rect -1260 26287 -1258 26307
rect -1140 26287 -1138 26307
rect -852 26287 -850 26307
rect -804 26287 -802 26307
rect -756 26287 -754 26307
rect -708 26287 -706 26307
rect -612 26287 -610 26307
rect -588 26287 -586 26307
rect -540 26287 -538 26307
rect -516 26288 -514 26307
rect -527 26287 -493 26288
rect -492 26287 -490 26307
rect -444 26287 -442 26307
rect -396 26287 -394 26307
rect -300 26287 -298 26307
rect -276 26287 -274 26307
rect -204 26287 -202 26307
rect -108 26287 -106 26307
rect 12 26287 14 26307
rect 108 26287 110 26307
rect 156 26287 158 26307
rect 204 26287 206 26307
rect 228 26287 230 26307
rect 252 26287 254 26307
rect 348 26287 350 26307
rect 468 26287 470 26307
rect 492 26287 494 26307
rect 564 26287 566 26307
rect 588 26287 590 26307
rect 636 26287 638 26307
rect 660 26287 662 26307
rect 732 26287 734 26307
rect 756 26287 758 26307
rect 759 26304 773 26307
rect 780 26304 783 26307
rect 876 26287 878 26307
rect 972 26287 974 26307
rect 1020 26287 1022 26307
rect 1068 26287 1070 26307
rect 1092 26287 1094 26307
rect 1116 26287 1118 26307
rect 1164 26287 1166 26307
rect 1212 26287 1214 26307
rect 1308 26287 1310 26307
rect 1332 26287 1334 26307
rect 1380 26287 1382 26307
rect 1428 26287 1430 26307
rect 1524 26287 1526 26307
rect 1548 26287 1550 26307
rect 1596 26287 1598 26307
rect 1620 26287 1622 26307
rect 1644 26287 1646 26307
rect 1692 26287 1694 26307
rect 1716 26287 1718 26307
rect 1740 26287 1742 26307
rect 1788 26287 1790 26307
rect 1884 26287 1886 26307
rect 1911 26304 1925 26307
rect 1932 26304 1935 26307
rect 1980 26287 1982 26307
rect 2028 26287 2030 26307
rect 2076 26287 2078 26307
rect 2100 26287 2102 26307
rect 2124 26287 2126 26307
rect 2172 26287 2174 26307
rect 2196 26287 2198 26307
rect 2220 26287 2222 26307
rect 2268 26287 2270 26307
rect 2292 26287 2294 26307
rect 2316 26287 2318 26307
rect 2364 26287 2366 26307
rect 2412 26287 2414 26307
rect 2460 26287 2462 26307
rect 2508 26287 2510 26307
rect 2556 26287 2558 26307
rect 2580 26287 2582 26307
rect 2604 26287 2606 26307
rect 2652 26287 2654 26307
rect 2676 26287 2678 26307
rect 2700 26287 2702 26307
rect 2748 26287 2750 26307
rect 2772 26287 2774 26307
rect 2796 26287 2798 26307
rect 2844 26287 2846 26307
rect 2868 26287 2870 26307
rect 2892 26287 2894 26307
rect 2940 26287 2942 26307
rect 3012 26287 3014 26307
rect 3108 26287 3110 26307
rect 3156 26287 3158 26307
rect 3252 26287 3254 26307
rect 3348 26287 3350 26307
rect 3396 26287 3398 26307
rect 3468 26287 3470 26307
rect 3492 26287 3494 26307
rect 3588 26287 3590 26307
rect 3612 26287 3614 26307
rect 3636 26287 3638 26307
rect 3708 26287 3710 26307
rect 3732 26287 3734 26307
rect 3804 26287 3806 26307
rect 3828 26287 3830 26307
rect 3924 26287 3926 26307
rect 4020 26287 4022 26307
rect 4044 26287 4046 26307
rect 4092 26287 4094 26307
rect 4116 26287 4118 26307
rect 4140 26287 4142 26307
rect 4188 26287 4190 26307
rect 4212 26287 4214 26307
rect 4236 26287 4238 26307
rect 4308 26287 4310 26307
rect 4332 26287 4334 26307
rect 4404 26287 4406 26307
rect 4500 26287 4502 26307
rect 4596 26287 4598 26307
rect 4860 26287 4862 26307
rect 4956 26287 4958 26307
rect 4980 26287 4982 26307
rect 5004 26287 5006 26307
rect 5076 26287 5078 26307
rect 5100 26287 5102 26307
rect 5124 26287 5126 26307
rect 5172 26287 5174 26307
rect 5196 26287 5198 26307
rect 5220 26287 5222 26307
rect 5268 26287 5270 26307
rect 5292 26287 5294 26307
rect 5388 26287 5390 26307
rect 5484 26287 5486 26307
rect 5508 26287 5510 26307
rect 5532 26287 5534 26307
rect 5628 26287 5630 26307
rect 5631 26304 5645 26307
rect 5652 26307 8117 26311
rect 5652 26304 5669 26307
rect 5652 26287 5654 26304
rect 5748 26287 5750 26307
rect 5796 26287 5798 26307
rect 5844 26287 5846 26307
rect 5892 26287 5894 26307
rect 6132 26287 6134 26307
rect 6180 26287 6182 26307
rect 6228 26287 6230 26307
rect 6252 26287 6254 26307
rect 6276 26287 6278 26307
rect 6324 26287 6326 26307
rect 6372 26287 6374 26307
rect 6492 26287 6494 26307
rect 6588 26287 6590 26307
rect 6612 26287 6614 26307
rect 6660 26287 6662 26307
rect 6684 26287 6686 26307
rect 6708 26287 6710 26307
rect 6780 26287 6782 26307
rect 6804 26287 6806 26307
rect 6828 26287 6830 26307
rect 6900 26287 6902 26307
rect 6924 26287 6926 26307
rect 7020 26287 7022 26307
rect 7140 26287 7142 26307
rect 7236 26287 7238 26307
rect 7332 26287 7334 26307
rect 7380 26287 7382 26307
rect 7428 26287 7430 26307
rect 7452 26287 7454 26307
rect 7476 26287 7478 26307
rect 7524 26287 7526 26307
rect 7548 26287 7550 26307
rect 7572 26287 7574 26307
rect 7620 26287 7622 26307
rect 7644 26287 7646 26307
rect 7668 26287 7670 26307
rect 7716 26287 7718 26307
rect 7740 26287 7742 26307
rect 7836 26287 7838 26307
rect 7884 26287 7886 26307
rect 7932 26287 7934 26307
rect 7956 26287 7958 26307
rect 7980 26287 7982 26307
rect 8028 26287 8030 26307
rect 8103 26304 8117 26307
rect 8127 26307 15269 26311
rect 8127 26304 8141 26307
rect 8148 26304 8151 26307
rect 8196 26287 8198 26307
rect 8244 26287 8246 26307
rect 8268 26287 8270 26307
rect 8292 26287 8294 26307
rect 8340 26287 8342 26307
rect 8364 26287 8366 26307
rect 8388 26287 8390 26307
rect 8436 26287 8438 26307
rect 8460 26287 8462 26307
rect 8556 26287 8558 26307
rect 8604 26287 8606 26307
rect 8652 26287 8654 26307
rect 8700 26287 8702 26307
rect 8724 26287 8726 26307
rect 8748 26287 8750 26307
rect 8820 26287 8822 26307
rect 8844 26287 8846 26307
rect 8868 26287 8870 26307
rect 9516 26287 9518 26307
rect 9612 26287 9614 26307
rect 9660 26287 9662 26307
rect 9684 26287 9686 26307
rect 9708 26287 9710 26307
rect 9756 26287 9758 26307
rect 9780 26287 9782 26307
rect 9804 26287 9806 26307
rect 9852 26287 9854 26307
rect 9876 26287 9878 26307
rect 9900 26287 9902 26307
rect 9948 26287 9950 26307
rect 9972 26287 9974 26307
rect 9996 26287 9998 26307
rect 10068 26287 10070 26307
rect 10092 26287 10094 26307
rect 10116 26287 10118 26307
rect 10164 26287 10166 26307
rect 10188 26287 10190 26307
rect 10212 26287 10214 26307
rect 10249 26302 10252 26307
rect 10260 26302 10262 26307
rect 10259 26288 10262 26302
rect 10284 26287 10286 26307
rect 10308 26287 10310 26307
rect 10332 26287 10335 26304
rect 10380 26287 10382 26307
rect 10404 26287 10406 26307
rect 10428 26287 10430 26307
rect 10476 26287 10478 26307
rect 10500 26287 10502 26307
rect 10524 26287 10526 26307
rect 10572 26287 10574 26307
rect 10596 26287 10598 26307
rect 10620 26287 10622 26307
rect 10668 26287 10670 26307
rect 10692 26287 10694 26307
rect 10716 26287 10718 26307
rect 10788 26287 10790 26307
rect 10836 26287 10838 26307
rect 10956 26287 10958 26307
rect 11052 26287 11054 26307
rect 11076 26287 11078 26307
rect 11124 26287 11126 26307
rect 11172 26287 11174 26307
rect 11220 26287 11222 26307
rect 11340 26287 11342 26307
rect 11436 26287 11438 26307
rect 11532 26287 11534 26307
rect 11580 26287 11582 26307
rect 11628 26287 11630 26307
rect 11676 26287 11678 26307
rect 11713 26287 11771 26288
rect 11772 26287 11774 26307
rect 11796 26287 11798 26307
rect 11844 26287 11846 26307
rect 11892 26287 11894 26307
rect 11988 26287 11990 26307
rect 12060 26287 12062 26307
rect 12132 26287 12134 26307
rect 12228 26287 12230 26307
rect 12276 26287 12278 26307
rect 12324 26287 12326 26307
rect 12420 26287 12422 26307
rect 12444 26287 12446 26307
rect 12492 26287 12494 26307
rect 12516 26287 12518 26307
rect 12540 26287 12542 26307
rect 12588 26287 12590 26307
rect 12636 26287 12638 26307
rect 12732 26287 12734 26307
rect 12756 26287 12758 26307
rect 12804 26287 12806 26307
rect 12828 26287 12830 26307
rect 12852 26287 12854 26307
rect 12900 26287 12902 26307
rect 12948 26287 12950 26307
rect 13044 26287 13046 26307
rect 13068 26287 13070 26307
rect 13116 26287 13118 26307
rect 13284 26287 13286 26307
rect 13332 26287 13334 26307
rect 13428 26287 13430 26307
rect 13524 26287 13526 26307
rect 13572 26287 13574 26307
rect 13644 26287 13646 26307
rect 13668 26287 13670 26307
rect 13764 26287 13766 26307
rect 13812 26287 13814 26307
rect 13860 26287 13862 26307
rect 13908 26287 13910 26307
rect 13956 26287 13958 26307
rect 14004 26287 14006 26307
rect 14100 26287 14102 26307
rect 14137 26287 14171 26288
rect 14196 26287 14198 26307
rect 14244 26287 14246 26307
rect 14292 26287 14294 26307
rect 15132 26287 15134 26307
rect 15180 26287 15182 26307
rect 15228 26287 15230 26307
rect 15252 26287 15254 26307
rect 15255 26304 15269 26307
rect 15279 26307 31115 26311
rect 15279 26304 15293 26307
rect 15300 26304 15303 26307
rect 15324 26287 15326 26307
rect 15396 26287 15398 26307
rect 15420 26287 15422 26307
rect 15492 26287 15494 26307
rect 15540 26287 15542 26307
rect 15636 26287 15638 26307
rect 15660 26287 15662 26307
rect 15708 26287 15710 26307
rect 15732 26287 15734 26307
rect 15756 26287 15758 26307
rect 15804 26287 15806 26307
rect 15828 26287 15830 26307
rect 15852 26287 15854 26307
rect 15900 26287 15902 26307
rect 15948 26287 15950 26307
rect 15996 26287 15998 26307
rect 16044 26287 16046 26307
rect 16092 26287 16094 26307
rect 16140 26287 16142 26307
rect 16236 26287 16238 26307
rect 16260 26287 16262 26307
rect 16308 26287 16310 26307
rect 16332 26287 16334 26307
rect 16356 26287 16358 26307
rect 16404 26287 16406 26307
rect 16452 26287 16454 26307
rect 16548 26287 16550 26307
rect 16572 26287 16574 26307
rect 16620 26287 16622 26307
rect 16668 26287 16670 26307
rect 16716 26287 16718 26307
rect 16764 26287 16766 26307
rect 16836 26287 16838 26307
rect 16884 26287 16886 26307
rect 16980 26287 16982 26307
rect 17052 26287 17054 26307
rect 17196 26287 17198 26307
rect 17220 26287 17222 26307
rect 17292 26287 17294 26307
rect 17316 26287 17318 26307
rect 18084 26287 18086 26307
rect 18132 26287 18134 26307
rect 18396 26287 18398 26307
rect 18492 26287 18494 26307
rect 18516 26287 18518 26307
rect 18564 26287 18566 26307
rect 18612 26287 18614 26307
rect 18660 26287 18662 26307
rect 18708 26287 18710 26307
rect 18756 26287 18758 26307
rect 18804 26287 18806 26307
rect 18852 26287 18854 26307
rect 18900 26287 18902 26307
rect 18996 26287 18998 26307
rect 19020 26287 19022 26307
rect 19092 26287 19094 26307
rect 19116 26287 19118 26307
rect 19140 26287 19142 26307
rect 19188 26287 19190 26307
rect 19236 26287 19238 26307
rect 19332 26287 19334 26307
rect 19476 26287 19478 26307
rect 19620 26287 19622 26307
rect 19716 26287 19718 26307
rect 19788 26287 19790 26307
rect 19836 26287 19838 26307
rect 19860 26287 19862 26307
rect 19884 26287 19886 26307
rect 19932 26287 19934 26307
rect 19956 26287 19958 26307
rect 19980 26287 19982 26307
rect 20028 26287 20030 26307
rect 20052 26287 20054 26307
rect 20076 26287 20078 26307
rect 20148 26287 20150 26307
rect 20172 26287 20174 26307
rect 20196 26287 20198 26307
rect 20268 26287 20270 26307
rect 20292 26287 20294 26307
rect 20388 26287 20390 26307
rect 20412 26287 20414 26307
rect 20508 26287 20510 26307
rect 20556 26287 20558 26307
rect 20604 26287 20606 26307
rect 20916 26287 20918 26307
rect 20964 26287 20966 26307
rect 21012 26287 21014 26307
rect 21060 26287 21062 26307
rect 21084 26287 21086 26307
rect 21108 26287 21110 26307
rect 21204 26287 21206 26307
rect 21300 26287 21302 26307
rect 21324 26287 21326 26307
rect 21444 26287 21446 26307
rect 21468 26287 21470 26307
rect 21564 26287 21566 26307
rect 21612 26287 21614 26307
rect 21684 26287 21686 26307
rect 21708 26287 21710 26307
rect 21804 26288 21806 26307
rect 21793 26287 21827 26288
rect 21828 26287 21830 26307
rect 21924 26287 21926 26307
rect 21948 26287 21950 26307
rect 22044 26287 22046 26307
rect 22068 26287 22070 26307
rect 22188 26287 22190 26307
rect 22212 26287 22214 26307
rect 23004 26287 23006 26307
rect 23052 26287 23054 26307
rect 23076 26287 23078 26307
rect 23100 26287 23102 26307
rect 23148 26287 23150 26307
rect 23220 26287 23222 26307
rect 23244 26287 23246 26307
rect 23316 26287 23318 26307
rect 23340 26287 23342 26307
rect 23412 26287 23414 26307
rect 23556 26287 23558 26307
rect 23628 26287 23630 26307
rect 23652 26287 23654 26307
rect 23676 26287 23678 26307
rect 23724 26287 23726 26307
rect 23772 26287 23774 26307
rect 23820 26287 23822 26307
rect 23868 26287 23870 26307
rect 23916 26287 23918 26307
rect 24012 26287 24014 26307
rect 24084 26287 24086 26307
rect 24372 26287 24374 26307
rect 24396 26287 24398 26307
rect 24492 26287 24494 26307
rect 24516 26287 24518 26307
rect 24588 26287 24590 26307
rect 24612 26287 24614 26307
rect 24708 26287 24710 26307
rect 24732 26287 24734 26307
rect 24756 26287 24758 26307
rect 24852 26287 24854 26307
rect 24876 26287 24878 26307
rect 24972 26287 24974 26307
rect 24996 26287 24998 26307
rect 25033 26287 25067 26288
rect 25092 26287 25094 26307
rect 25260 26287 25262 26307
rect 25297 26302 25300 26307
rect 25307 26288 25310 26302
rect 25308 26287 25310 26288
rect 25356 26287 25358 26307
rect 25380 26287 25382 26307
rect 25404 26287 25407 26304
rect 25452 26287 25454 26307
rect 25500 26287 25502 26307
rect 25596 26287 25598 26307
rect 27060 26287 27062 26307
rect 27108 26287 27110 26307
rect 27145 26302 27148 26307
rect 27169 26302 27172 26307
rect 27180 26302 27182 26307
rect 27155 26288 27158 26302
rect 27179 26288 27182 26302
rect 27156 26287 27158 26288
rect 27324 26287 27326 26307
rect 27396 26287 27398 26307
rect 27420 26287 27422 26307
rect 27540 26287 27542 26307
rect 27564 26287 27566 26307
rect 30564 26287 30566 26307
rect 30636 26287 30638 26307
rect 30660 26287 30662 26307
rect 30780 26287 30782 26307
rect 30804 26287 30806 26307
rect 30817 26287 30851 26288
rect 30924 26287 30926 26307
rect 30948 26287 30950 26307
rect 31068 26288 31070 26307
rect 31081 26302 31084 26307
rect 31092 26302 31094 26307
rect 31091 26288 31094 26302
rect 31057 26287 31091 26288
rect -16223 26283 -7771 26287
rect -16223 26278 -16220 26283
rect -16212 26278 -16210 26283
rect -16213 26264 -16210 26278
rect -16199 26270 -16195 26278
rect -16209 26264 -16199 26270
rect -15300 26263 -15298 26283
rect -15084 26263 -15082 26283
rect -15036 26263 -15034 26283
rect -14868 26263 -14866 26283
rect -14772 26263 -14770 26283
rect -14724 26263 -14722 26283
rect -14508 26263 -14506 26283
rect -14436 26263 -14434 26283
rect -14388 26264 -14386 26283
rect -14399 26263 -14365 26264
rect -14351 26263 -14293 26264
rect -14172 26263 -14170 26283
rect -14076 26263 -14074 26283
rect -13980 26263 -13978 26283
rect -13932 26263 -13930 26283
rect -13884 26263 -13882 26283
rect -13716 26263 -13714 26283
rect -13644 26263 -13642 26283
rect -13596 26263 -13594 26283
rect -13500 26263 -13498 26283
rect -13404 26263 -13402 26283
rect -13356 26263 -13354 26283
rect -13284 26263 -13282 26283
rect -13068 26263 -13066 26283
rect -13041 26280 -13027 26283
rect -12828 26263 -12826 26283
rect -12780 26263 -12778 26283
rect -12660 26263 -12658 26283
rect -12564 26263 -12562 26283
rect -12492 26263 -12490 26283
rect -12396 26263 -12394 26283
rect -12348 26263 -12346 26283
rect -12276 26263 -12274 26283
rect -12252 26263 -12250 26283
rect -12156 26263 -12154 26283
rect -12060 26263 -12058 26283
rect -11892 26263 -11890 26283
rect -11844 26263 -11842 26283
rect -11796 26263 -11794 26283
rect -11676 26263 -11674 26283
rect -11580 26263 -11578 26283
rect -11556 26263 -11554 26283
rect -11508 26263 -11506 26283
rect -11460 26263 -11458 26283
rect -11436 26263 -11434 26283
rect -11364 26263 -11362 26283
rect -11340 26263 -11338 26283
rect -11268 26263 -11266 26283
rect -11172 26263 -11170 26283
rect -11124 26263 -11122 26283
rect -11076 26263 -11074 26283
rect -11028 26263 -11026 26283
rect -10788 26263 -10786 26283
rect -10668 26263 -10666 26283
rect -9876 26263 -9874 26283
rect -9753 26280 -9739 26283
rect -9732 26280 -9729 26283
rect -9708 26263 -9706 26283
rect -9612 26263 -9610 26283
rect -9516 26263 -9514 26283
rect -9468 26263 -9466 26283
rect -9420 26263 -9418 26283
rect -9396 26263 -9394 26283
rect -9372 26263 -9370 26283
rect -9300 26263 -9298 26283
rect -9252 26263 -9250 26283
rect -9132 26263 -9130 26283
rect -9084 26263 -9082 26283
rect -9036 26263 -9034 26283
rect -8988 26263 -8986 26283
rect -8940 26263 -8938 26283
rect -8892 26263 -8890 26283
rect -8844 26263 -8842 26283
rect -8604 26263 -8602 26283
rect -8508 26263 -8506 26283
rect -8484 26263 -8482 26283
rect -8388 26263 -8386 26283
rect -8364 26263 -8362 26283
rect -8340 26263 -8338 26283
rect -8303 26278 -8300 26283
rect -8292 26278 -8290 26283
rect -8293 26264 -8290 26278
rect -8268 26263 -8266 26283
rect -8196 26280 -8194 26283
rect -8196 26263 -8193 26280
rect -8100 26263 -8098 26283
rect -8052 26263 -8050 26283
rect -7932 26263 -7930 26283
rect -7785 26280 -7771 26283
rect -7761 26283 10325 26287
rect -7761 26280 -7747 26283
rect -7740 26280 -7737 26283
rect -7692 26263 -7690 26283
rect -7620 26263 -7618 26283
rect -7404 26263 -7402 26283
rect -7356 26263 -7354 26283
rect -7308 26263 -7306 26283
rect -7212 26263 -7210 26283
rect -7188 26263 -7186 26283
rect -7116 26263 -7114 26283
rect -7068 26263 -7066 26283
rect -6972 26263 -6970 26283
rect -6948 26263 -6946 26283
rect -6876 26263 -6874 26283
rect -6852 26263 -6850 26283
rect -6804 26264 -6802 26283
rect -6839 26263 -6781 26264
rect -6780 26263 -6778 26283
rect -6756 26263 -6754 26283
rect -6708 26263 -6706 26283
rect -6695 26278 -6692 26283
rect -6684 26278 -6682 26283
rect -6685 26264 -6682 26278
rect -6660 26263 -6658 26283
rect -6612 26263 -6610 26283
rect -6588 26280 -6586 26283
rect -6588 26263 -6585 26280
rect -6564 26263 -6562 26283
rect -6516 26263 -6514 26283
rect -6492 26263 -6490 26283
rect -6468 26263 -6466 26283
rect -6420 26263 -6418 26283
rect -6396 26263 -6394 26283
rect -6372 26263 -6370 26283
rect -6324 26263 -6322 26283
rect -6300 26263 -6298 26283
rect -6276 26263 -6274 26283
rect -6228 26263 -6226 26283
rect -6180 26263 -6178 26283
rect -6060 26263 -6058 26283
rect -5940 26263 -5938 26283
rect -5892 26263 -5890 26283
rect -5652 26263 -5650 26283
rect -5316 26263 -5314 26283
rect -5268 26263 -5266 26283
rect -5196 26263 -5194 26283
rect -5172 26263 -5170 26283
rect -5100 26263 -5098 26283
rect -5076 26263 -5074 26283
rect -4980 26263 -4978 26283
rect -4956 26263 -4954 26283
rect -4884 26263 -4882 26283
rect -4860 26263 -4858 26283
rect -4788 26263 -4786 26283
rect -4692 26263 -4690 26283
rect -4644 26263 -4642 26283
rect -4596 26263 -4594 26283
rect -4548 26263 -4546 26283
rect -4439 26278 -4436 26283
rect -4428 26278 -4426 26283
rect -4429 26264 -4426 26278
rect -4332 26280 -4330 26283
rect -4332 26263 -4329 26280
rect -4308 26263 -4306 26283
rect -4260 26263 -4258 26283
rect -4212 26263 -4210 26283
rect -4116 26263 -4114 26283
rect -4092 26263 -4090 26283
rect -4020 26263 -4018 26283
rect -3876 26263 -3874 26283
rect -3732 26263 -3730 26283
rect -3588 26263 -3586 26283
rect -3564 26263 -3562 26283
rect -3516 26263 -3514 26283
rect -3492 26263 -3490 26283
rect -3468 26263 -3466 26283
rect -3420 26263 -3418 26283
rect -3324 26263 -3322 26283
rect -3252 26263 -3250 26283
rect -3228 26263 -3226 26283
rect -3156 26263 -3154 26283
rect -3132 26263 -3130 26283
rect -3060 26263 -3058 26283
rect -3012 26263 -3010 26283
rect -2964 26263 -2962 26283
rect -2916 26263 -2914 26283
rect -2892 26263 -2890 26283
rect -2820 26263 -2818 26283
rect -2796 26263 -2794 26283
rect -2748 26263 -2746 26283
rect -2700 26263 -2698 26283
rect -2604 26263 -2602 26283
rect -2580 26263 -2578 26283
rect -2364 26263 -2362 26283
rect -2292 26280 -2290 26283
rect -2292 26263 -2289 26280
rect -2268 26263 -2266 26283
rect -2244 26263 -2242 26283
rect -2172 26263 -2170 26283
rect -2148 26263 -2146 26283
rect -2076 26263 -2074 26283
rect -2052 26263 -2050 26283
rect -1980 26263 -1978 26283
rect -1884 26263 -1882 26283
rect -1836 26263 -1834 26283
rect -1716 26263 -1714 26283
rect -1596 26263 -1594 26283
rect -1572 26263 -1570 26283
rect -1476 26263 -1474 26283
rect -1380 26263 -1378 26283
rect -1356 26263 -1354 26283
rect -1308 26263 -1306 26283
rect -1260 26263 -1258 26283
rect -1140 26263 -1138 26283
rect -852 26263 -850 26283
rect -804 26263 -802 26283
rect -756 26263 -754 26283
rect -708 26263 -706 26283
rect -612 26263 -610 26283
rect -588 26263 -586 26283
rect -540 26263 -538 26283
rect -527 26278 -524 26283
rect -516 26278 -514 26283
rect -517 26264 -514 26278
rect -492 26263 -490 26283
rect -444 26263 -442 26283
rect -396 26263 -394 26283
rect -300 26263 -298 26283
rect -276 26263 -274 26283
rect -204 26263 -202 26283
rect -108 26263 -106 26283
rect 12 26263 14 26283
rect 108 26263 110 26283
rect 156 26263 158 26283
rect 204 26263 206 26283
rect 228 26263 230 26283
rect 252 26263 254 26283
rect 348 26263 350 26283
rect 468 26263 470 26283
rect 492 26263 494 26283
rect 564 26263 566 26283
rect 588 26263 590 26283
rect 636 26263 638 26283
rect 660 26263 662 26283
rect 732 26263 734 26283
rect 756 26263 758 26283
rect 876 26263 878 26283
rect 972 26263 974 26283
rect 1020 26263 1022 26283
rect 1068 26263 1070 26283
rect 1092 26263 1094 26283
rect 1116 26263 1118 26283
rect 1164 26263 1166 26283
rect 1212 26263 1214 26283
rect 1308 26263 1310 26283
rect 1332 26263 1334 26283
rect 1380 26263 1382 26283
rect 1428 26263 1430 26283
rect 1524 26263 1526 26283
rect 1548 26263 1550 26283
rect 1596 26263 1598 26283
rect 1620 26263 1622 26283
rect 1644 26263 1646 26283
rect 1692 26263 1694 26283
rect 1716 26263 1718 26283
rect 1740 26263 1742 26283
rect 1788 26263 1790 26283
rect 1884 26263 1886 26283
rect 1980 26263 1982 26283
rect 2028 26263 2030 26283
rect 2076 26263 2078 26283
rect 2100 26263 2102 26283
rect 2124 26263 2126 26283
rect 2172 26263 2174 26283
rect 2196 26263 2198 26283
rect 2220 26263 2222 26283
rect 2268 26263 2270 26283
rect 2292 26263 2294 26283
rect 2316 26263 2318 26283
rect 2364 26263 2366 26283
rect 2412 26263 2414 26283
rect 2460 26263 2462 26283
rect 2508 26263 2510 26283
rect 2556 26263 2558 26283
rect 2580 26263 2582 26283
rect 2604 26263 2606 26283
rect 2652 26263 2654 26283
rect 2676 26263 2678 26283
rect 2700 26263 2702 26283
rect 2748 26263 2750 26283
rect 2772 26263 2774 26283
rect 2796 26263 2798 26283
rect 2844 26263 2846 26283
rect 2868 26263 2870 26283
rect 2892 26263 2894 26283
rect 2940 26263 2942 26283
rect 3012 26263 3014 26283
rect 3108 26263 3110 26283
rect 3156 26263 3158 26283
rect 3252 26263 3254 26283
rect 3348 26263 3350 26283
rect 3396 26263 3398 26283
rect 3468 26263 3470 26283
rect 3492 26263 3494 26283
rect 3588 26263 3590 26283
rect 3612 26263 3614 26283
rect 3636 26263 3638 26283
rect 3708 26263 3710 26283
rect 3732 26263 3734 26283
rect 3804 26263 3806 26283
rect 3828 26263 3830 26283
rect 3924 26263 3926 26283
rect 4020 26263 4022 26283
rect 4044 26263 4046 26283
rect 4092 26263 4094 26283
rect 4116 26263 4118 26283
rect 4140 26263 4142 26283
rect 4188 26263 4190 26283
rect 4212 26263 4214 26283
rect 4236 26263 4238 26283
rect 4308 26263 4310 26283
rect 4332 26263 4334 26283
rect 4404 26263 4406 26283
rect 4500 26263 4502 26283
rect 4596 26263 4598 26283
rect 4860 26263 4862 26283
rect 4956 26263 4958 26283
rect 4980 26263 4982 26283
rect 5004 26263 5006 26283
rect 5076 26263 5078 26283
rect 5100 26263 5102 26283
rect 5124 26263 5126 26283
rect 5172 26263 5174 26283
rect 5196 26263 5198 26283
rect 5220 26263 5222 26283
rect 5268 26263 5270 26283
rect 5292 26263 5294 26283
rect 5388 26263 5390 26283
rect 5484 26263 5486 26283
rect 5508 26263 5510 26283
rect 5532 26263 5534 26283
rect 5628 26263 5630 26283
rect 5652 26263 5654 26283
rect 5748 26263 5750 26283
rect 5796 26263 5798 26283
rect 5844 26263 5846 26283
rect 5892 26263 5894 26283
rect 6132 26263 6134 26283
rect 6180 26263 6182 26283
rect 6228 26263 6230 26283
rect 6252 26263 6254 26283
rect 6276 26263 6278 26283
rect 6324 26263 6326 26283
rect 6372 26263 6374 26283
rect 6492 26263 6494 26283
rect 6588 26263 6590 26283
rect 6612 26263 6614 26283
rect 6660 26263 6662 26283
rect 6684 26263 6686 26283
rect 6708 26263 6710 26283
rect 6780 26263 6782 26283
rect 6804 26263 6806 26283
rect 6828 26263 6830 26283
rect 6900 26263 6902 26283
rect 6924 26263 6926 26283
rect 7020 26263 7022 26283
rect 7140 26263 7142 26283
rect 7236 26263 7238 26283
rect 7332 26263 7334 26283
rect 7380 26263 7382 26283
rect 7428 26263 7430 26283
rect 7452 26263 7454 26283
rect 7476 26263 7478 26283
rect 7524 26263 7526 26283
rect 7548 26263 7550 26283
rect 7572 26263 7574 26283
rect 7620 26263 7622 26283
rect 7644 26263 7646 26283
rect 7668 26263 7670 26283
rect 7716 26263 7718 26283
rect 7740 26263 7742 26283
rect 7836 26263 7838 26283
rect 7884 26263 7886 26283
rect 7932 26263 7934 26283
rect 7956 26263 7958 26283
rect 7980 26263 7982 26283
rect 8028 26263 8030 26283
rect 8196 26263 8198 26283
rect 8244 26263 8246 26283
rect 8268 26263 8270 26283
rect 8292 26263 8294 26283
rect 8340 26263 8342 26283
rect 8364 26263 8366 26283
rect 8388 26263 8390 26283
rect 8436 26263 8438 26283
rect 8460 26263 8462 26283
rect 8556 26263 8558 26283
rect 8604 26263 8606 26283
rect 8652 26263 8654 26283
rect 8700 26263 8702 26283
rect 8724 26263 8726 26283
rect 8748 26263 8750 26283
rect 8820 26263 8822 26283
rect 8844 26263 8846 26283
rect 8868 26263 8870 26283
rect 9516 26263 9518 26283
rect 9612 26263 9614 26283
rect 9660 26263 9662 26283
rect 9684 26263 9686 26283
rect 9708 26263 9710 26283
rect 9756 26263 9758 26283
rect 9780 26263 9782 26283
rect 9804 26263 9806 26283
rect 9852 26263 9854 26283
rect 9876 26263 9878 26283
rect 9900 26263 9902 26283
rect 9948 26263 9950 26283
rect 9972 26263 9974 26283
rect 9996 26263 9998 26283
rect 10068 26263 10070 26283
rect 10092 26263 10094 26283
rect 10116 26263 10118 26283
rect 10164 26263 10166 26283
rect 10188 26263 10190 26283
rect 10212 26263 10214 26283
rect 10284 26263 10286 26283
rect 10308 26263 10310 26283
rect 10311 26280 10325 26283
rect 10332 26283 25397 26287
rect 10332 26280 10349 26283
rect 10332 26263 10334 26280
rect 10380 26263 10382 26283
rect 10404 26263 10406 26283
rect 10428 26263 10430 26283
rect 10476 26263 10478 26283
rect 10500 26263 10502 26283
rect 10524 26263 10526 26283
rect 10572 26263 10574 26283
rect 10596 26263 10598 26283
rect 10620 26263 10622 26283
rect 10668 26263 10670 26283
rect 10692 26263 10694 26283
rect 10716 26263 10718 26283
rect 10788 26263 10790 26283
rect 10836 26263 10838 26283
rect 10956 26263 10958 26283
rect 11052 26263 11054 26283
rect 11076 26263 11078 26283
rect 11124 26263 11126 26283
rect 11172 26263 11174 26283
rect 11220 26263 11222 26283
rect 11340 26263 11342 26283
rect 11436 26263 11438 26283
rect 11532 26263 11534 26283
rect 11580 26263 11582 26283
rect 11628 26263 11630 26283
rect 11676 26263 11678 26283
rect 11713 26278 11716 26283
rect 11723 26264 11726 26278
rect 11724 26263 11726 26264
rect 11772 26263 11774 26283
rect 11796 26263 11798 26283
rect 11844 26280 11846 26283
rect 11844 26263 11847 26280
rect 11892 26263 11894 26283
rect 11988 26263 11990 26283
rect 12060 26263 12062 26283
rect 12132 26263 12134 26283
rect 12228 26263 12230 26283
rect 12276 26263 12278 26283
rect 12324 26263 12326 26283
rect 12420 26263 12422 26283
rect 12444 26263 12446 26283
rect 12492 26263 12494 26283
rect 12516 26263 12518 26283
rect 12540 26263 12542 26283
rect 12588 26263 12590 26283
rect 12636 26263 12638 26283
rect 12732 26263 12734 26283
rect 12756 26263 12758 26283
rect 12804 26263 12806 26283
rect 12828 26263 12830 26283
rect 12852 26263 12854 26283
rect 12900 26263 12902 26283
rect 12948 26263 12950 26283
rect 13044 26263 13046 26283
rect 13068 26263 13070 26283
rect 13116 26263 13118 26283
rect 13284 26263 13286 26283
rect 13332 26263 13334 26283
rect 13428 26263 13430 26283
rect 13524 26263 13526 26283
rect 13572 26263 13574 26283
rect 13644 26263 13646 26283
rect 13668 26263 13670 26283
rect 13764 26263 13766 26283
rect 13812 26263 13814 26283
rect 13860 26263 13862 26283
rect 13908 26263 13910 26283
rect 13956 26263 13958 26283
rect 14004 26263 14006 26283
rect 14100 26263 14102 26283
rect 14196 26263 14198 26283
rect 14244 26280 14246 26283
rect 14244 26263 14247 26280
rect 14292 26263 14294 26283
rect 15132 26263 15134 26283
rect 15180 26263 15182 26283
rect 15228 26263 15230 26283
rect 15252 26263 15254 26283
rect 15324 26263 15326 26283
rect 15396 26263 15398 26283
rect 15420 26263 15422 26283
rect 15492 26263 15494 26283
rect 15540 26263 15542 26283
rect 15636 26263 15638 26283
rect 15660 26263 15662 26283
rect 15708 26263 15710 26283
rect 15732 26263 15734 26283
rect 15756 26263 15758 26283
rect 15804 26263 15806 26283
rect 15828 26263 15830 26283
rect 15852 26263 15854 26283
rect 15900 26263 15902 26283
rect 15948 26263 15950 26283
rect 15996 26263 15998 26283
rect 16044 26263 16046 26283
rect 16092 26263 16094 26283
rect 16140 26264 16142 26283
rect 16129 26263 16163 26264
rect 16236 26263 16238 26283
rect 16260 26263 16262 26283
rect 16308 26263 16310 26283
rect 16332 26263 16334 26283
rect 16356 26263 16358 26283
rect 16404 26263 16406 26283
rect 16452 26263 16454 26283
rect 16548 26263 16550 26283
rect 16572 26263 16574 26283
rect 16620 26263 16622 26283
rect 16668 26263 16670 26283
rect 16716 26263 16718 26283
rect 16764 26263 16766 26283
rect 16836 26263 16838 26283
rect 16884 26263 16886 26283
rect 16980 26263 16982 26283
rect 17052 26263 17054 26283
rect 17196 26263 17198 26283
rect 17220 26263 17222 26283
rect 17292 26263 17294 26283
rect 17316 26263 17318 26283
rect 18084 26263 18086 26283
rect 18132 26263 18134 26283
rect 18396 26263 18398 26283
rect 18492 26263 18494 26283
rect 18516 26263 18518 26283
rect 18564 26263 18566 26283
rect 18612 26263 18614 26283
rect 18660 26263 18662 26283
rect 18708 26263 18710 26283
rect 18756 26263 18758 26283
rect 18804 26263 18806 26283
rect 18852 26263 18854 26283
rect 18900 26263 18902 26283
rect 18996 26263 18998 26283
rect 19020 26263 19022 26283
rect 19092 26263 19094 26283
rect 19116 26263 19118 26283
rect 19140 26263 19142 26283
rect 19188 26263 19190 26283
rect 19236 26263 19238 26283
rect 19332 26263 19334 26283
rect 19476 26263 19478 26283
rect 19620 26263 19622 26283
rect 19716 26263 19718 26283
rect 19788 26263 19790 26283
rect 19836 26263 19838 26283
rect 19860 26263 19862 26283
rect 19884 26263 19886 26283
rect 19932 26263 19934 26283
rect 19956 26263 19958 26283
rect 19980 26263 19982 26283
rect 20028 26263 20030 26283
rect 20052 26263 20054 26283
rect 20076 26263 20078 26283
rect 20148 26263 20150 26283
rect 20172 26263 20174 26283
rect 20196 26263 20198 26283
rect 20268 26263 20270 26283
rect 20292 26263 20294 26283
rect 20388 26263 20390 26283
rect 20412 26263 20414 26283
rect 20508 26263 20510 26283
rect 20556 26263 20558 26283
rect 20604 26263 20606 26283
rect 20916 26263 20918 26283
rect 20964 26263 20966 26283
rect 21012 26263 21014 26283
rect 21060 26263 21062 26283
rect 21084 26263 21086 26283
rect 21108 26263 21110 26283
rect 21204 26263 21206 26283
rect 21300 26263 21302 26283
rect 21324 26263 21326 26283
rect 21444 26263 21446 26283
rect 21468 26263 21470 26283
rect 21564 26263 21566 26283
rect 21612 26263 21614 26283
rect 21684 26263 21686 26283
rect 21708 26263 21710 26283
rect 21793 26278 21796 26283
rect 21804 26278 21806 26283
rect 21803 26264 21806 26278
rect 21828 26263 21830 26283
rect 21924 26263 21926 26283
rect 21948 26263 21950 26283
rect 22044 26263 22046 26283
rect 22068 26263 22070 26283
rect 22188 26263 22190 26283
rect 22212 26263 22214 26283
rect 23004 26263 23006 26283
rect 23052 26263 23054 26283
rect 23076 26263 23078 26283
rect 23100 26263 23102 26283
rect 23148 26263 23150 26283
rect 23220 26263 23222 26283
rect 23244 26263 23246 26283
rect 23316 26263 23318 26283
rect 23340 26263 23342 26283
rect 23412 26263 23414 26283
rect 23556 26263 23558 26283
rect 23628 26263 23630 26283
rect 23652 26263 23654 26283
rect 23676 26263 23678 26283
rect 23724 26263 23726 26283
rect 23772 26263 23774 26283
rect 23820 26263 23822 26283
rect 23868 26263 23870 26283
rect 23916 26263 23918 26283
rect 24012 26263 24014 26283
rect 24084 26263 24086 26283
rect 24372 26263 24374 26283
rect 24396 26263 24398 26283
rect 24492 26263 24494 26283
rect 24516 26263 24518 26283
rect 24588 26263 24590 26283
rect 24612 26263 24614 26283
rect 24708 26263 24710 26283
rect 24732 26263 24734 26283
rect 24756 26263 24758 26283
rect 24852 26263 24854 26283
rect 24876 26263 24878 26283
rect 24972 26263 24974 26283
rect 24996 26263 24998 26283
rect 25092 26263 25094 26283
rect 25260 26263 25262 26283
rect 25308 26263 25310 26283
rect 25356 26263 25358 26283
rect 25380 26263 25382 26283
rect 25383 26280 25397 26283
rect 25404 26283 27245 26287
rect 25404 26280 25421 26283
rect 25404 26263 25406 26280
rect 25452 26263 25454 26283
rect 25500 26263 25502 26283
rect 25596 26263 25598 26283
rect 27060 26263 27062 26283
rect 27108 26263 27110 26283
rect 27156 26263 27158 26283
rect 27231 26280 27245 26283
rect 27255 26283 31091 26287
rect 27255 26280 27269 26283
rect 27324 26263 27326 26283
rect 27396 26263 27398 26283
rect 27420 26263 27422 26283
rect 27540 26263 27542 26283
rect 27564 26263 27566 26283
rect 30564 26263 30566 26283
rect 30636 26263 30638 26283
rect 30660 26263 30662 26283
rect 30780 26263 30782 26283
rect 30804 26263 30806 26283
rect 30924 26280 30926 26283
rect 30924 26263 30927 26280
rect 30948 26263 30950 26283
rect 31057 26278 31060 26283
rect 31068 26278 31070 26283
rect 31067 26264 31070 26278
rect 30985 26263 31019 26264
rect -17337 26259 -16195 26263
rect -17337 26256 -17323 26259
rect -17457 26239 -17437 26240
rect -17436 26239 -17433 26256
rect -17388 26239 -17386 26256
rect -17292 26239 -17290 26259
rect -17196 26239 -17194 26259
rect -17028 26239 -17026 26259
rect -16932 26239 -16930 26259
rect -16860 26239 -16858 26259
rect -16836 26239 -16834 26259
rect -16764 26239 -16762 26259
rect -16740 26239 -16738 26259
rect -16668 26239 -16666 26259
rect -16500 26239 -16498 26259
rect -16380 26239 -16378 26259
rect -16356 26239 -16354 26259
rect -16284 26239 -16282 26259
rect -16260 26239 -16258 26259
rect -16236 26239 -16234 26259
rect -16209 26256 -16195 26259
rect -16137 26259 11813 26263
rect -16137 26256 -16123 26259
rect -15300 26239 -15298 26259
rect -15143 26239 -15109 26240
rect -15084 26239 -15082 26259
rect -15036 26239 -15034 26259
rect -14868 26239 -14866 26259
rect -14772 26239 -14770 26259
rect -14724 26239 -14722 26259
rect -14508 26239 -14506 26259
rect -14436 26239 -14434 26259
rect -14399 26254 -14396 26259
rect -14388 26254 -14386 26259
rect -14351 26254 -14348 26259
rect -14389 26240 -14386 26254
rect -14341 26240 -14338 26254
rect -14303 26246 -14299 26254
rect -14313 26240 -14303 26246
rect -14340 26239 -14338 26240
rect -14244 26239 -14241 26256
rect -14172 26239 -14170 26259
rect -14076 26239 -14074 26259
rect -13980 26239 -13978 26259
rect -13932 26239 -13930 26259
rect -13884 26239 -13882 26259
rect -13716 26239 -13714 26259
rect -13644 26239 -13642 26259
rect -13596 26239 -13594 26259
rect -13500 26239 -13498 26259
rect -13404 26240 -13402 26259
rect -13439 26239 -13381 26240
rect -13356 26239 -13354 26259
rect -13284 26239 -13282 26259
rect -13068 26239 -13066 26259
rect -12828 26239 -12826 26259
rect -12780 26239 -12778 26259
rect -12660 26239 -12658 26259
rect -12564 26239 -12562 26259
rect -12492 26239 -12490 26259
rect -12396 26239 -12394 26259
rect -12348 26239 -12346 26259
rect -12276 26239 -12274 26259
rect -12252 26239 -12250 26259
rect -12156 26239 -12154 26259
rect -12060 26239 -12058 26259
rect -11892 26239 -11890 26259
rect -11844 26239 -11842 26259
rect -11796 26239 -11794 26259
rect -11676 26239 -11674 26259
rect -11580 26239 -11578 26259
rect -11556 26239 -11554 26259
rect -11508 26239 -11506 26259
rect -11460 26239 -11458 26259
rect -11436 26239 -11434 26259
rect -11364 26239 -11362 26259
rect -11340 26239 -11338 26259
rect -11268 26239 -11266 26259
rect -11172 26239 -11170 26259
rect -11124 26239 -11122 26259
rect -11076 26239 -11074 26259
rect -11028 26239 -11026 26259
rect -10788 26239 -10786 26259
rect -10668 26239 -10666 26259
rect -10487 26239 -10429 26240
rect -9876 26239 -9874 26259
rect -9708 26239 -9706 26259
rect -9612 26239 -9610 26259
rect -9516 26239 -9514 26259
rect -9468 26239 -9466 26259
rect -9420 26239 -9418 26259
rect -9396 26239 -9394 26259
rect -9372 26239 -9370 26259
rect -9300 26239 -9298 26259
rect -9252 26239 -9250 26259
rect -9132 26239 -9130 26259
rect -9084 26239 -9082 26259
rect -9036 26239 -9034 26259
rect -8988 26239 -8986 26259
rect -8940 26239 -8938 26259
rect -8892 26239 -8890 26259
rect -8844 26239 -8842 26259
rect -8604 26239 -8602 26259
rect -8508 26239 -8506 26259
rect -8484 26239 -8482 26259
rect -8388 26239 -8386 26259
rect -8364 26239 -8362 26259
rect -8340 26239 -8338 26259
rect -8268 26239 -8266 26259
rect -8217 26256 -8203 26259
rect -8196 26256 -8193 26259
rect -8100 26239 -8098 26259
rect -8052 26239 -8050 26259
rect -7932 26239 -7930 26259
rect -7692 26239 -7690 26259
rect -7620 26239 -7618 26259
rect -7404 26239 -7402 26259
rect -7356 26239 -7354 26259
rect -7308 26239 -7306 26259
rect -7212 26239 -7210 26259
rect -7188 26239 -7186 26259
rect -7116 26239 -7114 26259
rect -7068 26239 -7066 26259
rect -6972 26239 -6970 26259
rect -6948 26239 -6946 26259
rect -6876 26239 -6874 26259
rect -6852 26239 -6850 26259
rect -6815 26254 -6812 26259
rect -6804 26254 -6802 26259
rect -6805 26240 -6802 26254
rect -6780 26239 -6778 26259
rect -6756 26239 -6754 26259
rect -6708 26256 -6706 26259
rect -6708 26239 -6705 26256
rect -6660 26239 -6658 26259
rect -6612 26239 -6610 26259
rect -6609 26256 -6595 26259
rect -6588 26256 -6585 26259
rect -6564 26239 -6562 26259
rect -6516 26239 -6514 26259
rect -6492 26239 -6490 26259
rect -6468 26239 -6466 26259
rect -6420 26239 -6418 26259
rect -6396 26239 -6394 26259
rect -6372 26239 -6370 26259
rect -6324 26239 -6322 26259
rect -6300 26239 -6298 26259
rect -6276 26239 -6274 26259
rect -6228 26239 -6226 26259
rect -6180 26239 -6178 26259
rect -6060 26239 -6058 26259
rect -5940 26239 -5938 26259
rect -5892 26239 -5890 26259
rect -5652 26239 -5650 26259
rect -5316 26240 -5314 26259
rect -5351 26239 -5293 26240
rect -5268 26239 -5266 26259
rect -5196 26239 -5194 26259
rect -5172 26239 -5170 26259
rect -5100 26239 -5098 26259
rect -5076 26239 -5074 26259
rect -4980 26239 -4978 26259
rect -4956 26239 -4954 26259
rect -4884 26239 -4882 26259
rect -4860 26239 -4858 26259
rect -4788 26239 -4786 26259
rect -4692 26239 -4690 26259
rect -4644 26239 -4642 26259
rect -4596 26239 -4594 26259
rect -4548 26239 -4546 26259
rect -4353 26256 -4339 26259
rect -4332 26256 -4329 26259
rect -4308 26239 -4306 26259
rect -4260 26239 -4258 26259
rect -4212 26239 -4210 26259
rect -4116 26239 -4114 26259
rect -4092 26239 -4090 26259
rect -4020 26239 -4018 26259
rect -3876 26239 -3874 26259
rect -3732 26239 -3730 26259
rect -3588 26239 -3586 26259
rect -3564 26239 -3562 26259
rect -3516 26239 -3514 26259
rect -3492 26239 -3490 26259
rect -3468 26239 -3466 26259
rect -3420 26239 -3418 26259
rect -3324 26239 -3322 26259
rect -3252 26239 -3250 26259
rect -3228 26239 -3226 26259
rect -3156 26239 -3154 26259
rect -3132 26239 -3130 26259
rect -3060 26239 -3058 26259
rect -3012 26239 -3010 26259
rect -2964 26239 -2962 26259
rect -2916 26239 -2914 26259
rect -2892 26239 -2890 26259
rect -2820 26239 -2818 26259
rect -2796 26239 -2794 26259
rect -2748 26239 -2746 26259
rect -2700 26239 -2698 26259
rect -2604 26239 -2602 26259
rect -2580 26239 -2578 26259
rect -2364 26239 -2362 26259
rect -2313 26256 -2299 26259
rect -2292 26256 -2289 26259
rect -2268 26239 -2266 26259
rect -2244 26239 -2242 26259
rect -2172 26239 -2170 26259
rect -2148 26239 -2146 26259
rect -2076 26239 -2074 26259
rect -2052 26239 -2050 26259
rect -1980 26239 -1978 26259
rect -1884 26239 -1882 26259
rect -1836 26239 -1834 26259
rect -1716 26239 -1714 26259
rect -1596 26239 -1594 26259
rect -1572 26239 -1570 26259
rect -1476 26239 -1474 26259
rect -1380 26239 -1378 26259
rect -1356 26239 -1354 26259
rect -1308 26239 -1306 26259
rect -1260 26239 -1258 26259
rect -1140 26239 -1138 26259
rect -852 26239 -850 26259
rect -804 26239 -802 26259
rect -756 26239 -754 26259
rect -708 26239 -706 26259
rect -612 26239 -610 26259
rect -588 26239 -586 26259
rect -540 26239 -538 26259
rect -492 26239 -490 26259
rect -444 26239 -442 26259
rect -441 26256 -427 26259
rect -396 26239 -394 26259
rect -300 26239 -298 26259
rect -276 26239 -274 26259
rect -204 26239 -202 26259
rect -108 26239 -106 26259
rect 12 26239 14 26259
rect 108 26239 110 26259
rect 156 26239 158 26259
rect 204 26239 206 26259
rect 228 26239 230 26259
rect 252 26239 254 26259
rect 348 26239 350 26259
rect 468 26239 470 26259
rect 492 26239 494 26259
rect 564 26239 566 26259
rect 588 26239 590 26259
rect 636 26239 638 26259
rect 660 26239 662 26259
rect 732 26239 734 26259
rect 756 26239 758 26259
rect 876 26239 878 26259
rect 972 26239 974 26259
rect 1020 26239 1022 26259
rect 1068 26239 1070 26259
rect 1092 26239 1094 26259
rect 1116 26239 1118 26259
rect 1164 26239 1166 26259
rect 1212 26239 1214 26259
rect 1308 26239 1310 26259
rect 1332 26239 1334 26259
rect 1380 26239 1382 26259
rect 1428 26239 1430 26259
rect 1524 26239 1526 26259
rect 1548 26239 1550 26259
rect 1596 26239 1598 26259
rect 1620 26239 1622 26259
rect 1644 26239 1646 26259
rect 1692 26239 1694 26259
rect 1716 26239 1718 26259
rect 1740 26239 1742 26259
rect 1788 26239 1790 26259
rect 1884 26239 1886 26259
rect 1980 26239 1982 26259
rect 2028 26239 2030 26259
rect 2076 26239 2078 26259
rect 2100 26239 2102 26259
rect 2124 26239 2126 26259
rect 2172 26239 2174 26259
rect 2196 26239 2198 26259
rect 2220 26239 2222 26259
rect 2268 26239 2270 26259
rect 2292 26239 2294 26259
rect 2316 26239 2318 26259
rect 2364 26239 2366 26259
rect 2412 26239 2414 26259
rect 2460 26239 2462 26259
rect 2508 26239 2510 26259
rect 2556 26239 2558 26259
rect 2580 26239 2582 26259
rect 2604 26239 2606 26259
rect 2652 26239 2654 26259
rect 2676 26239 2678 26259
rect 2700 26239 2702 26259
rect 2748 26239 2750 26259
rect 2772 26239 2774 26259
rect 2796 26239 2798 26259
rect 2844 26239 2846 26259
rect 2868 26239 2870 26259
rect 2892 26239 2894 26259
rect 2940 26239 2942 26259
rect 3012 26239 3014 26259
rect 3108 26239 3110 26259
rect 3156 26239 3158 26259
rect 3252 26239 3254 26259
rect 3348 26239 3350 26259
rect 3396 26239 3398 26259
rect 3468 26239 3470 26259
rect 3492 26239 3494 26259
rect 3588 26239 3590 26259
rect 3612 26239 3614 26259
rect 3636 26239 3638 26259
rect 3708 26239 3710 26259
rect 3732 26239 3734 26259
rect 3804 26239 3806 26259
rect 3828 26239 3830 26259
rect 3924 26239 3926 26259
rect 4020 26239 4022 26259
rect 4044 26239 4046 26259
rect 4092 26239 4094 26259
rect 4116 26239 4118 26259
rect 4140 26239 4142 26259
rect 4188 26239 4190 26259
rect 4212 26239 4214 26259
rect 4236 26239 4238 26259
rect 4308 26239 4310 26259
rect 4332 26239 4334 26259
rect 4404 26239 4406 26259
rect 4500 26239 4502 26259
rect 4596 26239 4598 26259
rect 4860 26239 4862 26259
rect 4956 26239 4958 26259
rect 4980 26239 4982 26259
rect 5004 26239 5006 26259
rect 5076 26239 5078 26259
rect 5100 26239 5102 26259
rect 5124 26239 5126 26259
rect 5172 26239 5174 26259
rect 5196 26239 5198 26259
rect 5220 26239 5222 26259
rect 5268 26239 5270 26259
rect 5292 26239 5294 26259
rect 5388 26239 5390 26259
rect 5484 26239 5486 26259
rect 5508 26239 5510 26259
rect 5532 26239 5534 26259
rect 5628 26239 5630 26259
rect 5652 26239 5654 26259
rect 5748 26239 5750 26259
rect 5796 26239 5798 26259
rect 5844 26239 5846 26259
rect 5892 26239 5894 26259
rect 6132 26239 6134 26259
rect 6180 26239 6182 26259
rect 6228 26239 6230 26259
rect 6252 26239 6254 26259
rect 6276 26239 6278 26259
rect 6324 26239 6326 26259
rect 6372 26239 6374 26259
rect 6492 26239 6494 26259
rect 6588 26239 6590 26259
rect 6612 26239 6614 26259
rect 6660 26239 6662 26259
rect 6684 26239 6686 26259
rect 6708 26239 6710 26259
rect 6780 26239 6782 26259
rect 6804 26239 6806 26259
rect 6828 26239 6830 26259
rect 6900 26239 6902 26259
rect 6924 26239 6926 26259
rect 7020 26239 7022 26259
rect 7140 26239 7142 26259
rect 7236 26239 7238 26259
rect 7332 26239 7334 26259
rect 7380 26239 7382 26259
rect 7428 26239 7430 26259
rect 7452 26239 7454 26259
rect 7476 26239 7478 26259
rect 7524 26239 7526 26259
rect 7548 26239 7550 26259
rect 7572 26239 7574 26259
rect 7620 26239 7622 26259
rect 7644 26239 7646 26259
rect 7668 26239 7670 26259
rect 7716 26239 7718 26259
rect 7740 26239 7742 26259
rect 7836 26239 7838 26259
rect 7884 26239 7886 26259
rect 7932 26239 7934 26259
rect 7956 26239 7958 26259
rect 7980 26239 7982 26259
rect 8028 26239 8030 26259
rect 8196 26239 8198 26259
rect 8244 26239 8246 26259
rect 8268 26239 8270 26259
rect 8292 26239 8294 26259
rect 8340 26239 8342 26259
rect 8364 26239 8366 26259
rect 8388 26239 8390 26259
rect 8436 26239 8438 26259
rect 8460 26239 8462 26259
rect 8556 26239 8558 26259
rect 8604 26239 8606 26259
rect 8652 26239 8654 26259
rect 8700 26239 8702 26259
rect 8724 26239 8726 26259
rect 8748 26239 8750 26259
rect 8820 26239 8822 26259
rect 8844 26239 8846 26259
rect 8868 26239 8870 26259
rect 9516 26239 9518 26259
rect 9612 26239 9614 26259
rect 9660 26239 9662 26259
rect 9684 26239 9686 26259
rect 9708 26239 9710 26259
rect 9756 26239 9758 26259
rect 9780 26239 9782 26259
rect 9804 26239 9806 26259
rect 9852 26239 9854 26259
rect 9876 26239 9878 26259
rect 9900 26239 9902 26259
rect 9948 26239 9950 26259
rect 9972 26239 9974 26259
rect 9996 26239 9998 26259
rect 10068 26239 10070 26259
rect 10092 26239 10094 26259
rect 10116 26239 10118 26259
rect 10164 26239 10166 26259
rect 10188 26239 10190 26259
rect 10212 26239 10214 26259
rect 10284 26239 10286 26259
rect 10308 26239 10310 26259
rect 10332 26239 10334 26259
rect 10380 26239 10382 26259
rect 10404 26239 10406 26259
rect 10428 26239 10430 26259
rect 10476 26239 10478 26259
rect 10500 26239 10502 26259
rect 10524 26239 10526 26259
rect 10572 26239 10574 26259
rect 10596 26239 10598 26259
rect 10620 26239 10622 26259
rect 10668 26239 10670 26259
rect 10692 26239 10694 26259
rect 10716 26239 10718 26259
rect 10788 26239 10790 26259
rect 10836 26239 10838 26259
rect 10956 26239 10958 26259
rect 11052 26239 11054 26259
rect 11076 26239 11078 26259
rect 11124 26239 11126 26259
rect 11172 26239 11174 26259
rect 11220 26239 11222 26259
rect 11340 26239 11342 26259
rect 11436 26239 11438 26259
rect 11532 26239 11534 26259
rect 11580 26239 11582 26259
rect 11628 26239 11630 26259
rect 11676 26239 11678 26259
rect 11724 26239 11726 26259
rect 11772 26239 11774 26259
rect 11796 26239 11798 26259
rect 11799 26256 11813 26259
rect 11823 26259 31019 26263
rect 11823 26256 11837 26259
rect 11844 26256 11847 26259
rect 11892 26239 11894 26259
rect 11988 26239 11990 26259
rect 12060 26239 12062 26259
rect 12132 26239 12134 26259
rect 12228 26239 12230 26259
rect 12276 26239 12278 26259
rect 12324 26239 12326 26259
rect 12420 26239 12422 26259
rect 12444 26239 12446 26259
rect 12492 26239 12494 26259
rect 12516 26239 12518 26259
rect 12540 26239 12542 26259
rect 12588 26239 12590 26259
rect 12636 26239 12638 26259
rect 12732 26239 12734 26259
rect 12756 26239 12758 26259
rect 12804 26239 12806 26259
rect 12828 26239 12830 26259
rect 12852 26239 12854 26259
rect 12900 26239 12902 26259
rect 12948 26239 12950 26259
rect 13044 26239 13046 26259
rect 13068 26239 13070 26259
rect 13116 26239 13118 26259
rect 13284 26239 13286 26259
rect 13332 26239 13334 26259
rect 13428 26239 13430 26259
rect 13524 26239 13526 26259
rect 13572 26239 13574 26259
rect 13644 26239 13646 26259
rect 13668 26239 13670 26259
rect 13764 26239 13766 26259
rect 13812 26239 13814 26259
rect 13860 26239 13862 26259
rect 13908 26239 13910 26259
rect 13956 26239 13958 26259
rect 14004 26239 14006 26259
rect 14100 26239 14102 26259
rect 14196 26239 14198 26259
rect 14223 26256 14237 26259
rect 14244 26256 14247 26259
rect 14292 26239 14294 26259
rect 15132 26239 15134 26259
rect 15180 26239 15182 26259
rect 15228 26239 15230 26259
rect 15252 26239 15254 26259
rect 15324 26239 15326 26259
rect 15396 26239 15398 26259
rect 15420 26239 15422 26259
rect 15492 26239 15494 26259
rect 15540 26239 15542 26259
rect 15636 26239 15638 26259
rect 15660 26239 15662 26259
rect 15708 26239 15710 26259
rect 15732 26239 15734 26259
rect 15756 26239 15758 26259
rect 15804 26239 15806 26259
rect 15828 26239 15830 26259
rect 15852 26239 15854 26259
rect 15900 26239 15902 26259
rect 15948 26239 15950 26259
rect 15996 26239 15998 26259
rect 16044 26239 16046 26259
rect 16092 26239 16094 26259
rect 16129 26254 16132 26259
rect 16140 26254 16142 26259
rect 16139 26240 16142 26254
rect 16236 26256 16238 26259
rect 16236 26239 16239 26256
rect 16260 26239 16262 26259
rect 16308 26239 16310 26259
rect 16332 26239 16334 26259
rect 16356 26239 16358 26259
rect 16404 26239 16406 26259
rect 16452 26239 16454 26259
rect 16548 26239 16550 26259
rect 16572 26239 16574 26259
rect 16620 26239 16622 26259
rect 16668 26239 16670 26259
rect 16716 26239 16718 26259
rect 16764 26239 16766 26259
rect 16836 26239 16838 26259
rect 16884 26239 16886 26259
rect 16980 26239 16982 26259
rect 17052 26239 17054 26259
rect 17196 26239 17198 26259
rect 17220 26239 17222 26259
rect 17292 26239 17294 26259
rect 17316 26239 17318 26259
rect 18084 26239 18086 26259
rect 18132 26239 18134 26259
rect 18396 26239 18398 26259
rect 18492 26239 18494 26259
rect 18516 26239 18518 26259
rect 18564 26239 18566 26259
rect 18612 26239 18614 26259
rect 18660 26239 18662 26259
rect 18708 26239 18710 26259
rect 18756 26239 18758 26259
rect 18804 26239 18806 26259
rect 18852 26239 18854 26259
rect 18900 26239 18902 26259
rect 18996 26239 18998 26259
rect 19020 26239 19022 26259
rect 19092 26239 19094 26259
rect 19116 26239 19118 26259
rect 19140 26239 19142 26259
rect 19188 26239 19190 26259
rect 19236 26239 19238 26259
rect 19332 26239 19334 26259
rect 19476 26239 19478 26259
rect 19620 26239 19622 26259
rect 19716 26239 19718 26259
rect 19788 26239 19790 26259
rect 19836 26239 19838 26259
rect 19860 26239 19862 26259
rect 19884 26239 19886 26259
rect 19932 26239 19934 26259
rect 19956 26239 19958 26259
rect 19980 26239 19982 26259
rect 20028 26239 20030 26259
rect 20052 26239 20054 26259
rect 20076 26239 20078 26259
rect 20148 26239 20150 26259
rect 20172 26239 20174 26259
rect 20196 26239 20198 26259
rect 20268 26239 20270 26259
rect 20292 26239 20294 26259
rect 20388 26239 20390 26259
rect 20412 26239 20414 26259
rect 20508 26239 20510 26259
rect 20556 26239 20558 26259
rect 20604 26239 20606 26259
rect 20916 26239 20918 26259
rect 20964 26239 20966 26259
rect 21012 26239 21014 26259
rect 21060 26239 21062 26259
rect 21084 26239 21086 26259
rect 21108 26239 21110 26259
rect 21204 26239 21206 26259
rect 21300 26239 21302 26259
rect 21324 26239 21326 26259
rect 21444 26239 21446 26259
rect 21468 26239 21470 26259
rect 21564 26239 21566 26259
rect 21612 26239 21614 26259
rect 21684 26239 21686 26259
rect 21708 26239 21710 26259
rect 21828 26239 21830 26259
rect 21879 26256 21893 26259
rect 21924 26239 21926 26259
rect 21948 26239 21950 26259
rect 22044 26239 22046 26259
rect 22068 26239 22070 26259
rect 22188 26239 22190 26259
rect 22212 26239 22214 26259
rect 23004 26239 23006 26259
rect 23052 26239 23054 26259
rect 23076 26239 23078 26259
rect 23100 26239 23102 26259
rect 23148 26239 23150 26259
rect 23220 26239 23222 26259
rect 23244 26239 23246 26259
rect 23316 26239 23318 26259
rect 23340 26239 23342 26259
rect 23412 26239 23414 26259
rect 23556 26239 23558 26259
rect 23628 26239 23630 26259
rect 23652 26239 23654 26259
rect 23676 26239 23678 26259
rect 23724 26239 23726 26259
rect 23772 26239 23774 26259
rect 23820 26239 23822 26259
rect 23868 26239 23870 26259
rect 23916 26239 23918 26259
rect 24012 26239 24014 26259
rect 24084 26239 24086 26259
rect 24372 26239 24374 26259
rect 24396 26239 24398 26259
rect 24492 26239 24494 26259
rect 24516 26239 24518 26259
rect 24588 26239 24590 26259
rect 24612 26239 24614 26259
rect 24708 26239 24710 26259
rect 24732 26239 24734 26259
rect 24756 26239 24758 26259
rect 24852 26239 24854 26259
rect 24876 26239 24878 26259
rect 24972 26239 24974 26259
rect 24996 26239 24998 26259
rect 25092 26239 25094 26259
rect 25119 26256 25133 26259
rect 25260 26239 25262 26259
rect 25308 26239 25310 26259
rect 25356 26239 25358 26259
rect 25380 26239 25382 26259
rect 25404 26239 25406 26259
rect 25452 26239 25454 26259
rect 25500 26239 25502 26259
rect 25596 26239 25598 26259
rect 27060 26239 27062 26259
rect 27108 26239 27110 26259
rect 27156 26239 27158 26259
rect 27324 26239 27326 26259
rect 27396 26239 27398 26259
rect 27420 26239 27422 26259
rect 27540 26239 27542 26259
rect 27564 26239 27566 26259
rect 30564 26239 30566 26259
rect 30636 26239 30638 26259
rect 30660 26239 30662 26259
rect 30780 26239 30782 26259
rect 30804 26239 30806 26259
rect 30903 26256 30917 26259
rect 30924 26256 30927 26259
rect 30948 26239 30950 26259
rect 30961 26239 30995 26240
rect -17457 26235 -14251 26239
rect -17457 26232 -17443 26235
rect -17436 26232 -17433 26235
rect -17461 26216 -17458 26230
rect -17913 26211 -17419 26215
rect -17913 26208 -17899 26211
rect -17844 26208 -17842 26211
rect -17844 26192 -17841 26208
rect -17855 26191 -17821 26192
rect -17508 26191 -17506 26211
rect -17484 26191 -17482 26211
rect -17433 26208 -17419 26211
rect -17388 26191 -17386 26235
rect -17292 26215 -17290 26235
rect -17196 26216 -17194 26235
rect -17207 26215 -17173 26216
rect -17028 26215 -17026 26235
rect -16932 26215 -16930 26235
rect -16860 26215 -16858 26235
rect -16836 26215 -16834 26235
rect -16764 26215 -16762 26235
rect -16740 26215 -16738 26235
rect -16668 26215 -16666 26235
rect -16500 26215 -16498 26235
rect -16380 26215 -16378 26235
rect -16356 26215 -16354 26235
rect -16284 26215 -16282 26235
rect -16260 26215 -16258 26235
rect -16236 26215 -16234 26235
rect -15300 26215 -15298 26235
rect -15084 26215 -15082 26235
rect -15036 26232 -15034 26235
rect -15036 26216 -15033 26232
rect -15047 26215 -15013 26216
rect -14868 26215 -14866 26235
rect -14772 26215 -14770 26235
rect -14724 26215 -14722 26235
rect -14508 26215 -14506 26235
rect -14436 26215 -14434 26235
rect -14340 26215 -14338 26235
rect -14313 26232 -14299 26235
rect -14265 26232 -14251 26235
rect -14244 26235 -6739 26239
rect -14244 26232 -14227 26235
rect -14244 26215 -14242 26232
rect -14172 26215 -14170 26235
rect -14076 26215 -14074 26235
rect -13980 26215 -13978 26235
rect -13932 26215 -13930 26235
rect -13884 26215 -13882 26235
rect -13716 26215 -13714 26235
rect -13703 26215 -13669 26216
rect -13644 26215 -13642 26235
rect -13596 26215 -13594 26235
rect -13500 26215 -13498 26235
rect -13415 26230 -13412 26235
rect -13404 26230 -13402 26235
rect -13405 26216 -13402 26230
rect -13356 26215 -13354 26235
rect -13284 26215 -13282 26235
rect -13068 26215 -13066 26235
rect -12828 26215 -12826 26235
rect -12780 26215 -12778 26235
rect -12660 26215 -12658 26235
rect -12564 26215 -12562 26235
rect -12492 26215 -12490 26235
rect -12396 26215 -12394 26235
rect -12348 26215 -12346 26235
rect -12276 26215 -12274 26235
rect -12252 26215 -12250 26235
rect -12156 26215 -12154 26235
rect -12060 26215 -12058 26235
rect -11892 26215 -11890 26235
rect -11844 26215 -11842 26235
rect -11796 26215 -11794 26235
rect -11676 26215 -11674 26235
rect -11580 26215 -11578 26235
rect -11556 26215 -11554 26235
rect -11508 26215 -11506 26235
rect -11460 26215 -11458 26235
rect -11436 26215 -11434 26235
rect -11364 26215 -11362 26235
rect -11340 26215 -11338 26235
rect -11268 26215 -11266 26235
rect -11172 26215 -11170 26235
rect -11124 26215 -11122 26235
rect -11076 26215 -11074 26235
rect -11028 26215 -11026 26235
rect -10788 26215 -10786 26235
rect -10668 26215 -10666 26235
rect -10007 26215 -9949 26216
rect -9876 26215 -9874 26235
rect -9708 26215 -9706 26235
rect -9612 26215 -9610 26235
rect -9516 26215 -9514 26235
rect -9468 26215 -9466 26235
rect -9420 26215 -9418 26235
rect -9396 26215 -9394 26235
rect -9372 26215 -9370 26235
rect -9300 26215 -9298 26235
rect -9252 26215 -9250 26235
rect -9132 26215 -9130 26235
rect -9084 26215 -9082 26235
rect -9036 26215 -9034 26235
rect -8988 26215 -8986 26235
rect -8940 26215 -8938 26235
rect -8892 26215 -8890 26235
rect -8844 26216 -8842 26235
rect -8879 26215 -8821 26216
rect -8604 26215 -8602 26235
rect -8508 26215 -8506 26235
rect -8484 26215 -8482 26235
rect -8388 26215 -8386 26235
rect -8364 26215 -8362 26235
rect -8340 26215 -8338 26235
rect -8268 26215 -8266 26235
rect -8100 26215 -8098 26235
rect -8052 26215 -8050 26235
rect -7932 26215 -7930 26235
rect -7692 26215 -7690 26235
rect -7620 26215 -7618 26235
rect -7404 26215 -7402 26235
rect -7356 26215 -7354 26235
rect -7308 26215 -7306 26235
rect -7212 26215 -7210 26235
rect -7188 26215 -7186 26235
rect -7116 26215 -7114 26235
rect -7068 26215 -7066 26235
rect -6972 26215 -6970 26235
rect -6948 26215 -6946 26235
rect -6876 26215 -6874 26235
rect -6852 26215 -6850 26235
rect -6780 26215 -6778 26235
rect -6756 26215 -6754 26235
rect -6753 26232 -6739 26235
rect -6729 26235 30995 26239
rect -6729 26232 -6715 26235
rect -6708 26232 -6705 26235
rect -6660 26215 -6658 26235
rect -6612 26215 -6610 26235
rect -6564 26215 -6562 26235
rect -6516 26215 -6514 26235
rect -6492 26215 -6490 26235
rect -6468 26215 -6466 26235
rect -6420 26215 -6418 26235
rect -6396 26215 -6394 26235
rect -6372 26215 -6370 26235
rect -6324 26215 -6322 26235
rect -6300 26215 -6298 26235
rect -6276 26215 -6274 26235
rect -6228 26215 -6226 26235
rect -6180 26215 -6178 26235
rect -6060 26215 -6058 26235
rect -5940 26215 -5938 26235
rect -5892 26215 -5890 26235
rect -5652 26215 -5650 26235
rect -5327 26230 -5324 26235
rect -5316 26230 -5314 26235
rect -5317 26216 -5314 26230
rect -5268 26215 -5266 26235
rect -5196 26215 -5194 26235
rect -5172 26215 -5170 26235
rect -5100 26215 -5098 26235
rect -5076 26215 -5074 26235
rect -4980 26215 -4978 26235
rect -4956 26215 -4954 26235
rect -4884 26215 -4882 26235
rect -4860 26215 -4858 26235
rect -4788 26215 -4786 26235
rect -4692 26215 -4690 26235
rect -4644 26215 -4642 26235
rect -4596 26215 -4594 26235
rect -4548 26215 -4546 26235
rect -4308 26215 -4306 26235
rect -4260 26215 -4258 26235
rect -4212 26215 -4210 26235
rect -4199 26215 -4165 26216
rect -4116 26215 -4114 26235
rect -4092 26215 -4090 26235
rect -4020 26215 -4018 26235
rect -3876 26215 -3874 26235
rect -3732 26215 -3730 26235
rect -3588 26215 -3586 26235
rect -3564 26215 -3562 26235
rect -3516 26215 -3514 26235
rect -3492 26215 -3490 26235
rect -3468 26215 -3466 26235
rect -3420 26215 -3418 26235
rect -3324 26215 -3322 26235
rect -3252 26215 -3250 26235
rect -3228 26215 -3226 26235
rect -3156 26215 -3154 26235
rect -3132 26215 -3130 26235
rect -3060 26215 -3058 26235
rect -3012 26215 -3010 26235
rect -2964 26215 -2962 26235
rect -2916 26215 -2914 26235
rect -2892 26215 -2890 26235
rect -2820 26215 -2818 26235
rect -2796 26215 -2794 26235
rect -2748 26215 -2746 26235
rect -2700 26215 -2698 26235
rect -2604 26215 -2602 26235
rect -2580 26215 -2578 26235
rect -2364 26215 -2362 26235
rect -2268 26215 -2266 26235
rect -2244 26215 -2242 26235
rect -2172 26215 -2170 26235
rect -2148 26215 -2146 26235
rect -2076 26215 -2074 26235
rect -2052 26215 -2050 26235
rect -1980 26215 -1978 26235
rect -1884 26215 -1882 26235
rect -1836 26215 -1834 26235
rect -1716 26215 -1714 26235
rect -1596 26215 -1594 26235
rect -1572 26215 -1570 26235
rect -1476 26215 -1474 26235
rect -1380 26215 -1378 26235
rect -1356 26215 -1354 26235
rect -1308 26215 -1306 26235
rect -1260 26215 -1258 26235
rect -1140 26215 -1138 26235
rect -852 26215 -850 26235
rect -804 26215 -802 26235
rect -756 26215 -754 26235
rect -708 26215 -706 26235
rect -612 26215 -610 26235
rect -588 26215 -586 26235
rect -540 26215 -538 26235
rect -492 26215 -490 26235
rect -444 26215 -442 26235
rect -396 26215 -394 26235
rect -300 26215 -298 26235
rect -276 26215 -274 26235
rect -204 26216 -202 26235
rect -239 26215 -181 26216
rect -108 26215 -106 26235
rect 12 26215 14 26235
rect 108 26215 110 26235
rect 156 26215 158 26235
rect 204 26215 206 26235
rect 228 26215 230 26235
rect 252 26215 254 26235
rect 348 26215 350 26235
rect 468 26215 470 26235
rect 492 26215 494 26235
rect 564 26215 566 26235
rect 588 26215 590 26235
rect 636 26215 638 26235
rect 660 26215 662 26235
rect 732 26215 734 26235
rect 756 26215 758 26235
rect 876 26215 878 26235
rect 972 26215 974 26235
rect 1020 26215 1022 26235
rect 1068 26215 1070 26235
rect 1092 26215 1094 26235
rect 1116 26215 1118 26235
rect 1164 26215 1166 26235
rect 1212 26215 1214 26235
rect 1308 26215 1310 26235
rect 1332 26215 1334 26235
rect 1380 26215 1382 26235
rect 1428 26215 1430 26235
rect 1524 26215 1526 26235
rect 1548 26215 1550 26235
rect 1596 26215 1598 26235
rect 1620 26215 1622 26235
rect 1644 26215 1646 26235
rect 1692 26215 1694 26235
rect 1716 26215 1718 26235
rect 1740 26215 1742 26235
rect 1788 26215 1790 26235
rect 1884 26215 1886 26235
rect 1980 26215 1982 26235
rect 2028 26215 2030 26235
rect 2076 26215 2078 26235
rect 2100 26215 2102 26235
rect 2124 26215 2126 26235
rect 2172 26215 2174 26235
rect 2196 26215 2198 26235
rect 2220 26215 2222 26235
rect 2268 26215 2270 26235
rect 2292 26215 2294 26235
rect 2316 26215 2318 26235
rect 2364 26215 2366 26235
rect 2412 26215 2414 26235
rect 2460 26215 2462 26235
rect 2508 26215 2510 26235
rect 2556 26215 2558 26235
rect 2580 26215 2582 26235
rect 2604 26215 2606 26235
rect 2652 26215 2654 26235
rect 2676 26215 2678 26235
rect 2700 26215 2702 26235
rect 2748 26215 2750 26235
rect 2772 26215 2774 26235
rect 2796 26215 2798 26235
rect 2844 26215 2846 26235
rect 2868 26215 2870 26235
rect 2892 26215 2894 26235
rect 2940 26215 2942 26235
rect 3012 26215 3014 26235
rect 3108 26215 3110 26235
rect 3156 26215 3158 26235
rect 3252 26215 3254 26235
rect 3348 26215 3350 26235
rect 3396 26215 3398 26235
rect 3468 26215 3470 26235
rect 3492 26215 3494 26235
rect 3588 26215 3590 26235
rect 3612 26215 3614 26235
rect 3636 26215 3638 26235
rect 3708 26215 3710 26235
rect 3732 26215 3734 26235
rect 3804 26215 3806 26235
rect 3828 26215 3830 26235
rect 3924 26215 3926 26235
rect 4020 26215 4022 26235
rect 4044 26215 4046 26235
rect 4092 26215 4094 26235
rect 4116 26215 4118 26235
rect 4140 26215 4142 26235
rect 4188 26215 4190 26235
rect 4212 26215 4214 26235
rect 4236 26215 4238 26235
rect 4308 26215 4310 26235
rect 4332 26215 4334 26235
rect 4404 26215 4406 26235
rect 4500 26215 4502 26235
rect 4596 26215 4598 26235
rect 4860 26215 4862 26235
rect 4956 26215 4958 26235
rect 4980 26215 4982 26235
rect 5004 26215 5006 26235
rect 5076 26215 5078 26235
rect 5100 26215 5102 26235
rect 5124 26215 5126 26235
rect 5172 26215 5174 26235
rect 5196 26216 5198 26235
rect 5185 26215 5219 26216
rect 5220 26215 5222 26235
rect 5268 26215 5270 26235
rect 5292 26215 5294 26235
rect 5388 26215 5390 26235
rect 5484 26215 5486 26235
rect 5508 26215 5510 26235
rect 5532 26215 5534 26235
rect 5628 26215 5630 26235
rect 5652 26215 5654 26235
rect 5748 26215 5750 26235
rect 5796 26215 5798 26235
rect 5844 26215 5846 26235
rect 5892 26215 5894 26235
rect 6132 26215 6134 26235
rect 6180 26215 6182 26235
rect 6228 26215 6230 26235
rect 6252 26215 6254 26235
rect 6276 26215 6278 26235
rect 6324 26215 6326 26235
rect 6372 26215 6374 26235
rect 6492 26215 6494 26235
rect 6588 26215 6590 26235
rect 6612 26215 6614 26235
rect 6660 26215 6662 26235
rect 6684 26215 6686 26235
rect 6708 26215 6710 26235
rect 6780 26215 6782 26235
rect 6804 26215 6806 26235
rect 6828 26215 6830 26235
rect 6900 26215 6902 26235
rect 6924 26215 6926 26235
rect 7020 26215 7022 26235
rect 7140 26215 7142 26235
rect 7236 26215 7238 26235
rect 7332 26215 7334 26235
rect 7380 26215 7382 26235
rect 7428 26215 7430 26235
rect 7452 26215 7454 26235
rect 7476 26215 7478 26235
rect 7524 26215 7526 26235
rect 7548 26215 7550 26235
rect 7572 26215 7574 26235
rect 7620 26215 7622 26235
rect 7644 26215 7646 26235
rect 7668 26215 7670 26235
rect 7716 26215 7718 26235
rect 7740 26215 7742 26235
rect 7836 26215 7838 26235
rect 7884 26215 7886 26235
rect 7932 26215 7934 26235
rect 7956 26215 7958 26235
rect 7980 26215 7982 26235
rect 8028 26215 8030 26235
rect 8196 26215 8198 26235
rect 8244 26215 8246 26235
rect 8268 26215 8270 26235
rect 8292 26215 8294 26235
rect 8340 26215 8342 26235
rect 8364 26215 8366 26235
rect 8388 26215 8390 26235
rect 8436 26215 8438 26235
rect 8460 26215 8462 26235
rect 8556 26215 8558 26235
rect 8604 26215 8606 26235
rect 8652 26215 8654 26235
rect 8700 26215 8702 26235
rect 8724 26215 8726 26235
rect 8748 26215 8750 26235
rect 8820 26215 8822 26235
rect 8844 26215 8846 26235
rect 8868 26215 8870 26235
rect 9516 26215 9518 26235
rect 9612 26215 9614 26235
rect 9660 26215 9662 26235
rect 9684 26215 9686 26235
rect 9708 26215 9710 26235
rect 9756 26215 9758 26235
rect 9780 26215 9782 26235
rect 9804 26215 9806 26235
rect 9852 26215 9854 26235
rect 9876 26215 9878 26235
rect 9900 26215 9902 26235
rect 9948 26215 9950 26235
rect 9972 26215 9974 26235
rect 9996 26215 9998 26235
rect 10068 26215 10070 26235
rect 10092 26215 10094 26235
rect 10116 26215 10118 26235
rect 10164 26215 10166 26235
rect 10188 26215 10190 26235
rect 10212 26215 10214 26235
rect 10284 26215 10286 26235
rect 10308 26215 10310 26235
rect 10332 26215 10334 26235
rect 10380 26215 10382 26235
rect 10404 26215 10406 26235
rect 10428 26215 10430 26235
rect 10476 26215 10478 26235
rect 10500 26215 10502 26235
rect 10524 26215 10526 26235
rect 10572 26215 10574 26235
rect 10596 26215 10598 26235
rect 10620 26215 10622 26235
rect 10668 26215 10670 26235
rect 10692 26215 10694 26235
rect 10716 26215 10718 26235
rect 10788 26215 10790 26235
rect 10836 26215 10838 26235
rect 10956 26215 10958 26235
rect 11052 26215 11054 26235
rect 11076 26215 11078 26235
rect 11124 26215 11126 26235
rect 11172 26215 11174 26235
rect 11220 26215 11222 26235
rect 11340 26215 11342 26235
rect 11436 26215 11438 26235
rect 11532 26215 11534 26235
rect 11580 26215 11582 26235
rect 11628 26215 11630 26235
rect 11676 26215 11678 26235
rect 11724 26215 11726 26235
rect 11772 26215 11774 26235
rect 11796 26215 11798 26235
rect 11892 26215 11894 26235
rect 11988 26215 11990 26235
rect 12060 26215 12062 26235
rect 12132 26215 12134 26235
rect 12228 26215 12230 26235
rect 12276 26215 12278 26235
rect 12324 26215 12326 26235
rect 12420 26215 12422 26235
rect 12444 26215 12446 26235
rect 12492 26215 12494 26235
rect 12516 26215 12518 26235
rect 12540 26215 12542 26235
rect 12588 26215 12590 26235
rect 12636 26215 12638 26235
rect 12732 26215 12734 26235
rect 12756 26215 12758 26235
rect 12804 26215 12806 26235
rect 12828 26215 12830 26235
rect 12852 26215 12854 26235
rect 12900 26215 12902 26235
rect 12948 26215 12950 26235
rect 13044 26215 13046 26235
rect 13068 26215 13070 26235
rect 13116 26215 13118 26235
rect 13284 26215 13286 26235
rect 13332 26215 13334 26235
rect 13428 26215 13430 26235
rect 13524 26215 13526 26235
rect 13572 26215 13574 26235
rect 13644 26215 13646 26235
rect 13668 26215 13670 26235
rect 13764 26215 13766 26235
rect 13812 26215 13814 26235
rect 13860 26215 13862 26235
rect 13908 26215 13910 26235
rect 13956 26215 13958 26235
rect 14004 26215 14006 26235
rect 14100 26215 14102 26235
rect 14196 26215 14198 26235
rect 14292 26215 14294 26235
rect 15132 26215 15134 26235
rect 15180 26215 15182 26235
rect 15228 26215 15230 26235
rect 15252 26215 15254 26235
rect 15324 26215 15326 26235
rect 15396 26215 15398 26235
rect 15420 26215 15422 26235
rect 15492 26215 15494 26235
rect 15540 26215 15542 26235
rect 15636 26215 15638 26235
rect 15660 26215 15662 26235
rect 15708 26215 15710 26235
rect 15732 26215 15734 26235
rect 15756 26215 15758 26235
rect 15804 26215 15806 26235
rect 15828 26215 15830 26235
rect 15852 26215 15854 26235
rect 15900 26215 15902 26235
rect 15948 26215 15950 26235
rect 15996 26215 15998 26235
rect 16044 26215 16046 26235
rect 16092 26215 16094 26235
rect 16215 26232 16229 26235
rect 16236 26232 16239 26235
rect 16260 26215 16262 26235
rect 16308 26215 16310 26235
rect 16332 26215 16334 26235
rect 16356 26215 16358 26235
rect 16404 26215 16406 26235
rect 16452 26215 16454 26235
rect 16548 26215 16550 26235
rect 16572 26215 16574 26235
rect 16620 26215 16622 26235
rect 16668 26215 16670 26235
rect 16716 26215 16718 26235
rect 16764 26215 16766 26235
rect 16836 26215 16838 26235
rect 16884 26215 16886 26235
rect 16980 26215 16982 26235
rect 17052 26215 17054 26235
rect 17196 26215 17198 26235
rect 17220 26215 17222 26235
rect 17292 26215 17294 26235
rect 17316 26215 17318 26235
rect 18084 26215 18086 26235
rect 18132 26215 18134 26235
rect 18396 26215 18398 26235
rect 18492 26215 18494 26235
rect 18516 26215 18518 26235
rect 18564 26215 18566 26235
rect 18612 26215 18614 26235
rect 18660 26215 18662 26235
rect 18708 26215 18710 26235
rect 18756 26215 18758 26235
rect 18804 26215 18806 26235
rect 18852 26215 18854 26235
rect 18900 26215 18902 26235
rect 18996 26215 18998 26235
rect 19020 26215 19022 26235
rect 19092 26215 19094 26235
rect 19116 26215 19118 26235
rect 19140 26215 19142 26235
rect 19188 26215 19190 26235
rect 19236 26215 19238 26235
rect 19332 26215 19334 26235
rect 19476 26215 19478 26235
rect 19620 26215 19622 26235
rect 19716 26215 19718 26235
rect 19788 26215 19790 26235
rect 19836 26215 19838 26235
rect 19860 26215 19862 26235
rect 19884 26215 19886 26235
rect 19932 26215 19934 26235
rect 19956 26215 19958 26235
rect 19980 26215 19982 26235
rect 20028 26215 20030 26235
rect 20052 26215 20054 26235
rect 20076 26215 20078 26235
rect 20148 26215 20150 26235
rect 20172 26215 20174 26235
rect 20196 26215 20198 26235
rect 20268 26215 20270 26235
rect 20292 26215 20294 26235
rect 20388 26215 20390 26235
rect 20412 26215 20414 26235
rect 20508 26215 20510 26235
rect 20556 26215 20558 26235
rect 20604 26215 20606 26235
rect 20916 26215 20918 26235
rect 20964 26215 20966 26235
rect 21012 26215 21014 26235
rect 21060 26215 21062 26235
rect 21084 26215 21086 26235
rect 21108 26215 21110 26235
rect 21204 26215 21206 26235
rect 21300 26215 21302 26235
rect 21324 26215 21326 26235
rect 21444 26215 21446 26235
rect 21468 26215 21470 26235
rect 21564 26215 21566 26235
rect 21612 26215 21614 26235
rect 21684 26215 21686 26235
rect 21708 26215 21710 26235
rect 21828 26215 21830 26235
rect 21924 26215 21926 26235
rect 21948 26216 21950 26235
rect 21937 26215 21971 26216
rect 22044 26215 22046 26235
rect 22068 26215 22070 26235
rect 22188 26215 22190 26235
rect 22212 26215 22214 26235
rect 23004 26215 23006 26235
rect 23052 26215 23054 26235
rect 23076 26215 23078 26235
rect 23100 26215 23102 26235
rect 23148 26215 23150 26235
rect 23220 26216 23222 26235
rect 23209 26215 23243 26216
rect 23244 26215 23246 26235
rect 23316 26215 23318 26235
rect 23340 26215 23342 26235
rect 23412 26215 23414 26235
rect 23556 26215 23558 26235
rect 23628 26215 23630 26235
rect 23652 26215 23654 26235
rect 23676 26215 23678 26235
rect 23724 26215 23726 26235
rect 23772 26215 23774 26235
rect 23820 26215 23822 26235
rect 23868 26215 23870 26235
rect 23916 26215 23918 26235
rect 24012 26215 24014 26235
rect 24084 26215 24086 26235
rect 24372 26216 24374 26235
rect 24361 26215 24395 26216
rect 24396 26215 24398 26235
rect 24492 26215 24494 26235
rect 24516 26215 24518 26235
rect 24588 26215 24590 26235
rect 24612 26215 24614 26235
rect 24708 26215 24710 26235
rect 24732 26215 24734 26235
rect 24756 26215 24758 26235
rect 24852 26215 24854 26235
rect 24876 26215 24878 26235
rect 24972 26215 24974 26235
rect 24996 26215 24998 26235
rect 25092 26215 25094 26235
rect 25260 26215 25262 26235
rect 25308 26215 25310 26235
rect 25356 26215 25358 26235
rect 25380 26215 25382 26235
rect 25404 26215 25406 26235
rect 25452 26215 25454 26235
rect 25500 26215 25502 26235
rect 25596 26215 25598 26235
rect 27060 26215 27062 26235
rect 27108 26215 27110 26235
rect 27156 26215 27158 26235
rect 27324 26215 27326 26235
rect 27396 26215 27398 26235
rect 27420 26215 27422 26235
rect 27540 26215 27542 26235
rect 27564 26215 27566 26235
rect 30564 26215 30566 26235
rect 30636 26216 30638 26235
rect 30625 26215 30659 26216
rect 30660 26215 30662 26235
rect 30780 26215 30782 26235
rect 30804 26215 30806 26235
rect 30948 26216 30950 26235
rect 30937 26215 30971 26216
rect -17385 26211 -13339 26215
rect -17385 26208 -17371 26211
rect -17292 26191 -17290 26211
rect -17207 26206 -17204 26211
rect -17196 26206 -17194 26211
rect -17197 26192 -17194 26206
rect -17028 26191 -17026 26211
rect -16932 26191 -16930 26211
rect -16860 26191 -16858 26211
rect -16836 26191 -16834 26211
rect -16764 26191 -16762 26211
rect -16740 26191 -16738 26211
rect -16668 26191 -16666 26211
rect -16500 26191 -16498 26211
rect -16380 26191 -16378 26211
rect -16356 26191 -16354 26211
rect -16284 26191 -16282 26211
rect -16260 26191 -16258 26211
rect -16236 26191 -16234 26211
rect -15300 26192 -15298 26211
rect -15335 26191 -15277 26192
rect -15084 26191 -15082 26211
rect -15057 26208 -15043 26211
rect -15036 26208 -15033 26211
rect -14868 26191 -14866 26211
rect -14772 26191 -14770 26211
rect -14724 26191 -14722 26211
rect -14508 26191 -14506 26211
rect -14436 26191 -14434 26211
rect -14340 26191 -14338 26211
rect -14244 26191 -14242 26211
rect -14172 26191 -14170 26211
rect -14076 26191 -14074 26211
rect -13980 26191 -13978 26211
rect -13932 26191 -13930 26211
rect -13884 26191 -13882 26211
rect -13716 26191 -13714 26211
rect -13644 26191 -13642 26211
rect -13596 26208 -13594 26211
rect -13596 26191 -13593 26208
rect -13500 26191 -13498 26211
rect -13356 26191 -13354 26211
rect -13353 26208 -13339 26211
rect -13329 26211 -10387 26215
rect -13329 26208 -13315 26211
rect -13284 26191 -13282 26211
rect -13068 26191 -13066 26211
rect -12828 26191 -12826 26211
rect -12780 26191 -12778 26211
rect -12660 26191 -12658 26211
rect -12564 26191 -12562 26211
rect -12492 26191 -12490 26211
rect -12396 26191 -12394 26211
rect -12348 26191 -12346 26211
rect -12276 26191 -12274 26211
rect -12252 26191 -12250 26211
rect -12156 26191 -12154 26211
rect -12060 26191 -12058 26211
rect -11892 26191 -11890 26211
rect -11844 26191 -11842 26211
rect -11796 26191 -11794 26211
rect -11676 26191 -11674 26211
rect -11580 26191 -11578 26211
rect -11556 26191 -11554 26211
rect -11508 26191 -11506 26211
rect -11460 26191 -11458 26211
rect -11436 26191 -11434 26211
rect -11364 26191 -11362 26211
rect -11340 26191 -11338 26211
rect -11268 26192 -11266 26211
rect -11303 26191 -11245 26192
rect -11172 26191 -11170 26211
rect -11124 26191 -11122 26211
rect -11076 26191 -11074 26211
rect -11028 26191 -11026 26211
rect -10788 26191 -10786 26211
rect -10668 26191 -10666 26211
rect -10401 26208 -10387 26211
rect -10377 26211 -5251 26215
rect -10377 26208 -10363 26211
rect -10007 26206 -10004 26211
rect -9876 26208 -9874 26211
rect -9997 26192 -9994 26206
rect -9996 26191 -9994 26192
rect -9876 26191 -9873 26208
rect -9708 26191 -9706 26211
rect -9612 26191 -9610 26211
rect -9516 26191 -9514 26211
rect -9468 26191 -9466 26211
rect -9420 26191 -9418 26211
rect -9396 26191 -9394 26211
rect -9372 26191 -9370 26211
rect -9300 26191 -9298 26211
rect -9252 26191 -9250 26211
rect -9132 26191 -9130 26211
rect -9084 26191 -9082 26211
rect -9036 26191 -9034 26211
rect -8988 26191 -8986 26211
rect -8940 26191 -8938 26211
rect -8892 26191 -8890 26211
rect -8855 26206 -8852 26211
rect -8844 26206 -8842 26211
rect -8845 26192 -8842 26206
rect -8772 26191 -8769 26208
rect -8604 26191 -8602 26211
rect -8508 26191 -8506 26211
rect -8484 26191 -8482 26211
rect -8388 26191 -8386 26211
rect -8364 26191 -8362 26211
rect -8340 26191 -8338 26211
rect -8268 26191 -8266 26211
rect -8100 26191 -8098 26211
rect -8052 26191 -8050 26211
rect -7932 26191 -7930 26211
rect -7692 26191 -7690 26211
rect -7620 26191 -7618 26211
rect -7404 26191 -7402 26211
rect -7356 26191 -7354 26211
rect -7308 26191 -7306 26211
rect -7212 26191 -7210 26211
rect -7188 26191 -7186 26211
rect -7116 26191 -7114 26211
rect -7068 26191 -7066 26211
rect -6972 26191 -6970 26211
rect -6948 26191 -6946 26211
rect -6876 26191 -6874 26211
rect -6852 26191 -6850 26211
rect -6780 26191 -6778 26211
rect -6756 26191 -6754 26211
rect -6660 26191 -6658 26211
rect -6612 26191 -6610 26211
rect -6564 26192 -6562 26211
rect -6575 26191 -6541 26192
rect -6516 26191 -6514 26211
rect -6492 26191 -6490 26211
rect -6468 26191 -6466 26211
rect -6420 26191 -6418 26211
rect -6396 26191 -6394 26211
rect -6372 26191 -6370 26211
rect -6324 26191 -6322 26211
rect -6300 26191 -6298 26211
rect -6276 26192 -6274 26211
rect -6228 26192 -6226 26211
rect -6287 26191 -6205 26192
rect -6180 26191 -6178 26211
rect -6060 26191 -6058 26211
rect -5940 26191 -5938 26211
rect -5892 26191 -5890 26211
rect -5652 26191 -5650 26211
rect -5268 26191 -5266 26211
rect -5265 26208 -5251 26211
rect -5241 26211 30971 26215
rect -5241 26208 -5227 26211
rect -5196 26191 -5194 26211
rect -5172 26191 -5170 26211
rect -5100 26191 -5098 26211
rect -5076 26191 -5074 26211
rect -4980 26191 -4978 26211
rect -4956 26191 -4954 26211
rect -4884 26191 -4882 26211
rect -4860 26191 -4858 26211
rect -4788 26191 -4786 26211
rect -4692 26191 -4690 26211
rect -4644 26191 -4642 26211
rect -4596 26191 -4594 26211
rect -4548 26191 -4546 26211
rect -4308 26191 -4306 26211
rect -4260 26191 -4258 26211
rect -4212 26191 -4210 26211
rect -4116 26191 -4114 26211
rect -4092 26208 -4090 26211
rect -4092 26191 -4089 26208
rect -4020 26191 -4018 26211
rect -3876 26191 -3874 26211
rect -3732 26191 -3730 26211
rect -3588 26191 -3586 26211
rect -3564 26191 -3562 26211
rect -3516 26191 -3514 26211
rect -3492 26191 -3490 26211
rect -3468 26191 -3466 26211
rect -3420 26191 -3418 26211
rect -3324 26191 -3322 26211
rect -3252 26191 -3250 26211
rect -3228 26191 -3226 26211
rect -3156 26191 -3154 26211
rect -3132 26191 -3130 26211
rect -3060 26191 -3058 26211
rect -3012 26191 -3010 26211
rect -2964 26191 -2962 26211
rect -2916 26191 -2914 26211
rect -2892 26191 -2890 26211
rect -2820 26191 -2818 26211
rect -2796 26191 -2794 26211
rect -2748 26191 -2746 26211
rect -2700 26191 -2698 26211
rect -2604 26191 -2602 26211
rect -2580 26191 -2578 26211
rect -2364 26191 -2362 26211
rect -2268 26191 -2266 26211
rect -2244 26191 -2242 26211
rect -2172 26191 -2170 26211
rect -2148 26191 -2146 26211
rect -2076 26191 -2074 26211
rect -2052 26191 -2050 26211
rect -1980 26191 -1978 26211
rect -1884 26191 -1882 26211
rect -1836 26191 -1834 26211
rect -1716 26191 -1714 26211
rect -1596 26191 -1594 26211
rect -1572 26191 -1570 26211
rect -1476 26191 -1474 26211
rect -1380 26191 -1378 26211
rect -1356 26191 -1354 26211
rect -1308 26191 -1306 26211
rect -1260 26191 -1258 26211
rect -1140 26191 -1138 26211
rect -852 26191 -850 26211
rect -804 26191 -802 26211
rect -756 26191 -754 26211
rect -708 26191 -706 26211
rect -612 26191 -610 26211
rect -588 26191 -586 26211
rect -540 26191 -538 26211
rect -492 26191 -490 26211
rect -444 26191 -442 26211
rect -396 26191 -394 26211
rect -300 26191 -298 26211
rect -276 26191 -274 26211
rect -239 26206 -236 26211
rect -215 26206 -212 26211
rect -204 26206 -202 26211
rect -229 26192 -226 26206
rect -205 26192 -202 26206
rect -108 26208 -106 26211
rect -228 26191 -226 26192
rect -108 26191 -105 26208
rect 12 26191 14 26211
rect 108 26191 110 26211
rect 156 26191 158 26211
rect 204 26191 206 26211
rect 228 26191 230 26211
rect 252 26191 254 26211
rect 348 26191 350 26211
rect 468 26191 470 26211
rect 492 26191 494 26211
rect 564 26191 566 26211
rect 588 26191 590 26211
rect 636 26191 638 26211
rect 660 26191 662 26211
rect 732 26191 734 26211
rect 756 26191 758 26211
rect 876 26191 878 26211
rect 972 26191 974 26211
rect 1020 26191 1022 26211
rect 1068 26191 1070 26211
rect 1092 26191 1094 26211
rect 1116 26191 1118 26211
rect 1164 26191 1166 26211
rect 1212 26191 1214 26211
rect 1308 26191 1310 26211
rect 1332 26191 1334 26211
rect 1380 26191 1382 26211
rect 1428 26191 1430 26211
rect 1524 26191 1526 26211
rect 1548 26191 1550 26211
rect 1596 26191 1598 26211
rect 1620 26191 1622 26211
rect 1644 26191 1646 26211
rect 1692 26191 1694 26211
rect 1716 26191 1718 26211
rect 1740 26191 1742 26211
rect 1788 26191 1790 26211
rect 1884 26191 1886 26211
rect 1980 26191 1982 26211
rect 2028 26191 2030 26211
rect 2076 26191 2078 26211
rect 2100 26191 2102 26211
rect 2124 26191 2126 26211
rect 2172 26191 2174 26211
rect 2196 26191 2198 26211
rect 2220 26191 2222 26211
rect 2268 26191 2270 26211
rect 2292 26191 2294 26211
rect 2316 26191 2318 26211
rect 2364 26191 2366 26211
rect 2412 26191 2414 26211
rect 2460 26191 2462 26211
rect 2508 26191 2510 26211
rect 2556 26191 2558 26211
rect 2580 26191 2582 26211
rect 2604 26191 2606 26211
rect 2652 26191 2654 26211
rect 2676 26191 2678 26211
rect 2700 26191 2702 26211
rect 2748 26191 2750 26211
rect 2772 26191 2774 26211
rect 2796 26191 2798 26211
rect 2844 26191 2846 26211
rect 2868 26191 2870 26211
rect 2892 26191 2894 26211
rect 2940 26191 2942 26211
rect 3012 26191 3014 26211
rect 3108 26191 3110 26211
rect 3156 26191 3158 26211
rect 3252 26191 3254 26211
rect 3348 26191 3350 26211
rect 3396 26191 3398 26211
rect 3468 26191 3470 26211
rect 3492 26191 3494 26211
rect 3588 26191 3590 26211
rect 3612 26191 3614 26211
rect 3636 26191 3638 26211
rect 3708 26191 3710 26211
rect 3732 26191 3734 26211
rect 3804 26191 3806 26211
rect 3828 26191 3830 26211
rect 3924 26191 3926 26211
rect 4020 26191 4022 26211
rect 4044 26191 4046 26211
rect 4092 26191 4094 26211
rect 4116 26191 4118 26211
rect 4140 26191 4142 26211
rect 4188 26191 4190 26211
rect 4212 26191 4214 26211
rect 4236 26191 4238 26211
rect 4308 26191 4310 26211
rect 4332 26191 4334 26211
rect 4404 26191 4406 26211
rect 4500 26191 4502 26211
rect 4596 26191 4598 26211
rect 4860 26191 4862 26211
rect 4956 26191 4958 26211
rect 4980 26191 4982 26211
rect 5004 26191 5006 26211
rect 5076 26191 5078 26211
rect 5100 26191 5102 26211
rect 5124 26191 5126 26211
rect 5172 26191 5174 26211
rect 5185 26206 5188 26211
rect 5196 26206 5198 26211
rect 5195 26192 5198 26206
rect 5220 26191 5222 26211
rect 5268 26191 5270 26211
rect 5292 26208 5294 26211
rect 5292 26191 5295 26208
rect 5388 26191 5390 26211
rect 5484 26191 5486 26211
rect 5508 26191 5510 26211
rect 5532 26191 5534 26211
rect 5628 26191 5630 26211
rect 5652 26191 5654 26211
rect 5748 26191 5750 26211
rect 5796 26191 5798 26211
rect 5844 26191 5846 26211
rect 5892 26191 5894 26211
rect 6132 26191 6134 26211
rect 6180 26191 6182 26211
rect 6228 26191 6230 26211
rect 6252 26191 6254 26211
rect 6276 26191 6278 26211
rect 6324 26191 6326 26211
rect 6372 26191 6374 26211
rect 6492 26191 6494 26211
rect 6588 26191 6590 26211
rect 6612 26191 6614 26211
rect 6660 26191 6662 26211
rect 6684 26191 6686 26211
rect 6708 26191 6710 26211
rect 6780 26191 6782 26211
rect 6804 26191 6806 26211
rect 6828 26191 6830 26211
rect 6900 26191 6902 26211
rect 6924 26191 6926 26211
rect 7020 26191 7022 26211
rect 7140 26191 7142 26211
rect 7236 26191 7238 26211
rect 7332 26191 7334 26211
rect 7380 26191 7382 26211
rect 7428 26191 7430 26211
rect 7452 26191 7454 26211
rect 7476 26191 7478 26211
rect 7524 26191 7526 26211
rect 7548 26191 7550 26211
rect 7572 26191 7574 26211
rect 7620 26191 7622 26211
rect 7644 26191 7646 26211
rect 7668 26191 7670 26211
rect 7716 26191 7718 26211
rect 7740 26191 7742 26211
rect 7836 26191 7838 26211
rect 7884 26191 7886 26211
rect 7932 26191 7934 26211
rect 7956 26191 7958 26211
rect 7980 26191 7982 26211
rect 8028 26191 8030 26211
rect 8196 26191 8198 26211
rect 8244 26191 8246 26211
rect 8268 26191 8270 26211
rect 8292 26191 8294 26211
rect 8340 26191 8342 26211
rect 8364 26191 8366 26211
rect 8388 26191 8390 26211
rect 8436 26191 8438 26211
rect 8460 26191 8462 26211
rect 8556 26191 8558 26211
rect 8604 26191 8606 26211
rect 8652 26191 8654 26211
rect 8700 26191 8702 26211
rect 8724 26191 8726 26211
rect 8748 26191 8750 26211
rect 8820 26191 8822 26211
rect 8844 26191 8846 26211
rect 8868 26191 8870 26211
rect 9516 26191 9518 26211
rect 9612 26191 9614 26211
rect 9660 26191 9662 26211
rect 9684 26191 9686 26211
rect 9708 26191 9710 26211
rect 9756 26191 9758 26211
rect 9780 26191 9782 26211
rect 9804 26191 9806 26211
rect 9852 26191 9854 26211
rect 9876 26191 9878 26211
rect 9900 26191 9902 26211
rect 9948 26191 9950 26211
rect 9972 26191 9974 26211
rect 9996 26191 9998 26211
rect 10068 26191 10070 26211
rect 10092 26191 10094 26211
rect 10116 26191 10118 26211
rect 10164 26191 10166 26211
rect 10188 26191 10190 26211
rect 10212 26191 10214 26211
rect 10284 26191 10286 26211
rect 10308 26191 10310 26211
rect 10332 26191 10334 26211
rect 10380 26191 10382 26211
rect 10404 26191 10406 26211
rect 10428 26191 10430 26211
rect 10476 26191 10478 26211
rect 10500 26191 10502 26211
rect 10524 26191 10526 26211
rect 10572 26191 10574 26211
rect 10596 26191 10598 26211
rect 10620 26191 10622 26211
rect 10668 26191 10670 26211
rect 10692 26191 10694 26211
rect 10716 26191 10718 26211
rect 10788 26191 10790 26211
rect 10836 26191 10838 26211
rect 10956 26191 10958 26211
rect 11052 26191 11054 26211
rect 11076 26191 11078 26211
rect 11124 26191 11126 26211
rect 11172 26191 11174 26211
rect 11220 26191 11222 26211
rect 11340 26191 11342 26211
rect 11436 26191 11438 26211
rect 11532 26191 11534 26211
rect 11580 26191 11582 26211
rect 11628 26191 11630 26211
rect 11676 26191 11678 26211
rect 11724 26191 11726 26211
rect 11772 26191 11774 26211
rect 11796 26191 11798 26211
rect 11892 26191 11894 26211
rect 11988 26191 11990 26211
rect 12060 26191 12062 26211
rect 12132 26191 12134 26211
rect 12228 26191 12230 26211
rect 12276 26191 12278 26211
rect 12324 26191 12326 26211
rect 12420 26191 12422 26211
rect 12444 26191 12446 26211
rect 12492 26191 12494 26211
rect 12516 26191 12518 26211
rect 12540 26191 12542 26211
rect 12588 26191 12590 26211
rect 12636 26191 12638 26211
rect 12732 26191 12734 26211
rect 12756 26191 12758 26211
rect 12804 26191 12806 26211
rect 12828 26191 12830 26211
rect 12852 26191 12854 26211
rect 12900 26191 12902 26211
rect 12948 26191 12950 26211
rect 13044 26191 13046 26211
rect 13068 26191 13070 26211
rect 13116 26191 13118 26211
rect 13284 26191 13286 26211
rect 13332 26191 13334 26211
rect 13428 26191 13430 26211
rect 13524 26191 13526 26211
rect 13572 26191 13574 26211
rect 13644 26191 13646 26211
rect 13668 26191 13670 26211
rect 13764 26191 13766 26211
rect 13812 26191 13814 26211
rect 13860 26191 13862 26211
rect 13908 26191 13910 26211
rect 13956 26191 13958 26211
rect 14004 26191 14006 26211
rect 14100 26191 14102 26211
rect 14196 26191 14198 26211
rect 14292 26191 14294 26211
rect 15132 26191 15134 26211
rect 15180 26191 15182 26211
rect 15228 26191 15230 26211
rect 15252 26191 15254 26211
rect 15324 26191 15326 26211
rect 15396 26191 15398 26211
rect 15420 26191 15422 26211
rect 15492 26191 15494 26211
rect 15540 26191 15542 26211
rect 15636 26191 15638 26211
rect 15660 26191 15662 26211
rect 15708 26191 15710 26211
rect 15732 26191 15734 26211
rect 15756 26191 15758 26211
rect 15804 26191 15806 26211
rect 15828 26191 15830 26211
rect 15852 26191 15854 26211
rect 15900 26191 15902 26211
rect 15948 26191 15950 26211
rect 15996 26191 15998 26211
rect 16044 26191 16046 26211
rect 16092 26191 16094 26211
rect 16260 26191 16262 26211
rect 16308 26191 16310 26211
rect 16332 26191 16334 26211
rect 16356 26191 16358 26211
rect 16404 26191 16406 26211
rect 16452 26191 16454 26211
rect 16548 26191 16550 26211
rect 16572 26191 16574 26211
rect 16620 26191 16622 26211
rect 16668 26191 16670 26211
rect 16716 26191 16718 26211
rect 16764 26191 16766 26211
rect 16836 26192 16838 26211
rect 16801 26191 16859 26192
rect 16884 26191 16886 26211
rect 16980 26191 16982 26211
rect 17052 26191 17054 26211
rect 17196 26191 17198 26211
rect 17220 26191 17222 26211
rect 17292 26191 17294 26211
rect 17316 26191 17318 26211
rect 18084 26191 18086 26211
rect 18132 26191 18134 26211
rect 18396 26191 18398 26211
rect 18492 26191 18494 26211
rect 18516 26191 18518 26211
rect 18564 26191 18566 26211
rect 18612 26191 18614 26211
rect 18660 26191 18662 26211
rect 18708 26191 18710 26211
rect 18756 26191 18758 26211
rect 18804 26191 18806 26211
rect 18852 26191 18854 26211
rect 18900 26191 18902 26211
rect 18996 26191 18998 26211
rect 19020 26191 19022 26211
rect 19092 26191 19094 26211
rect 19116 26191 19118 26211
rect 19140 26191 19142 26211
rect 19188 26191 19190 26211
rect 19236 26191 19238 26211
rect 19332 26191 19334 26211
rect 19476 26191 19478 26211
rect 19620 26191 19622 26211
rect 19716 26191 19718 26211
rect 19788 26191 19790 26211
rect 19836 26191 19838 26211
rect 19860 26191 19862 26211
rect 19884 26191 19886 26211
rect 19932 26191 19934 26211
rect 19956 26191 19958 26211
rect 19980 26191 19982 26211
rect 20028 26191 20030 26211
rect 20052 26191 20054 26211
rect 20076 26191 20078 26211
rect 20148 26191 20150 26211
rect 20172 26191 20174 26211
rect 20196 26191 20198 26211
rect 20268 26191 20270 26211
rect 20292 26191 20294 26211
rect 20388 26191 20390 26211
rect 20412 26191 20414 26211
rect 20508 26191 20510 26211
rect 20556 26191 20558 26211
rect 20604 26191 20606 26211
rect 20916 26191 20918 26211
rect 20964 26191 20966 26211
rect 21012 26191 21014 26211
rect 21060 26191 21062 26211
rect 21084 26191 21086 26211
rect 21108 26191 21110 26211
rect 21204 26191 21206 26211
rect 21300 26191 21302 26211
rect 21324 26191 21326 26211
rect 21444 26191 21446 26211
rect 21468 26191 21470 26211
rect 21564 26191 21566 26211
rect 21612 26191 21614 26211
rect 21684 26191 21686 26211
rect 21708 26191 21710 26211
rect 21828 26191 21830 26211
rect 21924 26191 21926 26211
rect 21937 26206 21940 26211
rect 21948 26206 21950 26211
rect 21947 26192 21950 26206
rect 22044 26208 22046 26211
rect 22044 26191 22047 26208
rect 22068 26191 22070 26211
rect 22188 26191 22190 26211
rect 22212 26191 22214 26211
rect 22873 26191 22931 26192
rect 23004 26191 23006 26211
rect 23052 26191 23054 26211
rect 23076 26191 23078 26211
rect 23100 26191 23102 26211
rect 23148 26191 23150 26211
rect 23209 26206 23212 26211
rect 23220 26206 23222 26211
rect 23219 26192 23222 26206
rect 23244 26191 23246 26211
rect 23316 26208 23318 26211
rect 23316 26191 23319 26208
rect 23340 26191 23342 26211
rect 23412 26191 23414 26211
rect 23556 26191 23558 26211
rect 23628 26191 23630 26211
rect 23652 26191 23654 26211
rect 23676 26191 23678 26211
rect 23724 26191 23726 26211
rect 23772 26191 23774 26211
rect 23820 26191 23822 26211
rect 23868 26191 23870 26211
rect 23916 26191 23918 26211
rect 24012 26191 24014 26211
rect 24084 26191 24086 26211
rect 24361 26206 24364 26211
rect 24372 26206 24374 26211
rect 24371 26192 24374 26206
rect 24396 26191 24398 26211
rect 24492 26191 24494 26211
rect 24516 26191 24518 26211
rect 24588 26191 24590 26211
rect 24612 26191 24614 26211
rect 24708 26191 24710 26211
rect 24732 26191 24734 26211
rect 24756 26191 24758 26211
rect 24852 26191 24854 26211
rect 24876 26191 24878 26211
rect 24972 26191 24974 26211
rect 24996 26191 24998 26211
rect 25092 26191 25094 26211
rect 25260 26191 25262 26211
rect 25308 26191 25310 26211
rect 25356 26191 25358 26211
rect 25380 26191 25382 26211
rect 25404 26191 25406 26211
rect 25452 26191 25454 26211
rect 25500 26191 25502 26211
rect 25596 26191 25598 26211
rect 27060 26192 27062 26211
rect 27025 26191 27083 26192
rect 27108 26191 27110 26211
rect 27156 26191 27158 26211
rect 27324 26191 27326 26211
rect 27396 26191 27398 26211
rect 27420 26191 27422 26211
rect 27540 26191 27542 26211
rect 27564 26191 27566 26211
rect 30564 26191 30566 26211
rect 30625 26206 30628 26211
rect 30636 26206 30638 26211
rect 30635 26192 30638 26206
rect 30660 26191 30662 26211
rect 30780 26191 30782 26211
rect 30804 26191 30806 26211
rect 30937 26206 30940 26211
rect 30948 26206 30950 26211
rect 30947 26192 30950 26206
rect 30913 26191 30947 26192
rect -17855 26187 -9907 26191
rect -17855 26184 -17851 26187
rect -17844 26184 -17841 26187
rect -17735 26167 -17701 26168
rect -17508 26167 -17506 26187
rect -17484 26167 -17482 26187
rect -17471 26167 -17413 26168
rect -17388 26167 -17386 26187
rect -17292 26167 -17290 26187
rect -17121 26184 -17107 26187
rect -17028 26167 -17026 26187
rect -16932 26167 -16930 26187
rect -16860 26167 -16858 26187
rect -16836 26167 -16834 26187
rect -16764 26167 -16762 26187
rect -16740 26167 -16738 26187
rect -16668 26167 -16666 26187
rect -16500 26167 -16498 26187
rect -16380 26168 -16378 26187
rect -16391 26167 -16357 26168
rect -17735 26163 -16357 26167
rect -17615 26143 -17581 26144
rect -17508 26143 -17506 26163
rect -17484 26143 -17482 26163
rect -17471 26158 -17468 26163
rect -17461 26144 -17458 26158
rect -17460 26143 -17458 26144
rect -17388 26143 -17386 26163
rect -17292 26143 -17290 26163
rect -17028 26143 -17026 26163
rect -16967 26143 -16933 26144
rect -16932 26143 -16930 26163
rect -16860 26143 -16858 26163
rect -16836 26143 -16834 26163
rect -16764 26143 -16762 26163
rect -16740 26143 -16738 26163
rect -16668 26143 -16666 26163
rect -16631 26143 -16573 26144
rect -16500 26143 -16498 26163
rect -16391 26158 -16388 26163
rect -16380 26158 -16378 26163
rect -16381 26144 -16378 26158
rect -16380 26143 -16378 26144
rect -16356 26143 -16354 26187
rect -16319 26167 -16285 26168
rect -16284 26167 -16282 26187
rect -16260 26167 -16258 26187
rect -16236 26167 -16234 26187
rect -15335 26182 -15332 26187
rect -15311 26182 -15308 26187
rect -15300 26182 -15298 26187
rect -15325 26168 -15322 26182
rect -15301 26168 -15298 26182
rect -15324 26167 -15322 26168
rect -15084 26167 -15082 26187
rect -14961 26184 -14947 26187
rect -14868 26167 -14866 26187
rect -14772 26167 -14770 26187
rect -14724 26167 -14722 26187
rect -14508 26167 -14506 26187
rect -14436 26167 -14434 26187
rect -14340 26167 -14338 26187
rect -14244 26167 -14242 26187
rect -14172 26167 -14170 26187
rect -14076 26167 -14074 26187
rect -13980 26167 -13978 26187
rect -13932 26167 -13930 26187
rect -13884 26167 -13882 26187
rect -13716 26167 -13714 26187
rect -13644 26167 -13642 26187
rect -13617 26184 -13603 26187
rect -13596 26184 -13593 26187
rect -13500 26167 -13498 26187
rect -13356 26167 -13354 26187
rect -13284 26167 -13282 26187
rect -13068 26167 -13066 26187
rect -12828 26167 -12826 26187
rect -12780 26167 -12778 26187
rect -12660 26167 -12658 26187
rect -12564 26167 -12562 26187
rect -12492 26167 -12490 26187
rect -12396 26167 -12394 26187
rect -12348 26167 -12346 26187
rect -12276 26167 -12274 26187
rect -12252 26167 -12250 26187
rect -12156 26167 -12154 26187
rect -12060 26167 -12058 26187
rect -11927 26167 -11893 26168
rect -11892 26167 -11890 26187
rect -11844 26167 -11842 26187
rect -11796 26167 -11794 26187
rect -11676 26167 -11674 26187
rect -11580 26167 -11578 26187
rect -11556 26167 -11554 26187
rect -11508 26167 -11506 26187
rect -11460 26167 -11458 26187
rect -11436 26167 -11434 26187
rect -11364 26167 -11362 26187
rect -11340 26167 -11338 26187
rect -11303 26182 -11300 26187
rect -11279 26182 -11276 26187
rect -11268 26182 -11266 26187
rect -11293 26168 -11290 26182
rect -11269 26168 -11266 26182
rect -11172 26184 -11170 26187
rect -11292 26167 -11290 26168
rect -11172 26167 -11169 26184
rect -11124 26167 -11122 26187
rect -11076 26167 -11074 26187
rect -11028 26167 -11026 26187
rect -10788 26167 -10786 26187
rect -10751 26167 -10693 26168
rect -10668 26167 -10666 26187
rect -9996 26167 -9994 26187
rect -9921 26184 -9907 26187
rect -9897 26187 -8779 26191
rect -9897 26184 -9883 26187
rect -9876 26184 -9873 26187
rect -9708 26167 -9706 26187
rect -9612 26167 -9610 26187
rect -9516 26167 -9514 26187
rect -9468 26167 -9466 26187
rect -9420 26167 -9418 26187
rect -9396 26167 -9394 26187
rect -9372 26167 -9370 26187
rect -9300 26167 -9298 26187
rect -9252 26167 -9250 26187
rect -9132 26167 -9130 26187
rect -9084 26167 -9082 26187
rect -9036 26167 -9034 26187
rect -8988 26167 -8986 26187
rect -8940 26167 -8938 26187
rect -8892 26167 -8890 26187
rect -8793 26184 -8779 26187
rect -8772 26187 -139 26191
rect -8772 26184 -8755 26187
rect -8772 26167 -8770 26184
rect -8604 26167 -8602 26187
rect -8508 26167 -8506 26187
rect -8484 26167 -8482 26187
rect -8388 26167 -8386 26187
rect -8364 26167 -8362 26187
rect -8340 26167 -8338 26187
rect -8268 26167 -8266 26187
rect -8100 26167 -8098 26187
rect -8052 26167 -8050 26187
rect -7932 26167 -7930 26187
rect -7692 26167 -7690 26187
rect -7620 26167 -7618 26187
rect -7535 26167 -7477 26168
rect -7404 26167 -7402 26187
rect -7356 26167 -7354 26187
rect -7308 26167 -7306 26187
rect -7212 26167 -7210 26187
rect -7188 26167 -7186 26187
rect -7116 26167 -7114 26187
rect -7068 26167 -7066 26187
rect -6972 26167 -6970 26187
rect -6948 26167 -6946 26187
rect -6876 26167 -6874 26187
rect -6852 26167 -6850 26187
rect -6780 26167 -6778 26187
rect -6756 26167 -6754 26187
rect -6660 26167 -6658 26187
rect -6612 26167 -6610 26187
rect -6575 26182 -6572 26187
rect -6564 26182 -6562 26187
rect -6565 26168 -6562 26182
rect -6516 26167 -6514 26187
rect -6492 26167 -6490 26187
rect -6468 26184 -6466 26187
rect -6468 26167 -6465 26184
rect -6420 26167 -6418 26187
rect -6396 26167 -6394 26187
rect -6372 26167 -6370 26187
rect -6324 26167 -6322 26187
rect -6300 26167 -6298 26187
rect -6287 26182 -6284 26187
rect -6276 26182 -6274 26187
rect -6239 26182 -6236 26187
rect -6228 26182 -6226 26187
rect -6277 26168 -6274 26182
rect -6229 26168 -6226 26182
rect -6180 26184 -6178 26187
rect -6180 26167 -6177 26184
rect -6156 26167 -6153 26184
rect -6060 26167 -6058 26187
rect -5940 26167 -5938 26187
rect -5892 26167 -5890 26187
rect -5652 26167 -5650 26187
rect -5268 26167 -5266 26187
rect -5196 26167 -5194 26187
rect -5172 26167 -5170 26187
rect -5100 26167 -5098 26187
rect -5076 26167 -5074 26187
rect -4980 26167 -4978 26187
rect -4956 26167 -4954 26187
rect -4884 26167 -4882 26187
rect -4860 26167 -4858 26187
rect -4788 26167 -4786 26187
rect -4692 26167 -4690 26187
rect -4644 26167 -4642 26187
rect -4596 26167 -4594 26187
rect -4548 26167 -4546 26187
rect -4308 26167 -4306 26187
rect -4260 26167 -4258 26187
rect -4212 26167 -4210 26187
rect -4175 26167 -4117 26168
rect -4116 26167 -4114 26187
rect -4113 26184 -4099 26187
rect -4092 26184 -4089 26187
rect -4020 26167 -4018 26187
rect -3876 26167 -3874 26187
rect -3732 26167 -3730 26187
rect -3588 26167 -3586 26187
rect -3564 26167 -3562 26187
rect -3516 26167 -3514 26187
rect -3492 26167 -3490 26187
rect -3468 26167 -3466 26187
rect -3420 26167 -3418 26187
rect -3324 26167 -3322 26187
rect -3252 26167 -3250 26187
rect -3228 26167 -3226 26187
rect -3156 26167 -3154 26187
rect -3132 26167 -3130 26187
rect -3060 26167 -3058 26187
rect -3012 26167 -3010 26187
rect -2964 26167 -2962 26187
rect -2916 26167 -2914 26187
rect -2892 26167 -2890 26187
rect -2820 26167 -2818 26187
rect -2796 26167 -2794 26187
rect -2748 26167 -2746 26187
rect -2700 26167 -2698 26187
rect -2604 26167 -2602 26187
rect -2580 26167 -2578 26187
rect -2364 26167 -2362 26187
rect -2268 26167 -2266 26187
rect -2244 26167 -2242 26187
rect -2172 26167 -2170 26187
rect -2148 26167 -2146 26187
rect -2076 26167 -2074 26187
rect -2052 26167 -2050 26187
rect -1980 26167 -1978 26187
rect -1884 26167 -1882 26187
rect -1836 26167 -1834 26187
rect -1716 26167 -1714 26187
rect -1596 26167 -1594 26187
rect -1572 26167 -1570 26187
rect -1476 26167 -1474 26187
rect -1380 26167 -1378 26187
rect -1356 26167 -1354 26187
rect -1308 26167 -1306 26187
rect -1260 26167 -1258 26187
rect -1140 26167 -1138 26187
rect -852 26167 -850 26187
rect -804 26167 -802 26187
rect -756 26167 -754 26187
rect -708 26167 -706 26187
rect -612 26167 -610 26187
rect -588 26167 -586 26187
rect -540 26167 -538 26187
rect -492 26167 -490 26187
rect -444 26167 -442 26187
rect -396 26167 -394 26187
rect -300 26167 -298 26187
rect -276 26167 -274 26187
rect -228 26167 -226 26187
rect -153 26184 -139 26187
rect -129 26187 30947 26191
rect -129 26184 -115 26187
rect -108 26184 -105 26187
rect 12 26167 14 26187
rect 108 26167 110 26187
rect 156 26167 158 26187
rect 204 26167 206 26187
rect 228 26167 230 26187
rect 252 26167 254 26187
rect 348 26167 350 26187
rect 468 26167 470 26187
rect 492 26167 494 26187
rect 564 26167 566 26187
rect 588 26167 590 26187
rect 636 26167 638 26187
rect 660 26167 662 26187
rect 732 26167 734 26187
rect 756 26167 758 26187
rect 876 26167 878 26187
rect 972 26167 974 26187
rect 1020 26167 1022 26187
rect 1068 26167 1070 26187
rect 1092 26167 1094 26187
rect 1116 26167 1118 26187
rect 1164 26167 1166 26187
rect 1212 26167 1214 26187
rect 1308 26167 1310 26187
rect 1332 26167 1334 26187
rect 1380 26167 1382 26187
rect 1428 26167 1430 26187
rect 1524 26167 1526 26187
rect 1548 26167 1550 26187
rect 1596 26167 1598 26187
rect 1620 26167 1622 26187
rect 1644 26167 1646 26187
rect 1692 26167 1694 26187
rect 1716 26167 1718 26187
rect 1740 26167 1742 26187
rect 1788 26167 1790 26187
rect 1884 26167 1886 26187
rect 1980 26167 1982 26187
rect 2028 26167 2030 26187
rect 2076 26167 2078 26187
rect 2100 26167 2102 26187
rect 2124 26167 2126 26187
rect 2172 26167 2174 26187
rect 2196 26167 2198 26187
rect 2220 26167 2222 26187
rect 2268 26167 2270 26187
rect 2292 26167 2294 26187
rect 2316 26167 2318 26187
rect 2364 26167 2366 26187
rect 2412 26167 2414 26187
rect 2460 26167 2462 26187
rect 2508 26167 2510 26187
rect 2556 26168 2558 26187
rect 2521 26167 2579 26168
rect 2580 26167 2582 26187
rect 2604 26167 2606 26187
rect 2652 26167 2654 26187
rect 2676 26167 2678 26187
rect 2700 26167 2702 26187
rect 2748 26167 2750 26187
rect 2772 26167 2774 26187
rect 2796 26167 2798 26187
rect 2844 26167 2846 26187
rect 2868 26167 2870 26187
rect 2892 26167 2894 26187
rect 2940 26167 2942 26187
rect 3012 26167 3014 26187
rect 3108 26167 3110 26187
rect 3156 26167 3158 26187
rect 3252 26167 3254 26187
rect 3348 26167 3350 26187
rect 3396 26167 3398 26187
rect 3468 26167 3470 26187
rect 3492 26167 3494 26187
rect 3588 26167 3590 26187
rect 3612 26167 3614 26187
rect 3636 26167 3638 26187
rect 3708 26167 3710 26187
rect 3732 26167 3734 26187
rect 3804 26167 3806 26187
rect 3828 26167 3830 26187
rect 3924 26167 3926 26187
rect 4020 26167 4022 26187
rect 4044 26167 4046 26187
rect 4092 26167 4094 26187
rect 4116 26167 4118 26187
rect 4140 26167 4142 26187
rect 4188 26167 4190 26187
rect 4212 26167 4214 26187
rect 4236 26167 4238 26187
rect 4308 26167 4310 26187
rect 4332 26167 4334 26187
rect 4404 26167 4406 26187
rect 4500 26167 4502 26187
rect 4596 26167 4598 26187
rect 4860 26167 4862 26187
rect 4956 26167 4958 26187
rect 4980 26167 4982 26187
rect 5004 26167 5006 26187
rect 5076 26167 5078 26187
rect 5100 26167 5102 26187
rect 5124 26167 5126 26187
rect 5172 26167 5174 26187
rect 5220 26167 5222 26187
rect 5268 26167 5270 26187
rect 5271 26184 5285 26187
rect 5292 26184 5295 26187
rect 5388 26167 5390 26187
rect 5484 26167 5486 26187
rect 5508 26167 5510 26187
rect 5532 26167 5534 26187
rect 5628 26167 5630 26187
rect 5652 26167 5654 26187
rect 5748 26167 5750 26187
rect 5796 26167 5798 26187
rect 5844 26167 5846 26187
rect 5892 26167 5894 26187
rect 5953 26167 5987 26168
rect 6132 26167 6134 26187
rect 6180 26167 6182 26187
rect 6228 26167 6230 26187
rect 6252 26167 6254 26187
rect 6276 26167 6278 26187
rect 6324 26167 6326 26187
rect 6372 26167 6374 26187
rect 6492 26167 6494 26187
rect 6588 26167 6590 26187
rect 6612 26167 6614 26187
rect 6660 26167 6662 26187
rect 6684 26167 6686 26187
rect 6708 26167 6710 26187
rect 6780 26167 6782 26187
rect 6804 26167 6806 26187
rect 6828 26167 6830 26187
rect 6900 26167 6902 26187
rect 6924 26167 6926 26187
rect 7020 26167 7022 26187
rect 7140 26167 7142 26187
rect 7236 26167 7238 26187
rect 7332 26167 7334 26187
rect 7380 26167 7382 26187
rect 7428 26167 7430 26187
rect 7452 26167 7454 26187
rect 7476 26167 7478 26187
rect 7524 26167 7526 26187
rect 7548 26167 7550 26187
rect 7572 26167 7574 26187
rect 7620 26167 7622 26187
rect 7644 26167 7646 26187
rect 7668 26167 7670 26187
rect 7716 26167 7718 26187
rect 7740 26167 7742 26187
rect 7836 26167 7838 26187
rect 7884 26167 7886 26187
rect 7932 26167 7934 26187
rect 7956 26167 7958 26187
rect 7980 26167 7982 26187
rect 8028 26167 8030 26187
rect 8196 26167 8198 26187
rect 8244 26167 8246 26187
rect 8268 26167 8270 26187
rect 8292 26167 8294 26187
rect 8340 26167 8342 26187
rect 8364 26167 8366 26187
rect 8388 26167 8390 26187
rect 8436 26167 8438 26187
rect 8460 26167 8462 26187
rect 8556 26167 8558 26187
rect 8604 26167 8606 26187
rect 8652 26167 8654 26187
rect 8700 26167 8702 26187
rect 8724 26167 8726 26187
rect 8748 26167 8750 26187
rect 8820 26167 8822 26187
rect 8844 26167 8846 26187
rect 8868 26167 8870 26187
rect 9516 26167 9518 26187
rect 9612 26167 9614 26187
rect 9660 26167 9662 26187
rect 9684 26167 9686 26187
rect 9708 26167 9710 26187
rect 9756 26167 9758 26187
rect 9780 26167 9782 26187
rect 9804 26167 9806 26187
rect 9852 26167 9854 26187
rect 9876 26167 9878 26187
rect 9900 26167 9902 26187
rect 9948 26167 9950 26187
rect 9972 26167 9974 26187
rect 9996 26167 9998 26187
rect 10068 26167 10070 26187
rect 10092 26167 10094 26187
rect 10116 26167 10118 26187
rect 10164 26167 10166 26187
rect 10188 26167 10190 26187
rect 10212 26167 10214 26187
rect 10284 26167 10286 26187
rect 10308 26167 10310 26187
rect 10332 26167 10334 26187
rect 10380 26167 10382 26187
rect 10404 26167 10406 26187
rect 10428 26167 10430 26187
rect 10476 26167 10478 26187
rect 10500 26167 10502 26187
rect 10524 26167 10526 26187
rect 10572 26167 10574 26187
rect 10596 26167 10598 26187
rect 10620 26167 10622 26187
rect 10668 26167 10670 26187
rect 10692 26167 10694 26187
rect 10716 26167 10718 26187
rect 10788 26167 10790 26187
rect 10836 26167 10838 26187
rect 10956 26167 10958 26187
rect 11052 26167 11054 26187
rect 11076 26167 11078 26187
rect 11124 26167 11126 26187
rect 11172 26167 11174 26187
rect 11220 26167 11222 26187
rect 11340 26167 11342 26187
rect 11436 26167 11438 26187
rect 11532 26167 11534 26187
rect 11580 26167 11582 26187
rect 11628 26167 11630 26187
rect 11676 26167 11678 26187
rect 11724 26167 11726 26187
rect 11772 26167 11774 26187
rect 11796 26167 11798 26187
rect 11892 26167 11894 26187
rect 11988 26167 11990 26187
rect 12060 26167 12062 26187
rect 12132 26167 12134 26187
rect 12228 26167 12230 26187
rect 12276 26167 12278 26187
rect 12324 26167 12326 26187
rect 12420 26167 12422 26187
rect 12444 26167 12446 26187
rect 12492 26167 12494 26187
rect 12516 26167 12518 26187
rect 12540 26167 12542 26187
rect 12588 26167 12590 26187
rect 12636 26167 12638 26187
rect 12732 26167 12734 26187
rect 12756 26167 12758 26187
rect 12804 26167 12806 26187
rect 12828 26167 12830 26187
rect 12852 26167 12854 26187
rect 12900 26167 12902 26187
rect 12948 26167 12950 26187
rect 13044 26167 13046 26187
rect 13068 26167 13070 26187
rect 13116 26167 13118 26187
rect 13284 26167 13286 26187
rect 13332 26167 13334 26187
rect 13428 26167 13430 26187
rect 13524 26167 13526 26187
rect 13572 26167 13574 26187
rect 13644 26167 13646 26187
rect 13668 26167 13670 26187
rect 13764 26167 13766 26187
rect 13812 26167 13814 26187
rect 13860 26167 13862 26187
rect 13908 26167 13910 26187
rect 13956 26167 13958 26187
rect 14004 26167 14006 26187
rect 14100 26167 14102 26187
rect 14196 26167 14198 26187
rect 14292 26167 14294 26187
rect 15132 26167 15134 26187
rect 15180 26167 15182 26187
rect 15228 26167 15230 26187
rect 15252 26167 15254 26187
rect 15324 26167 15326 26187
rect 15396 26167 15398 26187
rect 15420 26167 15422 26187
rect 15492 26167 15494 26187
rect 15540 26167 15542 26187
rect 15636 26167 15638 26187
rect 15660 26167 15662 26187
rect 15708 26167 15710 26187
rect 15732 26167 15734 26187
rect 15756 26167 15758 26187
rect 15804 26167 15806 26187
rect 15828 26167 15830 26187
rect 15852 26167 15854 26187
rect 15900 26167 15902 26187
rect 15948 26167 15950 26187
rect 15996 26167 15998 26187
rect 16044 26167 16046 26187
rect 16092 26167 16094 26187
rect 16260 26167 16262 26187
rect 16308 26167 16310 26187
rect 16332 26167 16334 26187
rect 16356 26167 16358 26187
rect 16404 26167 16406 26187
rect 16452 26167 16454 26187
rect 16548 26167 16550 26187
rect 16572 26167 16574 26187
rect 16620 26167 16622 26187
rect 16668 26167 16670 26187
rect 16716 26167 16718 26187
rect 16764 26167 16766 26187
rect 16801 26182 16804 26187
rect 16825 26182 16828 26187
rect 16836 26182 16838 26187
rect 16811 26168 16814 26182
rect 16835 26168 16838 26182
rect 16812 26167 16814 26168
rect 16884 26167 16886 26187
rect 16908 26167 16911 26184
rect 16980 26167 16982 26187
rect 17052 26167 17054 26187
rect 17196 26167 17198 26187
rect 17220 26167 17222 26187
rect 17292 26167 17294 26187
rect 17316 26167 17318 26187
rect 18084 26167 18086 26187
rect 18132 26167 18134 26187
rect 18396 26167 18398 26187
rect 18492 26167 18494 26187
rect 18516 26167 18518 26187
rect 18564 26167 18566 26187
rect 18612 26167 18614 26187
rect 18660 26167 18662 26187
rect 18708 26167 18710 26187
rect 18756 26167 18758 26187
rect 18804 26167 18806 26187
rect 18852 26167 18854 26187
rect 18900 26167 18902 26187
rect 18996 26167 18998 26187
rect 19020 26167 19022 26187
rect 19092 26167 19094 26187
rect 19116 26167 19118 26187
rect 19140 26167 19142 26187
rect 19188 26167 19190 26187
rect 19236 26167 19238 26187
rect 19332 26167 19334 26187
rect 19476 26167 19478 26187
rect 19620 26167 19622 26187
rect 19716 26167 19718 26187
rect 19788 26167 19790 26187
rect 19836 26167 19838 26187
rect 19860 26167 19862 26187
rect 19884 26167 19886 26187
rect 19932 26167 19934 26187
rect 19956 26167 19958 26187
rect 19980 26167 19982 26187
rect 20028 26167 20030 26187
rect 20052 26167 20054 26187
rect 20076 26167 20078 26187
rect 20148 26167 20150 26187
rect 20172 26167 20174 26187
rect 20196 26167 20198 26187
rect 20268 26167 20270 26187
rect 20292 26167 20294 26187
rect 20388 26167 20390 26187
rect 20412 26167 20414 26187
rect 20508 26167 20510 26187
rect 20556 26167 20558 26187
rect 20604 26167 20606 26187
rect 20916 26167 20918 26187
rect 20964 26167 20966 26187
rect 21012 26167 21014 26187
rect 21060 26167 21062 26187
rect 21084 26167 21086 26187
rect 21108 26167 21110 26187
rect 21204 26167 21206 26187
rect 21300 26167 21302 26187
rect 21324 26167 21326 26187
rect 21444 26167 21446 26187
rect 21468 26167 21470 26187
rect 21564 26167 21566 26187
rect 21612 26167 21614 26187
rect 21684 26167 21686 26187
rect 21708 26167 21710 26187
rect 21828 26167 21830 26187
rect 21924 26167 21926 26187
rect 22023 26184 22037 26187
rect 22044 26184 22047 26187
rect 22068 26167 22070 26187
rect 22188 26167 22190 26187
rect 22212 26167 22214 26187
rect 22873 26182 22876 26187
rect 23004 26184 23006 26187
rect 22883 26168 22886 26182
rect 22884 26167 22886 26168
rect 22980 26167 22983 26184
rect 23004 26167 23007 26184
rect 23052 26167 23054 26187
rect 23076 26167 23078 26187
rect 23100 26167 23102 26187
rect 23148 26167 23150 26187
rect 23244 26167 23246 26187
rect 23295 26184 23309 26187
rect 23316 26184 23319 26187
rect 23340 26167 23342 26187
rect 23412 26167 23414 26187
rect 23556 26167 23558 26187
rect 23628 26167 23630 26187
rect 23652 26167 23654 26187
rect 23676 26167 23678 26187
rect 23724 26167 23726 26187
rect 23772 26167 23774 26187
rect 23820 26167 23822 26187
rect 23868 26167 23870 26187
rect 23916 26167 23918 26187
rect 24012 26167 24014 26187
rect 24084 26167 24086 26187
rect 24396 26167 24398 26187
rect 24447 26184 24461 26187
rect 24492 26167 24494 26187
rect 24516 26167 24518 26187
rect 24588 26167 24590 26187
rect 24612 26167 24614 26187
rect 24708 26167 24710 26187
rect 24732 26167 24734 26187
rect 24756 26167 24758 26187
rect 24852 26167 24854 26187
rect 24876 26167 24878 26187
rect 24972 26167 24974 26187
rect 24996 26167 24998 26187
rect 25092 26167 25094 26187
rect 25260 26167 25262 26187
rect 25308 26167 25310 26187
rect 25356 26167 25358 26187
rect 25380 26167 25382 26187
rect 25404 26167 25406 26187
rect 25452 26167 25454 26187
rect 25500 26167 25502 26187
rect 25596 26167 25598 26187
rect 27049 26182 27052 26187
rect 27060 26182 27062 26187
rect 27059 26168 27062 26182
rect 27108 26167 27110 26187
rect 27156 26184 27158 26187
rect 27156 26167 27159 26184
rect 27324 26167 27326 26187
rect 27396 26167 27398 26187
rect 27420 26167 27422 26187
rect 27540 26167 27542 26187
rect 27564 26167 27566 26187
rect 30564 26167 30566 26187
rect 30660 26167 30662 26187
rect 30711 26184 30725 26187
rect 30780 26167 30782 26187
rect 30804 26167 30806 26187
rect 30841 26167 30875 26168
rect -16319 26163 -15235 26167
rect -16284 26160 -16282 26163
rect -16295 26150 -16291 26158
rect -16305 26144 -16295 26150
rect -17615 26139 -17371 26143
rect -17508 26136 -17506 26139
rect -17508 26119 -17505 26136
rect -17484 26119 -17482 26139
rect -17460 26119 -17458 26139
rect -17388 26119 -17386 26139
rect -17385 26136 -17371 26139
rect -17361 26139 -16291 26143
rect -17361 26136 -17347 26139
rect -17292 26119 -17290 26139
rect -17028 26119 -17026 26139
rect -16932 26119 -16930 26139
rect -16860 26136 -16858 26139
rect -16860 26119 -16857 26136
rect -16836 26119 -16834 26139
rect -16764 26120 -16762 26139
rect -16775 26119 -16741 26120
rect -17529 26115 -16741 26119
rect -17529 26112 -17515 26115
rect -17508 26112 -17505 26115
rect -17484 26112 -17482 26115
rect -17484 26095 -17481 26112
rect -17460 26095 -17458 26115
rect -17388 26095 -17386 26115
rect -17292 26095 -17290 26115
rect -17028 26096 -17026 26115
rect -17063 26095 -17005 26096
rect -16932 26095 -16930 26115
rect -16881 26112 -16867 26115
rect -16860 26112 -16857 26115
rect -16836 26095 -16834 26115
rect -16775 26110 -16772 26115
rect -16764 26110 -16762 26115
rect -16765 26096 -16762 26110
rect -16764 26095 -16762 26096
rect -16740 26095 -16738 26139
rect -16727 26119 -16693 26120
rect -16668 26119 -16666 26139
rect -16631 26134 -16628 26139
rect -16500 26136 -16498 26139
rect -16621 26120 -16618 26134
rect -16620 26119 -16618 26120
rect -16500 26119 -16497 26136
rect -16380 26119 -16378 26139
rect -16356 26119 -16354 26139
rect -16305 26136 -16291 26139
rect -16284 26136 -16281 26160
rect -16284 26119 -16282 26136
rect -16260 26119 -16258 26163
rect -16236 26119 -16234 26163
rect -15324 26143 -15322 26163
rect -15249 26160 -15235 26163
rect -15225 26163 -11203 26167
rect -15225 26160 -15211 26163
rect -15084 26143 -15082 26163
rect -14868 26143 -14866 26163
rect -14772 26143 -14770 26163
rect -14724 26143 -14722 26163
rect -14508 26143 -14506 26163
rect -14436 26143 -14434 26163
rect -14340 26143 -14338 26163
rect -14244 26143 -14242 26163
rect -14172 26143 -14170 26163
rect -14076 26143 -14074 26163
rect -13980 26143 -13978 26163
rect -13932 26143 -13930 26163
rect -13884 26143 -13882 26163
rect -13823 26143 -13741 26144
rect -13716 26143 -13714 26163
rect -13644 26143 -13642 26163
rect -13500 26143 -13498 26163
rect -13356 26143 -13354 26163
rect -13284 26143 -13282 26163
rect -13068 26143 -13066 26163
rect -12828 26143 -12826 26163
rect -12780 26143 -12778 26163
rect -12660 26143 -12658 26163
rect -12564 26143 -12562 26163
rect -12492 26143 -12490 26163
rect -12396 26143 -12394 26163
rect -12348 26143 -12346 26163
rect -12276 26143 -12274 26163
rect -12252 26143 -12250 26163
rect -12156 26143 -12154 26163
rect -12060 26143 -12058 26163
rect -11892 26143 -11890 26163
rect -11844 26143 -11842 26163
rect -11796 26143 -11794 26163
rect -11676 26143 -11674 26163
rect -11580 26143 -11578 26163
rect -11556 26143 -11554 26163
rect -11508 26143 -11506 26163
rect -11460 26143 -11458 26163
rect -11436 26143 -11434 26163
rect -11364 26143 -11362 26163
rect -11340 26143 -11338 26163
rect -11292 26143 -11290 26163
rect -11217 26160 -11203 26163
rect -11193 26163 -6163 26167
rect -11193 26160 -11179 26163
rect -11172 26160 -11169 26163
rect -11207 26143 -11149 26144
rect -11124 26143 -11122 26163
rect -11076 26144 -11074 26163
rect -11111 26143 -11053 26144
rect -11028 26143 -11026 26163
rect -10788 26143 -10786 26163
rect -10751 26158 -10748 26163
rect -10741 26144 -10738 26158
rect -10740 26143 -10738 26144
rect -10668 26143 -10666 26163
rect -10644 26143 -10641 26160
rect -9996 26143 -9994 26163
rect -9708 26143 -9706 26163
rect -9612 26143 -9610 26163
rect -9516 26143 -9514 26163
rect -9468 26143 -9466 26163
rect -9420 26143 -9418 26163
rect -9396 26143 -9394 26163
rect -9372 26143 -9370 26163
rect -9300 26143 -9298 26163
rect -9252 26143 -9250 26163
rect -9132 26143 -9130 26163
rect -9084 26143 -9082 26163
rect -9036 26143 -9034 26163
rect -8988 26143 -8986 26163
rect -8940 26143 -8938 26163
rect -8892 26143 -8890 26163
rect -8772 26143 -8770 26163
rect -8604 26143 -8602 26163
rect -8508 26143 -8506 26163
rect -8484 26143 -8482 26163
rect -8388 26143 -8386 26163
rect -8364 26143 -8362 26163
rect -8340 26143 -8338 26163
rect -8268 26143 -8266 26163
rect -8100 26143 -8098 26163
rect -8052 26143 -8050 26163
rect -7932 26143 -7930 26163
rect -7692 26143 -7690 26163
rect -7620 26143 -7618 26163
rect -7535 26158 -7532 26163
rect -7404 26160 -7402 26163
rect -7525 26144 -7522 26158
rect -7524 26143 -7522 26144
rect -7404 26143 -7401 26160
rect -7356 26143 -7354 26163
rect -7308 26143 -7306 26163
rect -7212 26143 -7210 26163
rect -7188 26143 -7186 26163
rect -7116 26143 -7114 26163
rect -7068 26143 -7066 26163
rect -6972 26143 -6970 26163
rect -6948 26143 -6946 26163
rect -6876 26143 -6874 26163
rect -6852 26143 -6850 26163
rect -6780 26143 -6778 26163
rect -6756 26143 -6754 26163
rect -6660 26143 -6658 26163
rect -6612 26143 -6610 26163
rect -6516 26143 -6514 26163
rect -6492 26143 -6490 26163
rect -6489 26160 -6475 26163
rect -6468 26160 -6465 26163
rect -6420 26143 -6418 26163
rect -6396 26143 -6394 26163
rect -6372 26143 -6370 26163
rect -6324 26143 -6322 26163
rect -6300 26143 -6298 26163
rect -6201 26160 -6187 26163
rect -6180 26160 -6163 26163
rect -6156 26163 16901 26167
rect -6156 26160 -6139 26163
rect -6156 26143 -6154 26160
rect -6060 26143 -6058 26163
rect -5940 26143 -5938 26163
rect -5892 26143 -5890 26163
rect -5652 26143 -5650 26163
rect -5268 26143 -5266 26163
rect -5196 26143 -5194 26163
rect -5172 26143 -5170 26163
rect -5100 26143 -5098 26163
rect -5076 26143 -5074 26163
rect -4980 26143 -4978 26163
rect -4956 26143 -4954 26163
rect -4884 26143 -4882 26163
rect -4860 26143 -4858 26163
rect -4788 26143 -4786 26163
rect -4692 26143 -4690 26163
rect -4644 26143 -4642 26163
rect -4596 26143 -4594 26163
rect -4548 26143 -4546 26163
rect -4308 26143 -4306 26163
rect -4260 26143 -4258 26163
rect -4212 26143 -4210 26163
rect -4175 26158 -4172 26163
rect -4165 26144 -4162 26158
rect -4164 26143 -4162 26144
rect -4116 26143 -4114 26163
rect -4020 26143 -4018 26163
rect -3876 26143 -3874 26163
rect -3732 26143 -3730 26163
rect -3588 26143 -3586 26163
rect -3564 26143 -3562 26163
rect -3516 26143 -3514 26163
rect -3492 26143 -3490 26163
rect -3468 26143 -3466 26163
rect -3420 26143 -3418 26163
rect -3324 26143 -3322 26163
rect -3252 26143 -3250 26163
rect -3228 26143 -3226 26163
rect -3156 26143 -3154 26163
rect -3132 26143 -3130 26163
rect -3060 26143 -3058 26163
rect -3012 26143 -3010 26163
rect -2964 26143 -2962 26163
rect -2916 26143 -2914 26163
rect -2892 26143 -2890 26163
rect -2820 26143 -2818 26163
rect -2796 26143 -2794 26163
rect -2748 26143 -2746 26163
rect -2700 26143 -2698 26163
rect -2604 26143 -2602 26163
rect -2580 26143 -2578 26163
rect -2364 26143 -2362 26163
rect -2268 26143 -2266 26163
rect -2244 26143 -2242 26163
rect -2172 26143 -2170 26163
rect -2148 26143 -2146 26163
rect -2076 26143 -2074 26163
rect -2052 26143 -2050 26163
rect -1980 26143 -1978 26163
rect -1884 26143 -1882 26163
rect -1836 26143 -1834 26163
rect -1716 26143 -1714 26163
rect -1596 26143 -1594 26163
rect -1572 26143 -1570 26163
rect -1476 26143 -1474 26163
rect -1380 26143 -1378 26163
rect -1356 26143 -1354 26163
rect -1308 26143 -1306 26163
rect -1260 26143 -1258 26163
rect -1140 26143 -1138 26163
rect -852 26143 -850 26163
rect -804 26143 -802 26163
rect -756 26143 -754 26163
rect -708 26143 -706 26163
rect -612 26143 -610 26163
rect -588 26143 -586 26163
rect -540 26143 -538 26163
rect -492 26143 -490 26163
rect -444 26143 -442 26163
rect -396 26143 -394 26163
rect -300 26143 -298 26163
rect -276 26143 -274 26163
rect -228 26143 -226 26163
rect 12 26144 14 26163
rect -23 26143 35 26144
rect 108 26143 110 26163
rect 156 26143 158 26163
rect 204 26143 206 26163
rect 228 26143 230 26163
rect 252 26143 254 26163
rect 348 26143 350 26163
rect 468 26143 470 26163
rect 492 26143 494 26163
rect 564 26143 566 26163
rect 588 26143 590 26163
rect 636 26143 638 26163
rect 660 26143 662 26163
rect 732 26143 734 26163
rect 756 26143 758 26163
rect 876 26143 878 26163
rect 972 26143 974 26163
rect 1020 26143 1022 26163
rect 1068 26143 1070 26163
rect 1092 26143 1094 26163
rect 1116 26143 1118 26163
rect 1164 26143 1166 26163
rect 1212 26143 1214 26163
rect 1308 26143 1310 26163
rect 1332 26143 1334 26163
rect 1380 26143 1382 26163
rect 1428 26143 1430 26163
rect 1524 26143 1526 26163
rect 1548 26143 1550 26163
rect 1596 26143 1598 26163
rect 1620 26143 1622 26163
rect 1644 26143 1646 26163
rect 1692 26143 1694 26163
rect 1716 26143 1718 26163
rect 1740 26143 1742 26163
rect 1788 26143 1790 26163
rect 1884 26143 1886 26163
rect 1980 26143 1982 26163
rect 2028 26143 2030 26163
rect 2076 26143 2078 26163
rect 2100 26143 2102 26163
rect 2124 26143 2126 26163
rect 2172 26143 2174 26163
rect 2196 26143 2198 26163
rect 2220 26143 2222 26163
rect 2268 26143 2270 26163
rect 2292 26143 2294 26163
rect 2316 26143 2318 26163
rect 2364 26143 2366 26163
rect 2412 26143 2414 26163
rect 2460 26143 2462 26163
rect 2508 26143 2510 26163
rect 2545 26158 2548 26163
rect 2556 26158 2558 26163
rect 2555 26144 2558 26158
rect 2580 26143 2582 26163
rect 2604 26143 2606 26163
rect 2652 26160 2654 26163
rect 2652 26143 2655 26160
rect 2676 26143 2678 26163
rect 2700 26143 2702 26163
rect 2748 26143 2750 26163
rect 2772 26143 2774 26163
rect 2796 26143 2798 26163
rect 2844 26143 2846 26163
rect 2868 26143 2870 26163
rect 2892 26143 2894 26163
rect 2940 26143 2942 26163
rect 3012 26143 3014 26163
rect 3108 26143 3110 26163
rect 3156 26143 3158 26163
rect 3252 26143 3254 26163
rect 3348 26143 3350 26163
rect 3396 26143 3398 26163
rect 3468 26143 3470 26163
rect 3492 26143 3494 26163
rect 3588 26144 3590 26163
rect 3553 26143 3611 26144
rect 3612 26143 3614 26163
rect 3636 26143 3638 26163
rect 3708 26143 3710 26163
rect 3732 26143 3734 26163
rect 3804 26143 3806 26163
rect 3828 26143 3830 26163
rect 3924 26143 3926 26163
rect 4020 26143 4022 26163
rect 4044 26143 4046 26163
rect 4092 26143 4094 26163
rect 4116 26143 4118 26163
rect 4140 26143 4142 26163
rect 4188 26143 4190 26163
rect 4212 26143 4214 26163
rect 4236 26143 4238 26163
rect 4308 26143 4310 26163
rect 4332 26143 4334 26163
rect 4404 26143 4406 26163
rect 4500 26143 4502 26163
rect 4596 26143 4598 26163
rect 4860 26143 4862 26163
rect 4956 26143 4958 26163
rect 4980 26143 4982 26163
rect 5004 26143 5006 26163
rect 5076 26143 5078 26163
rect 5100 26143 5102 26163
rect 5124 26143 5126 26163
rect 5172 26143 5174 26163
rect 5220 26143 5222 26163
rect 5268 26143 5270 26163
rect 5388 26143 5390 26163
rect 5484 26143 5486 26163
rect 5508 26143 5510 26163
rect 5532 26143 5534 26163
rect 5628 26143 5630 26163
rect 5652 26143 5654 26163
rect 5748 26143 5750 26163
rect 5796 26143 5798 26163
rect 5844 26143 5846 26163
rect 5892 26143 5894 26163
rect 6132 26143 6134 26163
rect 6180 26143 6182 26163
rect 6228 26143 6230 26163
rect 6252 26143 6254 26163
rect 6276 26143 6278 26163
rect 6324 26143 6326 26163
rect 6372 26143 6374 26163
rect 6492 26143 6494 26163
rect 6588 26143 6590 26163
rect 6612 26143 6614 26163
rect 6660 26143 6662 26163
rect 6684 26143 6686 26163
rect 6708 26143 6710 26163
rect 6780 26143 6782 26163
rect 6804 26143 6806 26163
rect 6828 26143 6830 26163
rect 6900 26143 6902 26163
rect 6924 26143 6926 26163
rect 7020 26143 7022 26163
rect 7140 26143 7142 26163
rect 7236 26143 7238 26163
rect 7332 26143 7334 26163
rect 7380 26143 7382 26163
rect 7428 26143 7430 26163
rect 7452 26143 7454 26163
rect 7476 26143 7478 26163
rect 7524 26143 7526 26163
rect 7548 26143 7550 26163
rect 7572 26143 7574 26163
rect 7620 26143 7622 26163
rect 7644 26143 7646 26163
rect 7668 26143 7670 26163
rect 7716 26143 7718 26163
rect 7740 26143 7742 26163
rect 7836 26143 7838 26163
rect 7884 26143 7886 26163
rect 7932 26143 7934 26163
rect 7956 26143 7958 26163
rect 7980 26143 7982 26163
rect 8028 26143 8030 26163
rect 8196 26143 8198 26163
rect 8244 26143 8246 26163
rect 8268 26143 8270 26163
rect 8292 26143 8294 26163
rect 8340 26143 8342 26163
rect 8364 26143 8366 26163
rect 8388 26143 8390 26163
rect 8436 26143 8438 26163
rect 8460 26143 8462 26163
rect 8556 26143 8558 26163
rect 8604 26143 8606 26163
rect 8652 26143 8654 26163
rect 8700 26143 8702 26163
rect 8724 26143 8726 26163
rect 8748 26143 8750 26163
rect 8820 26143 8822 26163
rect 8844 26143 8846 26163
rect 8868 26143 8870 26163
rect 9516 26143 9518 26163
rect 9612 26143 9614 26163
rect 9660 26143 9662 26163
rect 9684 26143 9686 26163
rect 9708 26143 9710 26163
rect 9756 26143 9758 26163
rect 9780 26143 9782 26163
rect 9804 26143 9806 26163
rect 9852 26143 9854 26163
rect 9876 26143 9878 26163
rect 9900 26143 9902 26163
rect 9948 26143 9950 26163
rect 9972 26143 9974 26163
rect 9996 26143 9998 26163
rect 10068 26143 10070 26163
rect 10092 26143 10094 26163
rect 10116 26143 10118 26163
rect 10164 26143 10166 26163
rect 10188 26143 10190 26163
rect 10212 26143 10214 26163
rect 10284 26143 10286 26163
rect 10308 26143 10310 26163
rect 10332 26143 10334 26163
rect 10380 26143 10382 26163
rect 10404 26143 10406 26163
rect 10428 26143 10430 26163
rect 10476 26143 10478 26163
rect 10500 26143 10502 26163
rect 10524 26143 10526 26163
rect 10572 26143 10574 26163
rect 10596 26143 10598 26163
rect 10620 26143 10622 26163
rect 10668 26143 10670 26163
rect 10692 26143 10694 26163
rect 10716 26143 10718 26163
rect 10788 26143 10790 26163
rect 10836 26143 10838 26163
rect 10956 26143 10958 26163
rect 11052 26143 11054 26163
rect 11076 26143 11078 26163
rect 11124 26143 11126 26163
rect 11172 26143 11174 26163
rect 11220 26143 11222 26163
rect 11340 26143 11342 26163
rect 11436 26143 11438 26163
rect 11532 26143 11534 26163
rect 11580 26143 11582 26163
rect 11628 26143 11630 26163
rect 11676 26143 11678 26163
rect 11724 26143 11726 26163
rect 11772 26143 11774 26163
rect 11796 26143 11798 26163
rect 11892 26143 11894 26163
rect 11988 26143 11990 26163
rect 12060 26143 12062 26163
rect 12132 26143 12134 26163
rect 12228 26143 12230 26163
rect 12276 26143 12278 26163
rect 12324 26143 12326 26163
rect 12420 26143 12422 26163
rect 12444 26143 12446 26163
rect 12492 26143 12494 26163
rect 12516 26143 12518 26163
rect 12540 26143 12542 26163
rect 12588 26143 12590 26163
rect 12636 26143 12638 26163
rect 12732 26143 12734 26163
rect 12756 26143 12758 26163
rect 12804 26143 12806 26163
rect 12828 26143 12830 26163
rect 12852 26143 12854 26163
rect 12900 26143 12902 26163
rect 12948 26143 12950 26163
rect 13044 26143 13046 26163
rect 13068 26143 13070 26163
rect 13116 26143 13118 26163
rect 13284 26143 13286 26163
rect 13332 26143 13334 26163
rect 13428 26143 13430 26163
rect 13524 26143 13526 26163
rect 13572 26143 13574 26163
rect 13644 26143 13646 26163
rect 13668 26143 13670 26163
rect 13764 26143 13766 26163
rect 13812 26143 13814 26163
rect 13860 26143 13862 26163
rect 13908 26143 13910 26163
rect 13956 26143 13958 26163
rect 14004 26143 14006 26163
rect 14100 26143 14102 26163
rect 14196 26143 14198 26163
rect 14292 26143 14294 26163
rect 15132 26143 15134 26163
rect 15180 26143 15182 26163
rect 15228 26143 15230 26163
rect 15252 26143 15254 26163
rect 15324 26143 15326 26163
rect 15396 26143 15398 26163
rect 15420 26143 15422 26163
rect 15492 26143 15494 26163
rect 15540 26143 15542 26163
rect 15636 26143 15638 26163
rect 15660 26143 15662 26163
rect 15708 26143 15710 26163
rect 15732 26143 15734 26163
rect 15756 26143 15758 26163
rect 15804 26143 15806 26163
rect 15828 26143 15830 26163
rect 15852 26143 15854 26163
rect 15900 26143 15902 26163
rect 15948 26143 15950 26163
rect 15996 26143 15998 26163
rect 16044 26143 16046 26163
rect 16092 26143 16094 26163
rect 16260 26143 16262 26163
rect 16308 26143 16310 26163
rect 16332 26143 16334 26163
rect 16356 26143 16358 26163
rect 16404 26143 16406 26163
rect 16452 26143 16454 26163
rect 16548 26143 16550 26163
rect 16572 26143 16574 26163
rect 16620 26143 16622 26163
rect 16668 26143 16670 26163
rect 16716 26143 16718 26163
rect 16764 26143 16766 26163
rect 16812 26143 16814 26163
rect 16884 26143 16886 26163
rect 16887 26160 16901 26163
rect 16908 26163 22973 26167
rect 16908 26160 16925 26163
rect 16908 26143 16910 26160
rect 16980 26143 16982 26163
rect 17052 26143 17054 26163
rect 17196 26143 17198 26163
rect 17220 26143 17222 26163
rect 17292 26143 17294 26163
rect 17316 26143 17318 26163
rect 18084 26143 18086 26163
rect 18132 26143 18134 26163
rect 18396 26143 18398 26163
rect 18492 26143 18494 26163
rect 18516 26143 18518 26163
rect 18564 26143 18566 26163
rect 18612 26143 18614 26163
rect 18660 26143 18662 26163
rect 18708 26143 18710 26163
rect 18756 26143 18758 26163
rect 18804 26143 18806 26163
rect 18852 26143 18854 26163
rect 18900 26143 18902 26163
rect 18996 26143 18998 26163
rect 19020 26143 19022 26163
rect 19092 26143 19094 26163
rect 19116 26143 19118 26163
rect 19140 26143 19142 26163
rect 19188 26143 19190 26163
rect 19236 26143 19238 26163
rect 19332 26143 19334 26163
rect 19476 26143 19478 26163
rect 19620 26143 19622 26163
rect 19716 26143 19718 26163
rect 19788 26143 19790 26163
rect 19836 26143 19838 26163
rect 19860 26143 19862 26163
rect 19884 26143 19886 26163
rect 19932 26143 19934 26163
rect 19956 26143 19958 26163
rect 19980 26143 19982 26163
rect 20028 26143 20030 26163
rect 20052 26143 20054 26163
rect 20076 26143 20078 26163
rect 20148 26143 20150 26163
rect 20172 26143 20174 26163
rect 20196 26143 20198 26163
rect 20268 26143 20270 26163
rect 20292 26143 20294 26163
rect 20388 26143 20390 26163
rect 20412 26143 20414 26163
rect 20508 26143 20510 26163
rect 20556 26143 20558 26163
rect 20604 26143 20606 26163
rect 20916 26143 20918 26163
rect 20964 26143 20966 26163
rect 21012 26143 21014 26163
rect 21060 26143 21062 26163
rect 21084 26143 21086 26163
rect 21108 26143 21110 26163
rect 21204 26143 21206 26163
rect 21300 26143 21302 26163
rect 21324 26143 21326 26163
rect 21444 26143 21446 26163
rect 21468 26143 21470 26163
rect 21564 26143 21566 26163
rect 21612 26143 21614 26163
rect 21684 26143 21686 26163
rect 21708 26143 21710 26163
rect 21828 26143 21830 26163
rect 21924 26143 21926 26163
rect 22068 26143 22070 26163
rect 22188 26143 22190 26163
rect 22212 26143 22214 26163
rect 22884 26143 22886 26163
rect 22959 26160 22973 26163
rect 22980 26163 27125 26167
rect 22980 26160 22997 26163
rect 23004 26160 23007 26163
rect 22980 26143 22982 26160
rect 23052 26144 23054 26163
rect 23017 26143 23075 26144
rect 23076 26143 23078 26163
rect 23100 26143 23102 26163
rect 23148 26143 23150 26163
rect 23244 26143 23246 26163
rect 23340 26143 23342 26163
rect 23412 26143 23414 26163
rect 23556 26143 23558 26163
rect 23628 26143 23630 26163
rect 23652 26143 23654 26163
rect 23676 26143 23678 26163
rect 23724 26143 23726 26163
rect 23772 26143 23774 26163
rect 23820 26143 23822 26163
rect 23868 26143 23870 26163
rect 23916 26143 23918 26163
rect 24012 26143 24014 26163
rect 24084 26143 24086 26163
rect 24396 26143 24398 26163
rect 24492 26143 24494 26163
rect 24516 26143 24518 26163
rect 24588 26143 24590 26163
rect 24612 26143 24614 26163
rect 24708 26143 24710 26163
rect 24732 26143 24734 26163
rect 24756 26143 24758 26163
rect 24852 26143 24854 26163
rect 24876 26143 24878 26163
rect 24972 26143 24974 26163
rect 24996 26143 24998 26163
rect 25092 26144 25094 26163
rect 25057 26143 25115 26144
rect 25260 26143 25262 26163
rect 25308 26143 25310 26163
rect 25356 26143 25358 26163
rect 25380 26143 25382 26163
rect 25404 26143 25406 26163
rect 25452 26143 25454 26163
rect 25500 26143 25502 26163
rect 25596 26143 25598 26163
rect 27108 26143 27110 26163
rect 27111 26160 27125 26163
rect 27135 26163 30875 26167
rect 27135 26160 27149 26163
rect 27156 26160 27159 26163
rect 27324 26143 27326 26163
rect 27396 26143 27398 26163
rect 27420 26143 27422 26163
rect 27540 26143 27542 26163
rect 27564 26143 27566 26163
rect 30564 26143 30566 26163
rect 30660 26143 30662 26163
rect 30780 26143 30782 26163
rect 30804 26144 30806 26163
rect 30793 26143 30827 26144
rect -16233 26139 -10651 26143
rect -16233 26136 -16219 26139
rect -15324 26119 -15322 26139
rect -15084 26119 -15082 26139
rect -14868 26119 -14866 26139
rect -14772 26119 -14770 26139
rect -14724 26119 -14722 26139
rect -14508 26119 -14506 26139
rect -14436 26119 -14434 26139
rect -14340 26119 -14338 26139
rect -14244 26119 -14242 26139
rect -14172 26119 -14170 26139
rect -14076 26119 -14074 26139
rect -13980 26119 -13978 26139
rect -13932 26119 -13930 26139
rect -13884 26119 -13882 26139
rect -13799 26134 -13796 26139
rect -13716 26136 -13714 26139
rect -13789 26120 -13786 26134
rect -13788 26119 -13786 26120
rect -13716 26119 -13713 26136
rect -13644 26119 -13642 26139
rect -13500 26119 -13498 26139
rect -13356 26119 -13354 26139
rect -13284 26119 -13282 26139
rect -13247 26119 -13213 26120
rect -13068 26119 -13066 26139
rect -12828 26119 -12826 26139
rect -12780 26119 -12778 26139
rect -12660 26119 -12658 26139
rect -12564 26119 -12562 26139
rect -12492 26119 -12490 26139
rect -12396 26119 -12394 26139
rect -12348 26119 -12346 26139
rect -12276 26119 -12274 26139
rect -12252 26119 -12250 26139
rect -12156 26119 -12154 26139
rect -12060 26119 -12058 26139
rect -11999 26119 -11965 26120
rect -11892 26119 -11890 26139
rect -11844 26119 -11842 26139
rect -11841 26136 -11827 26139
rect -11796 26119 -11794 26139
rect -11676 26119 -11674 26139
rect -11580 26119 -11578 26139
rect -11556 26119 -11554 26139
rect -11508 26119 -11506 26139
rect -11460 26119 -11458 26139
rect -11436 26119 -11434 26139
rect -11364 26119 -11362 26139
rect -11340 26119 -11338 26139
rect -11292 26119 -11290 26139
rect -11207 26134 -11204 26139
rect -11197 26120 -11194 26134
rect -11196 26119 -11194 26120
rect -11124 26119 -11122 26139
rect -11087 26134 -11084 26139
rect -11076 26136 -11074 26139
rect -11076 26134 -11073 26136
rect -11101 26126 -11097 26134
rect -11087 26126 -11083 26134
rect -11101 26120 -11087 26126
rect -11077 26120 -11073 26134
rect -11100 26119 -11097 26120
rect -11028 26119 -11026 26139
rect -11004 26119 -11001 26136
rect -10788 26119 -10786 26139
rect -10740 26119 -10738 26139
rect -10668 26119 -10666 26139
rect -10665 26136 -10651 26139
rect -10644 26139 -7435 26143
rect -10644 26136 -10627 26139
rect -10644 26119 -10642 26136
rect -9996 26119 -9994 26139
rect -9708 26119 -9706 26139
rect -9612 26119 -9610 26139
rect -9516 26119 -9514 26139
rect -9468 26119 -9466 26139
rect -9420 26119 -9418 26139
rect -9396 26119 -9394 26139
rect -9372 26119 -9370 26139
rect -9300 26119 -9298 26139
rect -9252 26119 -9250 26139
rect -9132 26119 -9130 26139
rect -9084 26119 -9082 26139
rect -9036 26119 -9034 26139
rect -8988 26119 -8986 26139
rect -8940 26119 -8938 26139
rect -8892 26119 -8890 26139
rect -8772 26119 -8770 26139
rect -8604 26119 -8602 26139
rect -8508 26119 -8506 26139
rect -8484 26119 -8482 26139
rect -8388 26119 -8386 26139
rect -8364 26119 -8362 26139
rect -8340 26119 -8338 26139
rect -8268 26119 -8266 26139
rect -8100 26119 -8098 26139
rect -8052 26119 -8050 26139
rect -7932 26119 -7930 26139
rect -7692 26119 -7690 26139
rect -7620 26119 -7618 26139
rect -7524 26119 -7522 26139
rect -7449 26136 -7435 26139
rect -7425 26139 -4075 26143
rect -7425 26136 -7411 26139
rect -7404 26136 -7401 26139
rect -7356 26119 -7354 26139
rect -7308 26119 -7306 26139
rect -7212 26119 -7210 26139
rect -7188 26119 -7186 26139
rect -7116 26119 -7114 26139
rect -7068 26119 -7066 26139
rect -6972 26119 -6970 26139
rect -6948 26119 -6946 26139
rect -6876 26119 -6874 26139
rect -6852 26119 -6850 26139
rect -6780 26119 -6778 26139
rect -6756 26119 -6754 26139
rect -6660 26119 -6658 26139
rect -6612 26119 -6610 26139
rect -6516 26119 -6514 26139
rect -6492 26119 -6490 26139
rect -6420 26119 -6418 26139
rect -6396 26119 -6394 26139
rect -6372 26119 -6370 26139
rect -6324 26119 -6322 26139
rect -6300 26120 -6298 26139
rect -6311 26119 -6277 26120
rect -6156 26119 -6154 26139
rect -6060 26119 -6058 26139
rect -5940 26119 -5938 26139
rect -5892 26119 -5890 26139
rect -5652 26119 -5650 26139
rect -5268 26119 -5266 26139
rect -5196 26119 -5194 26139
rect -5172 26119 -5170 26139
rect -5100 26119 -5098 26139
rect -5076 26119 -5074 26139
rect -4980 26119 -4978 26139
rect -4956 26119 -4954 26139
rect -4884 26119 -4882 26139
rect -4860 26119 -4858 26139
rect -4788 26119 -4786 26139
rect -4692 26119 -4690 26139
rect -4679 26119 -4645 26120
rect -4644 26119 -4642 26139
rect -4596 26119 -4594 26139
rect -4548 26119 -4546 26139
rect -4308 26119 -4306 26139
rect -4260 26119 -4258 26139
rect -4212 26119 -4210 26139
rect -4164 26119 -4162 26139
rect -4116 26119 -4114 26139
rect -4089 26136 -4075 26139
rect -4065 26139 2621 26143
rect -4065 26136 -4051 26139
rect -4020 26119 -4018 26139
rect -3876 26119 -3874 26139
rect -3732 26119 -3730 26139
rect -3588 26119 -3586 26139
rect -3564 26119 -3562 26139
rect -3516 26119 -3514 26139
rect -3492 26119 -3490 26139
rect -3468 26119 -3466 26139
rect -3420 26119 -3418 26139
rect -3324 26119 -3322 26139
rect -3252 26119 -3250 26139
rect -3228 26119 -3226 26139
rect -3156 26119 -3154 26139
rect -3132 26119 -3130 26139
rect -3060 26119 -3058 26139
rect -3012 26119 -3010 26139
rect -2964 26119 -2962 26139
rect -2916 26119 -2914 26139
rect -2892 26119 -2890 26139
rect -2820 26119 -2818 26139
rect -2796 26119 -2794 26139
rect -2748 26120 -2746 26139
rect -2783 26119 -2725 26120
rect -2700 26119 -2698 26139
rect -2604 26119 -2602 26139
rect -2580 26119 -2578 26139
rect -2364 26119 -2362 26139
rect -2268 26119 -2266 26139
rect -2244 26119 -2242 26139
rect -2172 26119 -2170 26139
rect -2148 26119 -2146 26139
rect -2076 26119 -2074 26139
rect -2052 26119 -2050 26139
rect -1980 26119 -1978 26139
rect -1884 26119 -1882 26139
rect -1836 26119 -1834 26139
rect -1716 26119 -1714 26139
rect -1596 26119 -1594 26139
rect -1572 26119 -1570 26139
rect -1476 26119 -1474 26139
rect -1380 26119 -1378 26139
rect -1356 26119 -1354 26139
rect -1308 26119 -1306 26139
rect -1260 26119 -1258 26139
rect -1140 26119 -1138 26139
rect -852 26119 -850 26139
rect -804 26119 -802 26139
rect -756 26119 -754 26139
rect -708 26119 -706 26139
rect -612 26119 -610 26139
rect -588 26119 -586 26139
rect -540 26119 -538 26139
rect -492 26119 -490 26139
rect -444 26119 -442 26139
rect -396 26119 -394 26139
rect -300 26119 -298 26139
rect -276 26119 -274 26139
rect -228 26119 -226 26139
rect -23 26134 -20 26139
rect 1 26134 4 26139
rect 12 26134 14 26139
rect -13 26120 -10 26134
rect 11 26120 14 26134
rect 108 26136 110 26139
rect -12 26119 -10 26120
rect 108 26119 111 26136
rect 156 26119 158 26139
rect 204 26119 206 26139
rect 228 26119 230 26139
rect 252 26119 254 26139
rect 348 26119 350 26139
rect 468 26119 470 26139
rect 492 26119 494 26139
rect 564 26119 566 26139
rect 588 26119 590 26139
rect 636 26119 638 26139
rect 660 26119 662 26139
rect 732 26119 734 26139
rect 756 26119 758 26139
rect 876 26120 878 26139
rect 841 26119 899 26120
rect 972 26119 974 26139
rect 1020 26119 1022 26139
rect 1068 26119 1070 26139
rect 1092 26119 1094 26139
rect 1116 26119 1118 26139
rect 1164 26119 1166 26139
rect 1212 26119 1214 26139
rect 1308 26119 1310 26139
rect 1332 26119 1334 26139
rect 1380 26119 1382 26139
rect 1428 26119 1430 26139
rect 1465 26119 1523 26120
rect 1524 26119 1526 26139
rect 1548 26119 1550 26139
rect 1596 26119 1598 26139
rect 1620 26119 1622 26139
rect 1644 26119 1646 26139
rect 1692 26119 1694 26139
rect 1716 26119 1718 26139
rect 1740 26119 1742 26139
rect 1788 26119 1790 26139
rect 1884 26119 1886 26139
rect 1980 26119 1982 26139
rect 2028 26119 2030 26139
rect 2076 26119 2078 26139
rect 2100 26119 2102 26139
rect 2124 26119 2126 26139
rect 2172 26119 2174 26139
rect 2196 26119 2198 26139
rect 2220 26119 2222 26139
rect 2268 26119 2270 26139
rect 2292 26119 2294 26139
rect 2316 26119 2318 26139
rect 2364 26119 2366 26139
rect 2412 26119 2414 26139
rect 2460 26119 2462 26139
rect 2508 26119 2510 26139
rect 2580 26119 2582 26139
rect 2604 26119 2606 26139
rect 2607 26136 2621 26139
rect 2631 26139 30827 26143
rect 2631 26136 2645 26139
rect 2652 26136 2655 26139
rect 2676 26119 2678 26139
rect 2700 26119 2702 26139
rect 2748 26119 2750 26139
rect 2772 26119 2774 26139
rect 2796 26119 2798 26139
rect 2844 26119 2846 26139
rect 2868 26119 2870 26139
rect 2892 26119 2894 26139
rect 2940 26119 2942 26139
rect 3012 26119 3014 26139
rect 3108 26119 3110 26139
rect 3156 26119 3158 26139
rect 3252 26119 3254 26139
rect 3348 26119 3350 26139
rect 3396 26119 3398 26139
rect 3468 26119 3470 26139
rect 3492 26119 3494 26139
rect 3553 26134 3556 26139
rect 3577 26134 3580 26139
rect 3588 26134 3590 26139
rect 3563 26120 3566 26134
rect 3587 26120 3590 26134
rect 3564 26119 3566 26120
rect 3612 26119 3614 26139
rect 3636 26119 3638 26139
rect 3660 26119 3663 26136
rect 3708 26119 3710 26139
rect 3732 26119 3734 26139
rect 3804 26119 3806 26139
rect 3828 26119 3830 26139
rect 3924 26119 3926 26139
rect 4020 26119 4022 26139
rect 4044 26119 4046 26139
rect 4092 26119 4094 26139
rect 4116 26119 4118 26139
rect 4140 26119 4142 26139
rect 4188 26119 4190 26139
rect 4212 26119 4214 26139
rect 4236 26119 4238 26139
rect 4308 26119 4310 26139
rect 4332 26119 4334 26139
rect 4404 26119 4406 26139
rect 4500 26119 4502 26139
rect 4596 26119 4598 26139
rect 4860 26119 4862 26139
rect 4956 26119 4958 26139
rect 4980 26119 4982 26139
rect 5004 26119 5006 26139
rect 5076 26119 5078 26139
rect 5100 26119 5102 26139
rect 5124 26119 5126 26139
rect 5172 26119 5174 26139
rect 5220 26119 5222 26139
rect 5268 26119 5270 26139
rect 5388 26119 5390 26139
rect 5484 26119 5486 26139
rect 5508 26119 5510 26139
rect 5532 26119 5534 26139
rect 5628 26119 5630 26139
rect 5652 26119 5654 26139
rect 5748 26119 5750 26139
rect 5796 26119 5798 26139
rect 5844 26119 5846 26139
rect 5892 26119 5894 26139
rect 6039 26136 6053 26139
rect 6132 26119 6134 26139
rect 6180 26119 6182 26139
rect 6228 26119 6230 26139
rect 6252 26119 6254 26139
rect 6276 26119 6278 26139
rect 6324 26119 6326 26139
rect 6372 26119 6374 26139
rect 6492 26119 6494 26139
rect 6588 26119 6590 26139
rect 6612 26119 6614 26139
rect 6660 26119 6662 26139
rect 6684 26119 6686 26139
rect 6708 26119 6710 26139
rect 6780 26119 6782 26139
rect 6804 26119 6806 26139
rect 6828 26119 6830 26139
rect 6900 26119 6902 26139
rect 6924 26119 6926 26139
rect 7020 26119 7022 26139
rect 7140 26119 7142 26139
rect 7236 26119 7238 26139
rect 7332 26119 7334 26139
rect 7380 26119 7382 26139
rect 7428 26119 7430 26139
rect 7452 26119 7454 26139
rect 7476 26119 7478 26139
rect 7524 26119 7526 26139
rect 7548 26119 7550 26139
rect 7572 26119 7574 26139
rect 7620 26119 7622 26139
rect 7644 26119 7646 26139
rect 7668 26119 7670 26139
rect 7716 26119 7718 26139
rect 7740 26119 7742 26139
rect 7836 26119 7838 26139
rect 7884 26119 7886 26139
rect 7932 26119 7934 26139
rect 7956 26119 7958 26139
rect 7980 26119 7982 26139
rect 8028 26119 8030 26139
rect 8196 26119 8198 26139
rect 8244 26119 8246 26139
rect 8268 26119 8270 26139
rect 8292 26119 8294 26139
rect 8340 26119 8342 26139
rect 8364 26119 8366 26139
rect 8388 26119 8390 26139
rect 8436 26119 8438 26139
rect 8460 26119 8462 26139
rect 8556 26119 8558 26139
rect 8604 26119 8606 26139
rect 8652 26119 8654 26139
rect 8700 26119 8702 26139
rect 8724 26119 8726 26139
rect 8748 26119 8750 26139
rect 8820 26119 8822 26139
rect 8844 26119 8846 26139
rect 8868 26119 8870 26139
rect 9516 26119 9518 26139
rect 9612 26119 9614 26139
rect 9660 26119 9662 26139
rect 9684 26119 9686 26139
rect 9708 26119 9710 26139
rect 9756 26119 9758 26139
rect 9780 26119 9782 26139
rect 9804 26119 9806 26139
rect 9852 26119 9854 26139
rect 9876 26119 9878 26139
rect 9900 26119 9902 26139
rect 9948 26119 9950 26139
rect 9972 26119 9974 26139
rect 9996 26119 9998 26139
rect 10068 26119 10070 26139
rect 10092 26119 10094 26139
rect 10116 26119 10118 26139
rect 10164 26119 10166 26139
rect 10188 26119 10190 26139
rect 10212 26119 10214 26139
rect 10284 26119 10286 26139
rect 10308 26119 10310 26139
rect 10332 26119 10334 26139
rect 10380 26119 10382 26139
rect 10404 26119 10406 26139
rect 10428 26119 10430 26139
rect 10476 26119 10478 26139
rect 10500 26119 10502 26139
rect 10524 26119 10526 26139
rect 10572 26119 10574 26139
rect 10596 26119 10598 26139
rect 10620 26119 10622 26139
rect 10668 26119 10670 26139
rect 10692 26119 10694 26139
rect 10716 26119 10718 26139
rect 10788 26119 10790 26139
rect 10836 26119 10838 26139
rect 10956 26119 10958 26139
rect 11052 26119 11054 26139
rect 11076 26119 11078 26139
rect 11124 26119 11126 26139
rect 11172 26119 11174 26139
rect 11220 26119 11222 26139
rect 11340 26119 11342 26139
rect 11436 26119 11438 26139
rect 11532 26119 11534 26139
rect 11580 26119 11582 26139
rect 11628 26119 11630 26139
rect 11676 26119 11678 26139
rect 11724 26119 11726 26139
rect 11772 26119 11774 26139
rect 11796 26119 11798 26139
rect 11892 26119 11894 26139
rect 11988 26119 11990 26139
rect 12060 26119 12062 26139
rect 12132 26119 12134 26139
rect 12228 26119 12230 26139
rect 12276 26119 12278 26139
rect 12324 26119 12326 26139
rect 12420 26119 12422 26139
rect 12444 26119 12446 26139
rect 12492 26119 12494 26139
rect 12516 26119 12518 26139
rect 12540 26119 12542 26139
rect 12588 26119 12590 26139
rect 12636 26119 12638 26139
rect 12732 26119 12734 26139
rect 12756 26119 12758 26139
rect 12804 26119 12806 26139
rect 12828 26119 12830 26139
rect 12852 26119 12854 26139
rect 12900 26119 12902 26139
rect 12948 26119 12950 26139
rect 13044 26119 13046 26139
rect 13068 26119 13070 26139
rect 13116 26119 13118 26139
rect 13284 26119 13286 26139
rect 13332 26119 13334 26139
rect 13428 26119 13430 26139
rect 13524 26119 13526 26139
rect 13572 26119 13574 26139
rect 13644 26119 13646 26139
rect 13668 26119 13670 26139
rect 13764 26119 13766 26139
rect 13812 26119 13814 26139
rect 13860 26119 13862 26139
rect 13908 26119 13910 26139
rect 13956 26119 13958 26139
rect 14004 26119 14006 26139
rect 14100 26119 14102 26139
rect 14196 26119 14198 26139
rect 14292 26119 14294 26139
rect 15132 26119 15134 26139
rect 15180 26119 15182 26139
rect 15228 26119 15230 26139
rect 15252 26119 15254 26139
rect 15324 26119 15326 26139
rect 15396 26119 15398 26139
rect 15420 26119 15422 26139
rect 15492 26119 15494 26139
rect 15540 26119 15542 26139
rect 15636 26119 15638 26139
rect 15660 26119 15662 26139
rect 15708 26119 15710 26139
rect 15732 26119 15734 26139
rect 15756 26119 15758 26139
rect 15804 26119 15806 26139
rect 15828 26119 15830 26139
rect 15852 26119 15854 26139
rect 15900 26119 15902 26139
rect 15948 26119 15950 26139
rect 15996 26119 15998 26139
rect 16044 26119 16046 26139
rect 16092 26119 16094 26139
rect 16260 26119 16262 26139
rect 16308 26119 16310 26139
rect 16332 26119 16334 26139
rect 16356 26119 16358 26139
rect 16404 26119 16406 26139
rect 16452 26119 16454 26139
rect 16548 26119 16550 26139
rect 16572 26119 16574 26139
rect 16620 26119 16622 26139
rect 16668 26119 16670 26139
rect 16716 26119 16718 26139
rect 16764 26119 16766 26139
rect 16812 26119 16814 26139
rect 16884 26119 16886 26139
rect 16908 26119 16910 26139
rect 16980 26119 16982 26139
rect 17052 26119 17054 26139
rect 17196 26119 17198 26139
rect 17220 26119 17222 26139
rect 17292 26119 17294 26139
rect 17316 26119 17318 26139
rect 18084 26119 18086 26139
rect 18132 26119 18134 26139
rect 18396 26119 18398 26139
rect 18492 26119 18494 26139
rect 18516 26119 18518 26139
rect 18564 26119 18566 26139
rect 18612 26119 18614 26139
rect 18660 26119 18662 26139
rect 18708 26119 18710 26139
rect 18756 26119 18758 26139
rect 18804 26119 18806 26139
rect 18852 26119 18854 26139
rect 18900 26119 18902 26139
rect 18996 26119 18998 26139
rect 19020 26119 19022 26139
rect 19092 26119 19094 26139
rect 19116 26119 19118 26139
rect 19140 26119 19142 26139
rect 19188 26119 19190 26139
rect 19236 26119 19238 26139
rect 19332 26119 19334 26139
rect 19476 26119 19478 26139
rect 19620 26119 19622 26139
rect 19716 26119 19718 26139
rect 19788 26119 19790 26139
rect 19836 26119 19838 26139
rect 19860 26119 19862 26139
rect 19884 26119 19886 26139
rect 19932 26119 19934 26139
rect 19956 26119 19958 26139
rect 19980 26119 19982 26139
rect 20028 26119 20030 26139
rect 20052 26119 20054 26139
rect 20076 26119 20078 26139
rect 20148 26119 20150 26139
rect 20172 26119 20174 26139
rect 20196 26119 20198 26139
rect 20268 26119 20270 26139
rect 20292 26119 20294 26139
rect 20388 26119 20390 26139
rect 20412 26119 20414 26139
rect 20508 26119 20510 26139
rect 20556 26119 20558 26139
rect 20604 26119 20606 26139
rect 20916 26119 20918 26139
rect 20964 26119 20966 26139
rect 21012 26119 21014 26139
rect 21060 26119 21062 26139
rect 21084 26119 21086 26139
rect 21108 26119 21110 26139
rect 21204 26119 21206 26139
rect 21300 26119 21302 26139
rect 21324 26119 21326 26139
rect 21444 26119 21446 26139
rect 21468 26119 21470 26139
rect 21564 26119 21566 26139
rect 21612 26119 21614 26139
rect 21684 26119 21686 26139
rect 21708 26119 21710 26139
rect 21828 26119 21830 26139
rect 21924 26119 21926 26139
rect 22068 26119 22070 26139
rect 22188 26119 22190 26139
rect 22212 26119 22214 26139
rect 22884 26119 22886 26139
rect 22980 26119 22982 26139
rect 23041 26134 23044 26139
rect 23052 26134 23054 26139
rect 23051 26120 23054 26134
rect 23076 26119 23078 26139
rect 23100 26119 23102 26139
rect 23148 26136 23150 26139
rect 23124 26119 23127 26136
rect 23148 26119 23151 26136
rect 23244 26119 23246 26139
rect 23340 26119 23342 26139
rect 23412 26119 23414 26139
rect 23556 26119 23558 26139
rect 23628 26119 23630 26139
rect 23652 26119 23654 26139
rect 23676 26119 23678 26139
rect 23724 26119 23726 26139
rect 23772 26119 23774 26139
rect 23820 26119 23822 26139
rect 23868 26119 23870 26139
rect 23916 26119 23918 26139
rect 24012 26119 24014 26139
rect 24084 26119 24086 26139
rect 24396 26119 24398 26139
rect 24492 26119 24494 26139
rect 24516 26119 24518 26139
rect 24588 26119 24590 26139
rect 24612 26119 24614 26139
rect 24708 26119 24710 26139
rect 24732 26119 24734 26139
rect 24756 26119 24758 26139
rect 24852 26119 24854 26139
rect 24876 26119 24878 26139
rect 24972 26119 24974 26139
rect 24996 26119 24998 26139
rect 25057 26134 25060 26139
rect 25081 26134 25084 26139
rect 25092 26134 25094 26139
rect 25067 26120 25070 26134
rect 25091 26120 25094 26134
rect 25068 26119 25070 26120
rect 25164 26119 25167 26136
rect 25260 26119 25262 26139
rect 25308 26119 25310 26139
rect 25356 26119 25358 26139
rect 25380 26119 25382 26139
rect 25404 26119 25406 26139
rect 25452 26119 25454 26139
rect 25500 26119 25502 26139
rect 25596 26119 25598 26139
rect 27108 26119 27110 26139
rect 27324 26119 27326 26139
rect 27396 26119 27398 26139
rect 27420 26119 27422 26139
rect 27540 26119 27542 26139
rect 27564 26119 27566 26139
rect 30564 26119 30566 26139
rect 30660 26119 30662 26139
rect 30780 26120 30782 26139
rect 30793 26134 30796 26139
rect 30804 26134 30806 26139
rect 30803 26120 30806 26134
rect 30769 26119 30803 26120
rect -16727 26115 -16531 26119
rect -16668 26112 -16666 26115
rect -16620 26112 -16618 26115
rect -16545 26112 -16531 26115
rect -16521 26115 -13699 26119
rect -16521 26112 -16507 26115
rect -16500 26112 -16497 26115
rect -16703 26095 -16675 26096
rect -17505 26091 -16675 26095
rect -17505 26088 -17491 26091
rect -17484 26088 -17481 26091
rect -17460 26088 -17458 26091
rect -17460 26071 -17457 26088
rect -17388 26071 -17386 26091
rect -17292 26072 -17290 26091
rect -17039 26086 -17036 26091
rect -17028 26086 -17026 26091
rect -17029 26072 -17026 26086
rect -16932 26088 -16930 26091
rect -17303 26071 -17269 26072
rect -17159 26071 -17101 26072
rect -16932 26071 -16929 26088
rect -16836 26071 -16834 26091
rect -16764 26071 -16762 26091
rect -16740 26071 -16738 26091
rect -16689 26088 -16675 26091
rect -16668 26088 -16665 26112
rect -16620 26095 -16617 26112
rect -16380 26095 -16378 26115
rect -16356 26095 -16354 26115
rect -16284 26095 -16282 26115
rect -16260 26095 -16258 26115
rect -16236 26095 -16234 26115
rect -15324 26095 -15322 26115
rect -15084 26095 -15082 26115
rect -14868 26095 -14866 26115
rect -14772 26095 -14770 26115
rect -14724 26095 -14722 26115
rect -14508 26095 -14506 26115
rect -14436 26095 -14434 26115
rect -14340 26095 -14338 26115
rect -14244 26095 -14242 26115
rect -14172 26095 -14170 26115
rect -14076 26095 -14074 26115
rect -13980 26095 -13978 26115
rect -13932 26095 -13930 26115
rect -13884 26095 -13882 26115
rect -13788 26095 -13786 26115
rect -13737 26112 -13723 26115
rect -13716 26112 -13699 26115
rect -13689 26115 -11107 26119
rect -13689 26112 -13675 26115
rect -13644 26096 -13642 26115
rect -13679 26095 -13621 26096
rect -13500 26095 -13498 26115
rect -13356 26095 -13354 26115
rect -13284 26095 -13282 26115
rect -13068 26095 -13066 26115
rect -12828 26095 -12826 26115
rect -12780 26095 -12778 26115
rect -12660 26095 -12658 26115
rect -12564 26095 -12562 26115
rect -12492 26095 -12490 26115
rect -12396 26095 -12394 26115
rect -12348 26095 -12346 26115
rect -12276 26095 -12274 26115
rect -12252 26095 -12250 26115
rect -12156 26095 -12154 26115
rect -12060 26095 -12058 26115
rect -11892 26112 -11890 26115
rect -11892 26095 -11889 26112
rect -11844 26095 -11842 26115
rect -11796 26095 -11794 26115
rect -11676 26095 -11674 26115
rect -11580 26095 -11578 26115
rect -11556 26095 -11554 26115
rect -11508 26095 -11506 26115
rect -11460 26095 -11458 26115
rect -11436 26095 -11434 26115
rect -11364 26095 -11362 26115
rect -11340 26095 -11338 26115
rect -11292 26095 -11290 26115
rect -11196 26095 -11194 26115
rect -11124 26095 -11122 26115
rect -11121 26112 -11107 26115
rect -11100 26115 -11011 26119
rect -11100 26112 -11083 26115
rect -11100 26095 -11098 26112
rect -11028 26095 -11026 26115
rect -11025 26112 -11011 26115
rect -11004 26115 77 26119
rect -11004 26112 -10987 26115
rect -11004 26095 -11002 26112
rect -10788 26095 -10786 26115
rect -10740 26095 -10738 26115
rect -10668 26095 -10666 26115
rect -10644 26095 -10642 26115
rect -9996 26095 -9994 26115
rect -9708 26095 -9706 26115
rect -9612 26095 -9610 26115
rect -9516 26095 -9514 26115
rect -9468 26095 -9466 26115
rect -9420 26095 -9418 26115
rect -9396 26095 -9394 26115
rect -9372 26095 -9370 26115
rect -9300 26095 -9298 26115
rect -9252 26095 -9250 26115
rect -9132 26096 -9130 26115
rect -9143 26095 -9109 26096
rect -9084 26095 -9082 26115
rect -9036 26095 -9034 26115
rect -8988 26095 -8986 26115
rect -8940 26095 -8938 26115
rect -8892 26095 -8890 26115
rect -8772 26095 -8770 26115
rect -8604 26095 -8602 26115
rect -8508 26096 -8506 26115
rect -8543 26095 -8485 26096
rect -8484 26095 -8482 26115
rect -8388 26095 -8386 26115
rect -8364 26095 -8362 26115
rect -8340 26095 -8338 26115
rect -8268 26095 -8266 26115
rect -8100 26095 -8098 26115
rect -8052 26095 -8050 26115
rect -7932 26095 -7930 26115
rect -7692 26095 -7690 26115
rect -7620 26095 -7618 26115
rect -7524 26095 -7522 26115
rect -7356 26095 -7354 26115
rect -7308 26095 -7306 26115
rect -7212 26095 -7210 26115
rect -7188 26095 -7186 26115
rect -7116 26095 -7114 26115
rect -7068 26095 -7066 26115
rect -6972 26095 -6970 26115
rect -6948 26095 -6946 26115
rect -6876 26095 -6874 26115
rect -6852 26095 -6850 26115
rect -6780 26095 -6778 26115
rect -6756 26095 -6754 26115
rect -6660 26095 -6658 26115
rect -6612 26095 -6610 26115
rect -6516 26095 -6514 26115
rect -6492 26095 -6490 26115
rect -6420 26095 -6418 26115
rect -6396 26095 -6394 26115
rect -6372 26095 -6370 26115
rect -6324 26095 -6322 26115
rect -6311 26110 -6308 26115
rect -6300 26110 -6298 26115
rect -6301 26096 -6298 26110
rect -6156 26095 -6154 26115
rect -6060 26095 -6058 26115
rect -5940 26095 -5938 26115
rect -5892 26095 -5890 26115
rect -5652 26095 -5650 26115
rect -5268 26095 -5266 26115
rect -5196 26095 -5194 26115
rect -5172 26095 -5170 26115
rect -5100 26095 -5098 26115
rect -5076 26095 -5074 26115
rect -4980 26095 -4978 26115
rect -4956 26095 -4954 26115
rect -4884 26095 -4882 26115
rect -4860 26095 -4858 26115
rect -4788 26095 -4786 26115
rect -4692 26095 -4690 26115
rect -4644 26095 -4642 26115
rect -4596 26095 -4594 26115
rect -4548 26095 -4546 26115
rect -4308 26095 -4306 26115
rect -4260 26095 -4258 26115
rect -4212 26095 -4210 26115
rect -4164 26095 -4162 26115
rect -4116 26095 -4114 26115
rect -4020 26095 -4018 26115
rect -3876 26095 -3874 26115
rect -3732 26095 -3730 26115
rect -3588 26095 -3586 26115
rect -3564 26095 -3562 26115
rect -3516 26095 -3514 26115
rect -3492 26095 -3490 26115
rect -3468 26095 -3466 26115
rect -3420 26095 -3418 26115
rect -3324 26095 -3322 26115
rect -3252 26095 -3250 26115
rect -3228 26095 -3226 26115
rect -3156 26095 -3154 26115
rect -3132 26095 -3130 26115
rect -3060 26095 -3058 26115
rect -3012 26095 -3010 26115
rect -2964 26095 -2962 26115
rect -2916 26095 -2914 26115
rect -2892 26095 -2890 26115
rect -2820 26095 -2818 26115
rect -2796 26095 -2794 26115
rect -2759 26110 -2756 26115
rect -2748 26110 -2746 26115
rect -2749 26096 -2746 26110
rect -2700 26095 -2698 26115
rect -2676 26095 -2673 26112
rect -2604 26095 -2602 26115
rect -2580 26095 -2578 26115
rect -2364 26095 -2362 26115
rect -2268 26095 -2266 26115
rect -2244 26095 -2242 26115
rect -2172 26095 -2170 26115
rect -2148 26095 -2146 26115
rect -2076 26095 -2074 26115
rect -2052 26095 -2050 26115
rect -1980 26095 -1978 26115
rect -1884 26095 -1882 26115
rect -1836 26095 -1834 26115
rect -1716 26095 -1714 26115
rect -1596 26095 -1594 26115
rect -1572 26095 -1570 26115
rect -1476 26095 -1474 26115
rect -1380 26095 -1378 26115
rect -1356 26095 -1354 26115
rect -1308 26095 -1306 26115
rect -1260 26095 -1258 26115
rect -1140 26095 -1138 26115
rect -852 26095 -850 26115
rect -804 26095 -802 26115
rect -756 26095 -754 26115
rect -708 26095 -706 26115
rect -612 26095 -610 26115
rect -588 26095 -586 26115
rect -540 26095 -538 26115
rect -492 26095 -490 26115
rect -444 26095 -442 26115
rect -396 26095 -394 26115
rect -300 26095 -298 26115
rect -276 26095 -274 26115
rect -228 26095 -226 26115
rect -12 26095 -10 26115
rect 63 26112 77 26115
rect 87 26115 3653 26119
rect 87 26112 101 26115
rect 108 26112 111 26115
rect 156 26095 158 26115
rect 204 26095 206 26115
rect 228 26095 230 26115
rect 252 26095 254 26115
rect 348 26095 350 26115
rect 468 26095 470 26115
rect 492 26095 494 26115
rect 564 26095 566 26115
rect 588 26095 590 26115
rect 636 26095 638 26115
rect 660 26095 662 26115
rect 732 26095 734 26115
rect 756 26095 758 26115
rect 841 26110 844 26115
rect 865 26110 868 26115
rect 876 26110 878 26115
rect 851 26096 854 26110
rect 875 26096 878 26110
rect 972 26112 974 26115
rect 852 26095 854 26096
rect 972 26095 975 26112
rect 1020 26095 1022 26115
rect 1068 26095 1070 26115
rect 1092 26095 1094 26115
rect 1116 26095 1118 26115
rect 1164 26095 1166 26115
rect 1212 26095 1214 26115
rect 1308 26095 1310 26115
rect 1332 26095 1334 26115
rect 1380 26095 1382 26115
rect 1428 26095 1430 26115
rect 1465 26110 1468 26115
rect 1475 26096 1478 26110
rect 1476 26095 1478 26096
rect 1524 26095 1526 26115
rect 1548 26095 1550 26115
rect 1596 26112 1598 26115
rect 1596 26095 1599 26112
rect 1620 26095 1622 26115
rect 1644 26095 1646 26115
rect 1692 26095 1694 26115
rect 1716 26095 1718 26115
rect 1740 26095 1742 26115
rect 1788 26095 1790 26115
rect 1884 26095 1886 26115
rect 1980 26095 1982 26115
rect 2028 26095 2030 26115
rect 2076 26095 2078 26115
rect 2100 26095 2102 26115
rect 2124 26095 2126 26115
rect 2172 26095 2174 26115
rect 2196 26095 2198 26115
rect 2220 26095 2222 26115
rect 2268 26095 2270 26115
rect 2292 26095 2294 26115
rect 2316 26095 2318 26115
rect 2364 26095 2366 26115
rect 2412 26095 2414 26115
rect 2460 26095 2462 26115
rect 2508 26095 2510 26115
rect 2580 26095 2582 26115
rect 2604 26095 2606 26115
rect 2676 26095 2678 26115
rect 2700 26095 2702 26115
rect 2748 26095 2750 26115
rect 2772 26095 2774 26115
rect 2796 26095 2798 26115
rect 2844 26095 2846 26115
rect 2868 26095 2870 26115
rect 2892 26095 2894 26115
rect 2940 26095 2942 26115
rect 3012 26095 3014 26115
rect 3108 26095 3110 26115
rect 3156 26095 3158 26115
rect 3252 26095 3254 26115
rect 3348 26095 3350 26115
rect 3396 26095 3398 26115
rect 3468 26095 3470 26115
rect 3492 26095 3494 26115
rect 3564 26095 3566 26115
rect 3612 26095 3614 26115
rect 3636 26095 3638 26115
rect 3639 26112 3653 26115
rect 3660 26115 23117 26119
rect 3660 26112 3677 26115
rect 3660 26095 3662 26112
rect 3708 26095 3710 26115
rect 3732 26095 3734 26115
rect 3804 26095 3806 26115
rect 3828 26095 3830 26115
rect 3924 26095 3926 26115
rect 4020 26095 4022 26115
rect 4044 26095 4046 26115
rect 4092 26095 4094 26115
rect 4116 26095 4118 26115
rect 4140 26095 4142 26115
rect 4188 26095 4190 26115
rect 4212 26095 4214 26115
rect 4236 26095 4238 26115
rect 4308 26095 4310 26115
rect 4332 26095 4334 26115
rect 4404 26095 4406 26115
rect 4500 26095 4502 26115
rect 4596 26095 4598 26115
rect 4860 26095 4862 26115
rect 4956 26095 4958 26115
rect 4980 26095 4982 26115
rect 5004 26095 5006 26115
rect 5076 26095 5078 26115
rect 5100 26095 5102 26115
rect 5124 26095 5126 26115
rect 5172 26095 5174 26115
rect 5220 26095 5222 26115
rect 5268 26095 5270 26115
rect 5388 26095 5390 26115
rect 5484 26095 5486 26115
rect 5508 26095 5510 26115
rect 5532 26095 5534 26115
rect 5628 26095 5630 26115
rect 5652 26095 5654 26115
rect 5748 26095 5750 26115
rect 5796 26095 5798 26115
rect 5844 26095 5846 26115
rect 5892 26095 5894 26115
rect 6132 26095 6134 26115
rect 6180 26095 6182 26115
rect 6228 26095 6230 26115
rect 6252 26095 6254 26115
rect 6276 26095 6278 26115
rect 6324 26095 6326 26115
rect 6372 26095 6374 26115
rect 6492 26095 6494 26115
rect 6588 26095 6590 26115
rect 6612 26095 6614 26115
rect 6660 26095 6662 26115
rect 6684 26095 6686 26115
rect 6708 26095 6710 26115
rect 6780 26095 6782 26115
rect 6804 26095 6806 26115
rect 6828 26095 6830 26115
rect 6900 26095 6902 26115
rect 6924 26095 6926 26115
rect 7020 26095 7022 26115
rect 7140 26095 7142 26115
rect 7236 26095 7238 26115
rect 7332 26095 7334 26115
rect 7380 26095 7382 26115
rect 7428 26095 7430 26115
rect 7452 26095 7454 26115
rect 7476 26095 7478 26115
rect 7524 26095 7526 26115
rect 7548 26095 7550 26115
rect 7572 26095 7574 26115
rect 7620 26095 7622 26115
rect 7644 26095 7646 26115
rect 7668 26095 7670 26115
rect 7716 26096 7718 26115
rect 7681 26095 7739 26096
rect 7740 26095 7742 26115
rect 7836 26095 7838 26115
rect 7884 26095 7886 26115
rect 7932 26095 7934 26115
rect 7956 26095 7958 26115
rect 7980 26095 7982 26115
rect 8028 26095 8030 26115
rect 8196 26095 8198 26115
rect 8244 26095 8246 26115
rect 8268 26095 8270 26115
rect 8292 26095 8294 26115
rect 8340 26095 8342 26115
rect 8364 26095 8366 26115
rect 8388 26095 8390 26115
rect 8436 26095 8438 26115
rect 8460 26095 8462 26115
rect 8556 26095 8558 26115
rect 8604 26095 8606 26115
rect 8652 26095 8654 26115
rect 8700 26095 8702 26115
rect 8724 26095 8726 26115
rect 8748 26095 8750 26115
rect 8820 26095 8822 26115
rect 8844 26095 8846 26115
rect 8868 26095 8870 26115
rect 9516 26095 9518 26115
rect 9612 26095 9614 26115
rect 9660 26095 9662 26115
rect 9684 26095 9686 26115
rect 9708 26095 9710 26115
rect 9756 26095 9758 26115
rect 9780 26095 9782 26115
rect 9804 26095 9806 26115
rect 9852 26095 9854 26115
rect 9876 26095 9878 26115
rect 9900 26095 9902 26115
rect 9948 26095 9950 26115
rect 9972 26095 9974 26115
rect 9996 26095 9998 26115
rect 10068 26095 10070 26115
rect 10092 26095 10094 26115
rect 10116 26095 10118 26115
rect 10164 26095 10166 26115
rect 10188 26095 10190 26115
rect 10212 26095 10214 26115
rect 10284 26095 10286 26115
rect 10308 26095 10310 26115
rect 10332 26095 10334 26115
rect 10380 26095 10382 26115
rect 10404 26095 10406 26115
rect 10428 26095 10430 26115
rect 10476 26095 10478 26115
rect 10500 26095 10502 26115
rect 10524 26095 10526 26115
rect 10572 26095 10574 26115
rect 10596 26095 10598 26115
rect 10620 26095 10622 26115
rect 10668 26095 10670 26115
rect 10692 26095 10694 26115
rect 10716 26095 10718 26115
rect 10788 26095 10790 26115
rect 10836 26095 10838 26115
rect 10956 26095 10958 26115
rect 11052 26095 11054 26115
rect 11076 26095 11078 26115
rect 11124 26095 11126 26115
rect 11172 26095 11174 26115
rect 11220 26095 11222 26115
rect 11340 26095 11342 26115
rect 11436 26095 11438 26115
rect 11532 26095 11534 26115
rect 11580 26095 11582 26115
rect 11628 26095 11630 26115
rect 11676 26095 11678 26115
rect 11724 26095 11726 26115
rect 11772 26095 11774 26115
rect 11796 26095 11798 26115
rect 11892 26095 11894 26115
rect 11988 26095 11990 26115
rect 12060 26095 12062 26115
rect 12132 26095 12134 26115
rect 12228 26095 12230 26115
rect 12276 26095 12278 26115
rect 12324 26095 12326 26115
rect 12420 26095 12422 26115
rect 12444 26095 12446 26115
rect 12492 26095 12494 26115
rect 12516 26095 12518 26115
rect 12540 26095 12542 26115
rect 12588 26095 12590 26115
rect 12636 26095 12638 26115
rect 12732 26095 12734 26115
rect 12756 26095 12758 26115
rect 12804 26095 12806 26115
rect 12828 26095 12830 26115
rect 12852 26095 12854 26115
rect 12900 26095 12902 26115
rect 12948 26095 12950 26115
rect 13044 26095 13046 26115
rect 13068 26095 13070 26115
rect 13116 26095 13118 26115
rect 13284 26095 13286 26115
rect 13332 26095 13334 26115
rect 13428 26095 13430 26115
rect 13524 26095 13526 26115
rect 13572 26095 13574 26115
rect 13644 26095 13646 26115
rect 13668 26095 13670 26115
rect 13764 26095 13766 26115
rect 13812 26095 13814 26115
rect 13860 26095 13862 26115
rect 13908 26095 13910 26115
rect 13956 26095 13958 26115
rect 14004 26095 14006 26115
rect 14100 26095 14102 26115
rect 14196 26095 14198 26115
rect 14292 26095 14294 26115
rect 15132 26095 15134 26115
rect 15180 26095 15182 26115
rect 15228 26095 15230 26115
rect 15252 26095 15254 26115
rect 15324 26095 15326 26115
rect 15396 26095 15398 26115
rect 15420 26095 15422 26115
rect 15492 26095 15494 26115
rect 15540 26095 15542 26115
rect 15636 26095 15638 26115
rect 15660 26095 15662 26115
rect 15708 26095 15710 26115
rect 15732 26095 15734 26115
rect 15756 26095 15758 26115
rect 15804 26095 15806 26115
rect 15828 26095 15830 26115
rect 15852 26095 15854 26115
rect 15900 26095 15902 26115
rect 15948 26095 15950 26115
rect 15996 26095 15998 26115
rect 16044 26095 16046 26115
rect 16092 26095 16094 26115
rect 16260 26095 16262 26115
rect 16308 26095 16310 26115
rect 16332 26095 16334 26115
rect 16356 26095 16358 26115
rect 16404 26095 16406 26115
rect 16452 26095 16454 26115
rect 16548 26095 16550 26115
rect 16572 26095 16574 26115
rect 16620 26095 16622 26115
rect 16668 26095 16670 26115
rect 16716 26095 16718 26115
rect 16764 26095 16766 26115
rect 16812 26095 16814 26115
rect 16884 26095 16886 26115
rect 16908 26095 16910 26115
rect 16980 26095 16982 26115
rect 17052 26095 17054 26115
rect 17196 26095 17198 26115
rect 17220 26095 17222 26115
rect 17292 26095 17294 26115
rect 17316 26095 17318 26115
rect 18084 26095 18086 26115
rect 18132 26095 18134 26115
rect 18396 26095 18398 26115
rect 18492 26095 18494 26115
rect 18516 26095 18518 26115
rect 18564 26095 18566 26115
rect 18612 26095 18614 26115
rect 18660 26095 18662 26115
rect 18708 26095 18710 26115
rect 18756 26095 18758 26115
rect 18804 26095 18806 26115
rect 18852 26095 18854 26115
rect 18900 26095 18902 26115
rect 18996 26095 18998 26115
rect 19020 26095 19022 26115
rect 19092 26095 19094 26115
rect 19116 26095 19118 26115
rect 19140 26095 19142 26115
rect 19188 26095 19190 26115
rect 19236 26095 19238 26115
rect 19332 26095 19334 26115
rect 19476 26095 19478 26115
rect 19620 26095 19622 26115
rect 19716 26095 19718 26115
rect 19788 26095 19790 26115
rect 19836 26095 19838 26115
rect 19860 26095 19862 26115
rect 19884 26095 19886 26115
rect 19932 26095 19934 26115
rect 19956 26095 19958 26115
rect 19980 26095 19982 26115
rect 20028 26095 20030 26115
rect 20052 26095 20054 26115
rect 20076 26095 20078 26115
rect 20148 26095 20150 26115
rect 20172 26095 20174 26115
rect 20196 26095 20198 26115
rect 20268 26095 20270 26115
rect 20292 26095 20294 26115
rect 20388 26095 20390 26115
rect 20412 26095 20414 26115
rect 20508 26095 20510 26115
rect 20556 26095 20558 26115
rect 20604 26095 20606 26115
rect 20916 26095 20918 26115
rect 20964 26095 20966 26115
rect 21012 26095 21014 26115
rect 21060 26095 21062 26115
rect 21084 26095 21086 26115
rect 21108 26095 21110 26115
rect 21204 26095 21206 26115
rect 21300 26095 21302 26115
rect 21324 26095 21326 26115
rect 21444 26095 21446 26115
rect 21468 26095 21470 26115
rect 21564 26095 21566 26115
rect 21612 26095 21614 26115
rect 21684 26095 21686 26115
rect 21708 26095 21710 26115
rect 21828 26095 21830 26115
rect 21924 26095 21926 26115
rect 22068 26095 22070 26115
rect 22188 26095 22190 26115
rect 22212 26095 22214 26115
rect 22884 26095 22886 26115
rect 22980 26095 22982 26115
rect 23076 26095 23078 26115
rect 23100 26095 23102 26115
rect 23103 26112 23117 26115
rect 23124 26115 25157 26119
rect 23124 26112 23141 26115
rect 23148 26112 23151 26115
rect 23124 26095 23126 26112
rect 23244 26095 23246 26115
rect 23340 26095 23342 26115
rect 23412 26095 23414 26115
rect 23556 26095 23558 26115
rect 23628 26095 23630 26115
rect 23652 26095 23654 26115
rect 23676 26095 23678 26115
rect 23724 26095 23726 26115
rect 23772 26095 23774 26115
rect 23820 26095 23822 26115
rect 23868 26095 23870 26115
rect 23916 26095 23918 26115
rect 24012 26095 24014 26115
rect 24084 26095 24086 26115
rect 24217 26095 24251 26096
rect 24396 26095 24398 26115
rect 24492 26095 24494 26115
rect 24516 26095 24518 26115
rect 24588 26095 24590 26115
rect 24612 26095 24614 26115
rect 24708 26095 24710 26115
rect 24732 26095 24734 26115
rect 24756 26095 24758 26115
rect 24852 26095 24854 26115
rect 24876 26095 24878 26115
rect 24972 26095 24974 26115
rect 24996 26095 24998 26115
rect 25068 26095 25070 26115
rect 25143 26112 25157 26115
rect 25164 26115 30803 26119
rect 25164 26112 25181 26115
rect 25164 26095 25166 26112
rect 25260 26095 25262 26115
rect 25308 26095 25310 26115
rect 25356 26095 25358 26115
rect 25380 26095 25382 26115
rect 25404 26095 25406 26115
rect 25452 26095 25454 26115
rect 25500 26095 25502 26115
rect 25596 26095 25598 26115
rect 27108 26095 27110 26115
rect 27324 26095 27326 26115
rect 27396 26095 27398 26115
rect 27420 26095 27422 26115
rect 27540 26095 27542 26115
rect 27564 26095 27566 26115
rect 30564 26095 30566 26115
rect 30660 26095 30662 26115
rect 30769 26110 30772 26115
rect 30780 26110 30782 26115
rect 30779 26096 30782 26110
rect 30697 26095 30731 26096
rect -16641 26091 -2683 26095
rect -16641 26088 -16627 26091
rect -16620 26088 -16617 26091
rect -16679 26086 -16676 26088
rect -16668 26086 -16666 26088
rect -16669 26072 -16666 26086
rect -16380 26071 -16378 26091
rect -16356 26071 -16354 26091
rect -16284 26071 -16282 26091
rect -16260 26071 -16258 26091
rect -16236 26071 -16234 26091
rect -15324 26071 -15322 26091
rect -15084 26071 -15082 26091
rect -14868 26071 -14866 26091
rect -14772 26071 -14770 26091
rect -14724 26071 -14722 26091
rect -14508 26071 -14506 26091
rect -14436 26071 -14434 26091
rect -14340 26071 -14338 26091
rect -14244 26071 -14242 26091
rect -14172 26072 -14170 26091
rect -14207 26071 -14149 26072
rect -14076 26071 -14074 26091
rect -13980 26071 -13978 26091
rect -13932 26071 -13930 26091
rect -13884 26071 -13882 26091
rect -13788 26071 -13786 26091
rect -13655 26086 -13652 26091
rect -13644 26086 -13642 26091
rect -13645 26072 -13642 26086
rect -13572 26071 -13569 26088
rect -13500 26071 -13498 26091
rect -13356 26071 -13354 26091
rect -13284 26071 -13282 26091
rect -13161 26088 -13147 26091
rect -13068 26071 -13066 26091
rect -12828 26071 -12826 26091
rect -12780 26071 -12778 26091
rect -12660 26071 -12658 26091
rect -12564 26071 -12562 26091
rect -12492 26071 -12490 26091
rect -12396 26071 -12394 26091
rect -12348 26071 -12346 26091
rect -12276 26071 -12274 26091
rect -12252 26071 -12250 26091
rect -12156 26071 -12154 26091
rect -12060 26071 -12058 26091
rect -11913 26088 -11899 26091
rect -11892 26088 -11889 26091
rect -11844 26071 -11842 26091
rect -11796 26071 -11794 26091
rect -11676 26071 -11674 26091
rect -11580 26071 -11578 26091
rect -11556 26071 -11554 26091
rect -11508 26071 -11506 26091
rect -11460 26071 -11458 26091
rect -11436 26071 -11434 26091
rect -11364 26071 -11362 26091
rect -11340 26071 -11338 26091
rect -11292 26071 -11290 26091
rect -11196 26071 -11194 26091
rect -11124 26071 -11122 26091
rect -11100 26071 -11098 26091
rect -11028 26071 -11026 26091
rect -11004 26071 -11002 26091
rect -10788 26071 -10786 26091
rect -10740 26071 -10738 26091
rect -10668 26071 -10666 26091
rect -10644 26071 -10642 26091
rect -9996 26071 -9994 26091
rect -9708 26071 -9706 26091
rect -9612 26071 -9610 26091
rect -9516 26071 -9514 26091
rect -9468 26071 -9466 26091
rect -9420 26071 -9418 26091
rect -9396 26071 -9394 26091
rect -9372 26071 -9370 26091
rect -9300 26071 -9298 26091
rect -9252 26071 -9250 26091
rect -9143 26086 -9140 26091
rect -9132 26086 -9130 26091
rect -9133 26072 -9130 26086
rect -9084 26071 -9082 26091
rect -9036 26088 -9034 26091
rect -9036 26071 -9033 26088
rect -8988 26071 -8986 26091
rect -8940 26071 -8938 26091
rect -8892 26071 -8890 26091
rect -8772 26071 -8770 26091
rect -8604 26071 -8602 26091
rect -8519 26086 -8516 26091
rect -8508 26086 -8506 26091
rect -8509 26072 -8506 26086
rect -8484 26071 -8482 26091
rect -8436 26071 -8433 26088
rect -8388 26071 -8386 26091
rect -8364 26071 -8362 26091
rect -8340 26071 -8338 26091
rect -8268 26071 -8266 26091
rect -8100 26071 -8098 26091
rect -8052 26071 -8050 26091
rect -7932 26071 -7930 26091
rect -7692 26071 -7690 26091
rect -7620 26071 -7618 26091
rect -7524 26071 -7522 26091
rect -7356 26071 -7354 26091
rect -7308 26071 -7306 26091
rect -7212 26071 -7210 26091
rect -7188 26071 -7186 26091
rect -7116 26071 -7114 26091
rect -7068 26071 -7066 26091
rect -6972 26071 -6970 26091
rect -6948 26071 -6946 26091
rect -6876 26071 -6874 26091
rect -6852 26071 -6850 26091
rect -6780 26071 -6778 26091
rect -6756 26071 -6754 26091
rect -6660 26071 -6658 26091
rect -6612 26071 -6610 26091
rect -6516 26071 -6514 26091
rect -6492 26071 -6490 26091
rect -6420 26071 -6418 26091
rect -6396 26071 -6394 26091
rect -6372 26071 -6370 26091
rect -6324 26071 -6322 26091
rect -6225 26088 -6211 26091
rect -6156 26071 -6154 26091
rect -6060 26071 -6058 26091
rect -5940 26071 -5938 26091
rect -5892 26071 -5890 26091
rect -5652 26071 -5650 26091
rect -5268 26071 -5266 26091
rect -5196 26071 -5194 26091
rect -5172 26071 -5170 26091
rect -5100 26071 -5098 26091
rect -5076 26071 -5074 26091
rect -4980 26071 -4978 26091
rect -4956 26071 -4954 26091
rect -4884 26071 -4882 26091
rect -4860 26071 -4858 26091
rect -4788 26071 -4786 26091
rect -4692 26071 -4690 26091
rect -4644 26071 -4642 26091
rect -4596 26071 -4594 26091
rect -4593 26088 -4579 26091
rect -4548 26071 -4546 26091
rect -4308 26071 -4306 26091
rect -4260 26071 -4258 26091
rect -4212 26071 -4210 26091
rect -4164 26071 -4162 26091
rect -4116 26071 -4114 26091
rect -4020 26071 -4018 26091
rect -3876 26071 -3874 26091
rect -3732 26071 -3730 26091
rect -3588 26071 -3586 26091
rect -3564 26071 -3562 26091
rect -3516 26071 -3514 26091
rect -3492 26071 -3490 26091
rect -3468 26071 -3466 26091
rect -3420 26071 -3418 26091
rect -3324 26071 -3322 26091
rect -3252 26071 -3250 26091
rect -3228 26071 -3226 26091
rect -3156 26071 -3154 26091
rect -3132 26071 -3130 26091
rect -3060 26071 -3058 26091
rect -3012 26071 -3010 26091
rect -2964 26071 -2962 26091
rect -2916 26071 -2914 26091
rect -2892 26071 -2890 26091
rect -2879 26071 -2821 26072
rect -2820 26071 -2818 26091
rect -2796 26071 -2794 26091
rect -2700 26071 -2698 26091
rect -2697 26088 -2683 26091
rect -2676 26091 941 26095
rect -2676 26088 -2659 26091
rect -2676 26071 -2674 26088
rect -2604 26071 -2602 26091
rect -2580 26071 -2578 26091
rect -2364 26071 -2362 26091
rect -2268 26071 -2266 26091
rect -2244 26071 -2242 26091
rect -2172 26071 -2170 26091
rect -2148 26071 -2146 26091
rect -2076 26071 -2074 26091
rect -2052 26071 -2050 26091
rect -1980 26071 -1978 26091
rect -1884 26071 -1882 26091
rect -1836 26071 -1834 26091
rect -1716 26071 -1714 26091
rect -1596 26071 -1594 26091
rect -1572 26071 -1570 26091
rect -1476 26071 -1474 26091
rect -1380 26071 -1378 26091
rect -1356 26071 -1354 26091
rect -1308 26071 -1306 26091
rect -1260 26071 -1258 26091
rect -1140 26071 -1138 26091
rect -911 26071 -877 26072
rect -852 26071 -850 26091
rect -804 26071 -802 26091
rect -756 26071 -754 26091
rect -708 26071 -706 26091
rect -612 26071 -610 26091
rect -588 26071 -586 26091
rect -540 26071 -538 26091
rect -492 26071 -490 26091
rect -444 26071 -442 26091
rect -396 26071 -394 26091
rect -300 26071 -298 26091
rect -276 26071 -274 26091
rect -228 26071 -226 26091
rect -12 26071 -10 26091
rect 156 26071 158 26091
rect 204 26071 206 26091
rect 228 26071 230 26091
rect 252 26071 254 26091
rect 348 26071 350 26091
rect 468 26071 470 26091
rect 492 26071 494 26091
rect 564 26071 566 26091
rect 588 26071 590 26091
rect 636 26071 638 26091
rect 660 26071 662 26091
rect 732 26071 734 26091
rect 756 26071 758 26091
rect 852 26071 854 26091
rect 927 26088 941 26091
rect 951 26091 1565 26095
rect 951 26088 965 26091
rect 972 26088 975 26091
rect 1020 26071 1022 26091
rect 1068 26072 1070 26091
rect 1033 26071 1091 26072
rect 1092 26071 1094 26091
rect 1116 26071 1118 26091
rect 1164 26071 1166 26091
rect 1212 26071 1214 26091
rect 1308 26071 1310 26091
rect 1332 26071 1334 26091
rect 1380 26071 1382 26091
rect 1428 26071 1430 26091
rect 1476 26071 1478 26091
rect 1524 26071 1526 26091
rect 1548 26071 1550 26091
rect 1551 26088 1565 26091
rect 1575 26091 30731 26095
rect 1575 26088 1589 26091
rect 1596 26088 1599 26091
rect 1620 26071 1622 26091
rect 1644 26071 1646 26091
rect 1692 26071 1694 26091
rect 1716 26071 1718 26091
rect 1740 26071 1742 26091
rect 1788 26071 1790 26091
rect 1884 26071 1886 26091
rect 1980 26071 1982 26091
rect 2028 26071 2030 26091
rect 2076 26071 2078 26091
rect 2100 26071 2102 26091
rect 2124 26071 2126 26091
rect 2172 26071 2174 26091
rect 2196 26071 2198 26091
rect 2220 26071 2222 26091
rect 2268 26071 2270 26091
rect 2292 26071 2294 26091
rect 2316 26071 2318 26091
rect 2364 26071 2366 26091
rect 2412 26071 2414 26091
rect 2460 26071 2462 26091
rect 2508 26071 2510 26091
rect 2580 26071 2582 26091
rect 2604 26071 2606 26091
rect 2676 26071 2678 26091
rect 2700 26071 2702 26091
rect 2748 26071 2750 26091
rect 2772 26071 2774 26091
rect 2796 26071 2798 26091
rect 2844 26071 2846 26091
rect 2868 26071 2870 26091
rect 2892 26071 2894 26091
rect 2940 26071 2942 26091
rect 3012 26071 3014 26091
rect 3108 26071 3110 26091
rect 3156 26071 3158 26091
rect 3252 26071 3254 26091
rect 3348 26071 3350 26091
rect 3396 26071 3398 26091
rect 3468 26071 3470 26091
rect 3492 26071 3494 26091
rect 3564 26071 3566 26091
rect 3612 26071 3614 26091
rect 3636 26071 3638 26091
rect 3660 26071 3662 26091
rect 3708 26071 3710 26091
rect 3732 26071 3734 26091
rect 3804 26071 3806 26091
rect 3828 26071 3830 26091
rect 3924 26071 3926 26091
rect 4020 26071 4022 26091
rect 4044 26071 4046 26091
rect 4092 26071 4094 26091
rect 4116 26071 4118 26091
rect 4140 26071 4142 26091
rect 4188 26071 4190 26091
rect 4212 26071 4214 26091
rect 4236 26071 4238 26091
rect 4308 26071 4310 26091
rect 4332 26071 4334 26091
rect 4404 26071 4406 26091
rect 4500 26071 4502 26091
rect 4596 26071 4598 26091
rect 4860 26071 4862 26091
rect 4956 26071 4958 26091
rect 4980 26071 4982 26091
rect 5004 26071 5006 26091
rect 5076 26071 5078 26091
rect 5100 26071 5102 26091
rect 5124 26071 5126 26091
rect 5172 26071 5174 26091
rect 5220 26071 5222 26091
rect 5268 26071 5270 26091
rect 5388 26071 5390 26091
rect 5484 26071 5486 26091
rect 5508 26071 5510 26091
rect 5532 26071 5534 26091
rect 5628 26071 5630 26091
rect 5652 26071 5654 26091
rect 5748 26071 5750 26091
rect 5796 26071 5798 26091
rect 5844 26071 5846 26091
rect 5892 26071 5894 26091
rect 6132 26071 6134 26091
rect 6180 26071 6182 26091
rect 6228 26071 6230 26091
rect 6252 26071 6254 26091
rect 6276 26071 6278 26091
rect 6324 26071 6326 26091
rect 6372 26071 6374 26091
rect 6492 26071 6494 26091
rect 6588 26071 6590 26091
rect 6612 26071 6614 26091
rect 6660 26071 6662 26091
rect 6684 26071 6686 26091
rect 6708 26071 6710 26091
rect 6780 26071 6782 26091
rect 6804 26071 6806 26091
rect 6828 26071 6830 26091
rect 6900 26071 6902 26091
rect 6924 26071 6926 26091
rect 7020 26071 7022 26091
rect 7140 26071 7142 26091
rect 7236 26071 7238 26091
rect 7332 26071 7334 26091
rect 7380 26071 7382 26091
rect 7428 26071 7430 26091
rect 7452 26071 7454 26091
rect 7476 26071 7478 26091
rect 7524 26071 7526 26091
rect 7548 26071 7550 26091
rect 7572 26071 7574 26091
rect 7620 26071 7622 26091
rect 7644 26071 7646 26091
rect 7668 26071 7670 26091
rect 7705 26086 7708 26091
rect 7716 26086 7718 26091
rect 7715 26072 7718 26086
rect 7740 26071 7742 26091
rect 7788 26071 7791 26088
rect 7836 26072 7838 26091
rect 7801 26071 7859 26072
rect 7884 26071 7886 26091
rect 7932 26071 7934 26091
rect 7956 26071 7958 26091
rect 7980 26071 7982 26091
rect 8028 26071 8030 26091
rect 8196 26071 8198 26091
rect 8244 26071 8246 26091
rect 8268 26071 8270 26091
rect 8292 26071 8294 26091
rect 8340 26071 8342 26091
rect 8364 26071 8366 26091
rect 8388 26071 8390 26091
rect 8436 26071 8438 26091
rect 8460 26071 8462 26091
rect 8556 26071 8558 26091
rect 8604 26071 8606 26091
rect 8652 26071 8654 26091
rect 8700 26071 8702 26091
rect 8724 26071 8726 26091
rect 8748 26071 8750 26091
rect 8820 26071 8822 26091
rect 8844 26071 8846 26091
rect 8868 26071 8870 26091
rect 9516 26071 9518 26091
rect 9612 26071 9614 26091
rect 9660 26071 9662 26091
rect 9684 26071 9686 26091
rect 9708 26071 9710 26091
rect 9756 26071 9758 26091
rect 9780 26071 9782 26091
rect 9804 26071 9806 26091
rect 9852 26071 9854 26091
rect 9876 26071 9878 26091
rect 9900 26071 9902 26091
rect 9948 26071 9950 26091
rect 9972 26071 9974 26091
rect 9996 26071 9998 26091
rect 10068 26071 10070 26091
rect 10092 26071 10094 26091
rect 10116 26071 10118 26091
rect 10164 26071 10166 26091
rect 10188 26071 10190 26091
rect 10212 26071 10214 26091
rect 10284 26071 10286 26091
rect 10308 26071 10310 26091
rect 10332 26071 10334 26091
rect 10380 26071 10382 26091
rect 10404 26071 10406 26091
rect 10428 26071 10430 26091
rect 10476 26071 10478 26091
rect 10500 26071 10502 26091
rect 10524 26071 10526 26091
rect 10572 26071 10574 26091
rect 10596 26071 10598 26091
rect 10620 26071 10622 26091
rect 10668 26071 10670 26091
rect 10692 26071 10694 26091
rect 10716 26071 10718 26091
rect 10788 26071 10790 26091
rect 10836 26071 10838 26091
rect 10956 26071 10958 26091
rect 11052 26071 11054 26091
rect 11076 26071 11078 26091
rect 11124 26071 11126 26091
rect 11172 26071 11174 26091
rect 11220 26071 11222 26091
rect 11340 26071 11342 26091
rect 11436 26071 11438 26091
rect 11532 26071 11534 26091
rect 11580 26071 11582 26091
rect 11628 26071 11630 26091
rect 11676 26071 11678 26091
rect 11724 26071 11726 26091
rect 11772 26071 11774 26091
rect 11796 26071 11798 26091
rect 11892 26071 11894 26091
rect 11988 26071 11990 26091
rect 12060 26071 12062 26091
rect 12132 26071 12134 26091
rect 12228 26071 12230 26091
rect 12276 26071 12278 26091
rect 12324 26071 12326 26091
rect 12420 26071 12422 26091
rect 12444 26071 12446 26091
rect 12492 26071 12494 26091
rect 12516 26071 12518 26091
rect 12540 26071 12542 26091
rect 12588 26071 12590 26091
rect 12636 26071 12638 26091
rect 12732 26071 12734 26091
rect 12756 26071 12758 26091
rect 12804 26071 12806 26091
rect 12828 26071 12830 26091
rect 12852 26071 12854 26091
rect 12900 26071 12902 26091
rect 12948 26071 12950 26091
rect 13044 26071 13046 26091
rect 13068 26071 13070 26091
rect 13116 26071 13118 26091
rect 13284 26071 13286 26091
rect 13332 26071 13334 26091
rect 13428 26071 13430 26091
rect 13524 26071 13526 26091
rect 13572 26071 13574 26091
rect 13644 26071 13646 26091
rect 13668 26071 13670 26091
rect 13764 26071 13766 26091
rect 13812 26071 13814 26091
rect 13860 26071 13862 26091
rect 13908 26071 13910 26091
rect 13956 26071 13958 26091
rect 14004 26071 14006 26091
rect 14100 26071 14102 26091
rect 14196 26071 14198 26091
rect 14292 26071 14294 26091
rect 15132 26071 15134 26091
rect 15180 26071 15182 26091
rect 15228 26071 15230 26091
rect 15252 26071 15254 26091
rect 15324 26071 15326 26091
rect 15396 26071 15398 26091
rect 15420 26071 15422 26091
rect 15492 26071 15494 26091
rect 15540 26071 15542 26091
rect 15636 26071 15638 26091
rect 15660 26071 15662 26091
rect 15708 26071 15710 26091
rect 15732 26071 15734 26091
rect 15756 26071 15758 26091
rect 15804 26071 15806 26091
rect 15828 26071 15830 26091
rect 15852 26071 15854 26091
rect 15900 26071 15902 26091
rect 15948 26071 15950 26091
rect 15996 26071 15998 26091
rect 16044 26071 16046 26091
rect 16092 26072 16094 26091
rect 16057 26071 16115 26072
rect 16260 26071 16262 26091
rect 16308 26071 16310 26091
rect 16332 26071 16334 26091
rect 16356 26071 16358 26091
rect 16404 26071 16406 26091
rect 16452 26071 16454 26091
rect 16548 26071 16550 26091
rect 16572 26071 16574 26091
rect 16620 26071 16622 26091
rect 16668 26071 16670 26091
rect 16716 26071 16718 26091
rect 16764 26071 16766 26091
rect 16812 26071 16814 26091
rect 16884 26071 16886 26091
rect 16908 26071 16910 26091
rect 16980 26071 16982 26091
rect 17052 26071 17054 26091
rect 17196 26071 17198 26091
rect 17220 26071 17222 26091
rect 17292 26071 17294 26091
rect 17316 26071 17318 26091
rect 18084 26071 18086 26091
rect 18132 26071 18134 26091
rect 18396 26071 18398 26091
rect 18492 26071 18494 26091
rect 18516 26071 18518 26091
rect 18564 26071 18566 26091
rect 18612 26071 18614 26091
rect 18660 26071 18662 26091
rect 18708 26071 18710 26091
rect 18756 26071 18758 26091
rect 18804 26071 18806 26091
rect 18852 26071 18854 26091
rect 18900 26071 18902 26091
rect 18996 26071 18998 26091
rect 19020 26071 19022 26091
rect 19092 26071 19094 26091
rect 19116 26071 19118 26091
rect 19140 26071 19142 26091
rect 19188 26071 19190 26091
rect 19236 26071 19238 26091
rect 19332 26071 19334 26091
rect 19476 26071 19478 26091
rect 19620 26072 19622 26091
rect 19609 26071 19643 26072
rect 19716 26071 19718 26091
rect 19788 26071 19790 26091
rect 19836 26071 19838 26091
rect 19860 26071 19862 26091
rect 19884 26071 19886 26091
rect 19932 26071 19934 26091
rect 19956 26071 19958 26091
rect 19980 26071 19982 26091
rect 20028 26071 20030 26091
rect 20052 26071 20054 26091
rect 20076 26071 20078 26091
rect 20148 26071 20150 26091
rect 20172 26071 20174 26091
rect 20196 26071 20198 26091
rect 20268 26071 20270 26091
rect 20292 26071 20294 26091
rect 20388 26071 20390 26091
rect 20412 26071 20414 26091
rect 20508 26071 20510 26091
rect 20556 26071 20558 26091
rect 20604 26071 20606 26091
rect 20916 26071 20918 26091
rect 20964 26071 20966 26091
rect 21012 26071 21014 26091
rect 21060 26071 21062 26091
rect 21084 26071 21086 26091
rect 21108 26071 21110 26091
rect 21204 26071 21206 26091
rect 21300 26071 21302 26091
rect 21324 26071 21326 26091
rect 21444 26071 21446 26091
rect 21468 26071 21470 26091
rect 21564 26071 21566 26091
rect 21612 26071 21614 26091
rect 21684 26071 21686 26091
rect 21708 26071 21710 26091
rect 21828 26071 21830 26091
rect 21924 26071 21926 26091
rect 22068 26071 22070 26091
rect 22188 26071 22190 26091
rect 22212 26071 22214 26091
rect 22884 26071 22886 26091
rect 22980 26071 22982 26091
rect 23076 26071 23078 26091
rect 23100 26071 23102 26091
rect 23124 26071 23126 26091
rect 23244 26071 23246 26091
rect 23340 26071 23342 26091
rect 23412 26071 23414 26091
rect 23556 26071 23558 26091
rect 23628 26071 23630 26091
rect 23652 26071 23654 26091
rect 23676 26071 23678 26091
rect 23724 26071 23726 26091
rect 23772 26071 23774 26091
rect 23820 26071 23822 26091
rect 23868 26071 23870 26091
rect 23916 26071 23918 26091
rect 24012 26071 24014 26091
rect 24084 26071 24086 26091
rect 24396 26071 24398 26091
rect 24492 26071 24494 26091
rect 24516 26071 24518 26091
rect 24588 26071 24590 26091
rect 24612 26071 24614 26091
rect 24708 26071 24710 26091
rect 24732 26071 24734 26091
rect 24756 26071 24758 26091
rect 24852 26071 24854 26091
rect 24876 26071 24878 26091
rect 24972 26071 24974 26091
rect 24996 26071 24998 26091
rect 25068 26071 25070 26091
rect 25164 26071 25166 26091
rect 25260 26071 25262 26091
rect 25308 26071 25310 26091
rect 25356 26071 25358 26091
rect 25380 26071 25382 26091
rect 25404 26071 25406 26091
rect 25452 26071 25454 26091
rect 25500 26071 25502 26091
rect 25596 26071 25598 26091
rect 27108 26071 27110 26091
rect 27324 26071 27326 26091
rect 27396 26071 27398 26091
rect 27420 26071 27422 26091
rect 27540 26071 27542 26091
rect 27564 26071 27566 26091
rect 30564 26071 30566 26091
rect 30660 26071 30662 26091
rect 30673 26071 30707 26072
rect -17481 26067 -16963 26071
rect -17481 26064 -17467 26067
rect -17460 26064 -17457 26067
rect -17388 26047 -17386 26067
rect -17303 26062 -17300 26067
rect -17292 26062 -17290 26067
rect -16977 26064 -16963 26067
rect -16953 26067 -16603 26071
rect -16953 26064 -16939 26067
rect -16932 26064 -16929 26067
rect -17293 26048 -17290 26062
rect -17052 26047 -17049 26064
rect -16895 26047 -16861 26048
rect -16836 26047 -16834 26067
rect -16764 26047 -16762 26067
rect -16740 26047 -16738 26067
rect -16617 26064 -16603 26067
rect -16593 26067 -13579 26071
rect -16593 26064 -16579 26067
rect -16380 26047 -16378 26067
rect -16356 26047 -16354 26067
rect -16284 26047 -16282 26067
rect -16260 26047 -16258 26067
rect -16236 26047 -16234 26067
rect -15324 26047 -15322 26067
rect -15084 26047 -15082 26067
rect -14868 26047 -14866 26067
rect -14772 26047 -14770 26067
rect -14724 26048 -14722 26067
rect -14735 26047 -14701 26048
rect -14508 26047 -14506 26067
rect -14436 26047 -14434 26067
rect -14340 26047 -14338 26067
rect -14244 26047 -14242 26067
rect -14183 26062 -14180 26067
rect -14172 26062 -14170 26067
rect -14173 26048 -14170 26062
rect -14076 26064 -14074 26067
rect -14076 26047 -14073 26064
rect -13980 26047 -13978 26067
rect -13932 26047 -13930 26067
rect -13884 26047 -13882 26067
rect -13788 26047 -13786 26067
rect -13593 26064 -13579 26067
rect -13572 26067 -8443 26071
rect -13572 26064 -13555 26067
rect -13572 26047 -13570 26064
rect -13500 26047 -13498 26067
rect -13356 26047 -13354 26067
rect -13284 26047 -13282 26067
rect -13068 26047 -13066 26067
rect -12828 26047 -12826 26067
rect -12780 26047 -12778 26067
rect -12660 26047 -12658 26067
rect -12564 26047 -12562 26067
rect -12492 26047 -12490 26067
rect -12396 26047 -12394 26067
rect -12383 26047 -12349 26048
rect -12348 26047 -12346 26067
rect -12276 26047 -12274 26067
rect -12252 26047 -12250 26067
rect -12156 26047 -12154 26067
rect -12060 26047 -12058 26067
rect -11844 26047 -11842 26067
rect -11796 26047 -11794 26067
rect -11676 26047 -11674 26067
rect -11580 26047 -11578 26067
rect -11556 26047 -11554 26067
rect -11508 26047 -11506 26067
rect -11460 26047 -11458 26067
rect -11436 26047 -11434 26067
rect -11364 26047 -11362 26067
rect -11340 26047 -11338 26067
rect -11292 26047 -11290 26067
rect -11196 26047 -11194 26067
rect -11124 26047 -11122 26067
rect -11100 26047 -11098 26067
rect -11028 26047 -11026 26067
rect -11004 26047 -11002 26067
rect -10788 26047 -10786 26067
rect -10740 26047 -10738 26067
rect -10668 26047 -10666 26067
rect -10644 26047 -10642 26067
rect -9996 26047 -9994 26067
rect -9708 26047 -9706 26067
rect -9612 26047 -9610 26067
rect -9516 26047 -9514 26067
rect -9468 26047 -9466 26067
rect -9420 26047 -9418 26067
rect -9396 26047 -9394 26067
rect -9372 26047 -9370 26067
rect -9300 26047 -9298 26067
rect -9252 26047 -9250 26067
rect -9084 26047 -9082 26067
rect -9057 26064 -9043 26067
rect -9036 26064 -9033 26067
rect -8988 26047 -8986 26067
rect -8940 26047 -8938 26067
rect -8892 26047 -8890 26067
rect -8772 26047 -8770 26067
rect -8604 26047 -8602 26067
rect -8484 26047 -8482 26067
rect -8457 26064 -8443 26067
rect -8436 26067 7781 26071
rect -8436 26064 -8419 26067
rect -8436 26047 -8434 26064
rect -8388 26047 -8386 26067
rect -8364 26047 -8362 26067
rect -8340 26047 -8338 26067
rect -8268 26047 -8266 26067
rect -8100 26047 -8098 26067
rect -8052 26047 -8050 26067
rect -7932 26047 -7930 26067
rect -7692 26047 -7690 26067
rect -7620 26047 -7618 26067
rect -7524 26047 -7522 26067
rect -7356 26047 -7354 26067
rect -7308 26047 -7306 26067
rect -7212 26047 -7210 26067
rect -7188 26047 -7186 26067
rect -7116 26047 -7114 26067
rect -7068 26047 -7066 26067
rect -6972 26047 -6970 26067
rect -6948 26047 -6946 26067
rect -6876 26047 -6874 26067
rect -6852 26047 -6850 26067
rect -6780 26047 -6778 26067
rect -6756 26047 -6754 26067
rect -6660 26047 -6658 26067
rect -6612 26047 -6610 26067
rect -6516 26047 -6514 26067
rect -6492 26047 -6490 26067
rect -6420 26047 -6418 26067
rect -6396 26047 -6394 26067
rect -6372 26047 -6370 26067
rect -6324 26047 -6322 26067
rect -6156 26047 -6154 26067
rect -6143 26047 -6085 26048
rect -6060 26047 -6058 26067
rect -5940 26047 -5938 26067
rect -5892 26047 -5890 26067
rect -5652 26047 -5650 26067
rect -5268 26047 -5266 26067
rect -5196 26047 -5194 26067
rect -5172 26047 -5170 26067
rect -5100 26047 -5098 26067
rect -5076 26047 -5074 26067
rect -4980 26047 -4978 26067
rect -4956 26047 -4954 26067
rect -4884 26047 -4882 26067
rect -4860 26047 -4858 26067
rect -4788 26047 -4786 26067
rect -4692 26048 -4690 26067
rect -4727 26047 -4669 26048
rect -4644 26047 -4642 26067
rect -4596 26047 -4594 26067
rect -4548 26047 -4546 26067
rect -4308 26047 -4306 26067
rect -4260 26047 -4258 26067
rect -4212 26047 -4210 26067
rect -4164 26047 -4162 26067
rect -4116 26047 -4114 26067
rect -4020 26047 -4018 26067
rect -3876 26047 -3874 26067
rect -3732 26047 -3730 26067
rect -3588 26047 -3586 26067
rect -3564 26047 -3562 26067
rect -3516 26047 -3514 26067
rect -3492 26047 -3490 26067
rect -3468 26047 -3466 26067
rect -3420 26047 -3418 26067
rect -3324 26047 -3322 26067
rect -3252 26047 -3250 26067
rect -3228 26047 -3226 26067
rect -3156 26047 -3154 26067
rect -3132 26047 -3130 26067
rect -3060 26047 -3058 26067
rect -3012 26047 -3010 26067
rect -2964 26047 -2962 26067
rect -2916 26047 -2914 26067
rect -2892 26047 -2890 26067
rect -2879 26062 -2876 26067
rect -2869 26048 -2866 26062
rect -2868 26047 -2866 26048
rect -2820 26047 -2818 26067
rect -2796 26047 -2794 26067
rect -2772 26047 -2769 26064
rect -2700 26047 -2698 26067
rect -2676 26047 -2674 26067
rect -2604 26047 -2602 26067
rect -2580 26047 -2578 26067
rect -2364 26047 -2362 26067
rect -2268 26047 -2266 26067
rect -2244 26047 -2242 26067
rect -2172 26047 -2170 26067
rect -2148 26047 -2146 26067
rect -2076 26047 -2074 26067
rect -2052 26047 -2050 26067
rect -1980 26047 -1978 26067
rect -1884 26047 -1882 26067
rect -1836 26047 -1834 26067
rect -1716 26047 -1714 26067
rect -1596 26047 -1594 26067
rect -1572 26047 -1570 26067
rect -1476 26047 -1474 26067
rect -1380 26047 -1378 26067
rect -1356 26047 -1354 26067
rect -1308 26047 -1306 26067
rect -1260 26047 -1258 26067
rect -1140 26047 -1138 26067
rect -852 26047 -850 26067
rect -804 26064 -802 26067
rect -804 26047 -801 26064
rect -756 26047 -754 26067
rect -708 26047 -706 26067
rect -612 26047 -610 26067
rect -588 26047 -586 26067
rect -540 26047 -538 26067
rect -492 26047 -490 26067
rect -444 26047 -442 26067
rect -396 26047 -394 26067
rect -300 26047 -298 26067
rect -276 26047 -274 26067
rect -228 26047 -226 26067
rect -12 26047 -10 26067
rect 156 26047 158 26067
rect 204 26047 206 26067
rect 228 26047 230 26067
rect 252 26047 254 26067
rect 348 26047 350 26067
rect 468 26047 470 26067
rect 492 26047 494 26067
rect 564 26047 566 26067
rect 588 26047 590 26067
rect 636 26047 638 26067
rect 660 26047 662 26067
rect 732 26047 734 26067
rect 756 26047 758 26067
rect 852 26047 854 26067
rect 1020 26047 1022 26067
rect 1057 26062 1060 26067
rect 1068 26062 1070 26067
rect 1067 26048 1070 26062
rect 1092 26047 1094 26067
rect 1116 26047 1118 26067
rect 1164 26064 1166 26067
rect 1164 26047 1167 26064
rect 1212 26047 1214 26067
rect 1308 26047 1310 26067
rect 1332 26047 1334 26067
rect 1380 26047 1382 26067
rect 1428 26047 1430 26067
rect 1476 26047 1478 26067
rect 1524 26047 1526 26067
rect 1548 26047 1550 26067
rect 1620 26047 1622 26067
rect 1644 26047 1646 26067
rect 1692 26047 1694 26067
rect 1716 26047 1718 26067
rect 1740 26047 1742 26067
rect 1788 26047 1790 26067
rect 1884 26047 1886 26067
rect 1980 26047 1982 26067
rect 2028 26047 2030 26067
rect 2076 26047 2078 26067
rect 2100 26047 2102 26067
rect 2124 26047 2126 26067
rect 2172 26047 2174 26067
rect 2196 26047 2198 26067
rect 2220 26047 2222 26067
rect 2268 26047 2270 26067
rect 2292 26047 2294 26067
rect 2316 26047 2318 26067
rect 2364 26047 2366 26067
rect 2412 26047 2414 26067
rect 2460 26047 2462 26067
rect 2508 26047 2510 26067
rect 2580 26047 2582 26067
rect 2604 26047 2606 26067
rect 2676 26047 2678 26067
rect 2700 26047 2702 26067
rect 2748 26047 2750 26067
rect 2772 26047 2774 26067
rect 2796 26047 2798 26067
rect 2844 26047 2846 26067
rect 2868 26047 2870 26067
rect 2892 26047 2894 26067
rect 2940 26047 2942 26067
rect 3012 26047 3014 26067
rect 3108 26047 3110 26067
rect 3156 26047 3158 26067
rect 3252 26047 3254 26067
rect 3348 26047 3350 26067
rect 3396 26047 3398 26067
rect 3468 26047 3470 26067
rect 3492 26047 3494 26067
rect 3564 26047 3566 26067
rect 3612 26047 3614 26067
rect 3636 26047 3638 26067
rect 3660 26047 3662 26067
rect 3708 26047 3710 26067
rect 3732 26047 3734 26067
rect 3804 26047 3806 26067
rect 3828 26047 3830 26067
rect 3924 26047 3926 26067
rect 4020 26047 4022 26067
rect 4044 26047 4046 26067
rect 4092 26047 4094 26067
rect 4116 26047 4118 26067
rect 4140 26047 4142 26067
rect 4188 26047 4190 26067
rect 4212 26047 4214 26067
rect 4236 26047 4238 26067
rect 4308 26047 4310 26067
rect 4332 26047 4334 26067
rect 4404 26047 4406 26067
rect 4500 26047 4502 26067
rect 4596 26047 4598 26067
rect 4860 26047 4862 26067
rect 4956 26047 4958 26067
rect 4980 26047 4982 26067
rect 5004 26047 5006 26067
rect 5076 26047 5078 26067
rect 5100 26047 5102 26067
rect 5124 26047 5126 26067
rect 5172 26047 5174 26067
rect 5220 26047 5222 26067
rect 5268 26047 5270 26067
rect 5388 26047 5390 26067
rect 5484 26047 5486 26067
rect 5508 26047 5510 26067
rect 5532 26047 5534 26067
rect 5628 26047 5630 26067
rect 5652 26047 5654 26067
rect 5748 26047 5750 26067
rect 5796 26047 5798 26067
rect 5844 26047 5846 26067
rect 5892 26047 5894 26067
rect 6132 26047 6134 26067
rect 6180 26047 6182 26067
rect 6228 26047 6230 26067
rect 6252 26047 6254 26067
rect 6276 26047 6278 26067
rect 6324 26047 6326 26067
rect 6372 26047 6374 26067
rect 6492 26047 6494 26067
rect 6588 26047 6590 26067
rect 6612 26047 6614 26067
rect 6660 26047 6662 26067
rect 6684 26047 6686 26067
rect 6708 26047 6710 26067
rect 6780 26047 6782 26067
rect 6804 26047 6806 26067
rect 6828 26047 6830 26067
rect 6900 26047 6902 26067
rect 6924 26047 6926 26067
rect 7020 26047 7022 26067
rect 7140 26047 7142 26067
rect 7236 26047 7238 26067
rect 7332 26047 7334 26067
rect 7380 26047 7382 26067
rect 7428 26047 7430 26067
rect 7452 26047 7454 26067
rect 7476 26047 7478 26067
rect 7524 26047 7526 26067
rect 7548 26047 7550 26067
rect 7572 26047 7574 26067
rect 7620 26047 7622 26067
rect 7644 26047 7646 26067
rect 7668 26047 7670 26067
rect 7740 26047 7742 26067
rect 7767 26064 7781 26067
rect 7788 26067 30707 26071
rect 7788 26064 7805 26067
rect 7788 26047 7790 26064
rect 7825 26062 7828 26067
rect 7836 26062 7838 26067
rect 7835 26048 7838 26062
rect 7884 26047 7886 26067
rect 7932 26064 7934 26067
rect 7932 26047 7935 26064
rect 7956 26047 7958 26067
rect 7980 26047 7982 26067
rect 8028 26047 8030 26067
rect 8196 26047 8198 26067
rect 8244 26047 8246 26067
rect 8268 26047 8270 26067
rect 8292 26047 8294 26067
rect 8340 26047 8342 26067
rect 8364 26047 8366 26067
rect 8388 26047 8390 26067
rect 8436 26047 8438 26067
rect 8460 26047 8462 26067
rect 8556 26047 8558 26067
rect 8604 26047 8606 26067
rect 8652 26047 8654 26067
rect 8700 26047 8702 26067
rect 8724 26047 8726 26067
rect 8748 26047 8750 26067
rect 8820 26047 8822 26067
rect 8844 26047 8846 26067
rect 8868 26047 8870 26067
rect 9516 26047 9518 26067
rect 9612 26047 9614 26067
rect 9660 26047 9662 26067
rect 9684 26047 9686 26067
rect 9708 26047 9710 26067
rect 9756 26047 9758 26067
rect 9780 26047 9782 26067
rect 9804 26047 9806 26067
rect 9852 26047 9854 26067
rect 9876 26047 9878 26067
rect 9900 26047 9902 26067
rect 9948 26047 9950 26067
rect 9972 26047 9974 26067
rect 9996 26047 9998 26067
rect 10068 26047 10070 26067
rect 10092 26047 10094 26067
rect 10116 26047 10118 26067
rect 10164 26047 10166 26067
rect 10188 26047 10190 26067
rect 10212 26047 10214 26067
rect 10284 26047 10286 26067
rect 10308 26047 10310 26067
rect 10332 26047 10334 26067
rect 10380 26047 10382 26067
rect 10404 26047 10406 26067
rect 10428 26047 10430 26067
rect 10476 26047 10478 26067
rect 10500 26047 10502 26067
rect 10524 26047 10526 26067
rect 10572 26047 10574 26067
rect 10596 26047 10598 26067
rect 10620 26047 10622 26067
rect 10668 26047 10670 26067
rect 10692 26047 10694 26067
rect 10716 26047 10718 26067
rect 10788 26047 10790 26067
rect 10836 26047 10838 26067
rect 10956 26047 10958 26067
rect 11052 26047 11054 26067
rect 11076 26047 11078 26067
rect 11124 26047 11126 26067
rect 11172 26047 11174 26067
rect 11220 26047 11222 26067
rect 11340 26047 11342 26067
rect 11436 26047 11438 26067
rect 11532 26047 11534 26067
rect 11580 26047 11582 26067
rect 11628 26047 11630 26067
rect 11676 26047 11678 26067
rect 11724 26047 11726 26067
rect 11772 26047 11774 26067
rect 11796 26047 11798 26067
rect 11892 26047 11894 26067
rect 11988 26047 11990 26067
rect 12060 26047 12062 26067
rect 12132 26047 12134 26067
rect 12228 26047 12230 26067
rect 12276 26047 12278 26067
rect 12324 26047 12326 26067
rect 12420 26047 12422 26067
rect 12444 26047 12446 26067
rect 12492 26047 12494 26067
rect 12516 26047 12518 26067
rect 12540 26047 12542 26067
rect 12588 26047 12590 26067
rect 12636 26047 12638 26067
rect 12732 26047 12734 26067
rect 12756 26047 12758 26067
rect 12804 26047 12806 26067
rect 12828 26047 12830 26067
rect 12852 26047 12854 26067
rect 12900 26047 12902 26067
rect 12948 26047 12950 26067
rect 13044 26047 13046 26067
rect 13068 26047 13070 26067
rect 13116 26047 13118 26067
rect 13284 26047 13286 26067
rect 13332 26047 13334 26067
rect 13428 26047 13430 26067
rect 13524 26047 13526 26067
rect 13572 26047 13574 26067
rect 13644 26047 13646 26067
rect 13668 26047 13670 26067
rect 13764 26047 13766 26067
rect 13812 26047 13814 26067
rect 13860 26047 13862 26067
rect 13908 26047 13910 26067
rect 13956 26047 13958 26067
rect 14004 26047 14006 26067
rect 14100 26047 14102 26067
rect 14196 26047 14198 26067
rect 14292 26047 14294 26067
rect 15132 26047 15134 26067
rect 15180 26047 15182 26067
rect 15228 26047 15230 26067
rect 15252 26047 15254 26067
rect 15324 26047 15326 26067
rect 15396 26047 15398 26067
rect 15420 26047 15422 26067
rect 15492 26047 15494 26067
rect 15540 26047 15542 26067
rect 15636 26047 15638 26067
rect 15660 26047 15662 26067
rect 15708 26047 15710 26067
rect 15732 26047 15734 26067
rect 15756 26047 15758 26067
rect 15804 26047 15806 26067
rect 15828 26047 15830 26067
rect 15852 26047 15854 26067
rect 15900 26047 15902 26067
rect 15948 26047 15950 26067
rect 15996 26047 15998 26067
rect 16044 26047 16046 26067
rect 16081 26062 16084 26067
rect 16092 26062 16094 26067
rect 16091 26048 16094 26062
rect 16164 26047 16167 26064
rect 16260 26047 16262 26067
rect 16308 26047 16310 26067
rect 16332 26047 16334 26067
rect 16356 26047 16358 26067
rect 16404 26047 16406 26067
rect 16452 26047 16454 26067
rect 16548 26047 16550 26067
rect 16572 26047 16574 26067
rect 16620 26047 16622 26067
rect 16668 26047 16670 26067
rect 16716 26047 16718 26067
rect 16764 26047 16766 26067
rect 16812 26047 16814 26067
rect 16884 26047 16886 26067
rect 16908 26047 16910 26067
rect 16980 26047 16982 26067
rect 17052 26047 17054 26067
rect 17196 26047 17198 26067
rect 17220 26047 17222 26067
rect 17292 26047 17294 26067
rect 17316 26047 17318 26067
rect 18084 26047 18086 26067
rect 18132 26047 18134 26067
rect 18396 26047 18398 26067
rect 18492 26047 18494 26067
rect 18516 26047 18518 26067
rect 18564 26047 18566 26067
rect 18612 26047 18614 26067
rect 18660 26047 18662 26067
rect 18708 26047 18710 26067
rect 18756 26047 18758 26067
rect 18804 26047 18806 26067
rect 18852 26047 18854 26067
rect 18900 26047 18902 26067
rect 18996 26047 18998 26067
rect 19020 26047 19022 26067
rect 19092 26047 19094 26067
rect 19116 26047 19118 26067
rect 19140 26047 19142 26067
rect 19188 26047 19190 26067
rect 19236 26047 19238 26067
rect 19332 26047 19334 26067
rect 19476 26047 19478 26067
rect 19609 26062 19612 26067
rect 19620 26062 19622 26067
rect 19619 26048 19622 26062
rect 19716 26064 19718 26067
rect 19716 26047 19719 26064
rect 19788 26047 19790 26067
rect 19836 26047 19838 26067
rect 19860 26047 19862 26067
rect 19884 26047 19886 26067
rect 19932 26047 19934 26067
rect 19956 26047 19958 26067
rect 19980 26047 19982 26067
rect 20028 26047 20030 26067
rect 20052 26047 20054 26067
rect 20076 26047 20078 26067
rect 20148 26047 20150 26067
rect 20172 26047 20174 26067
rect 20196 26047 20198 26067
rect 20268 26047 20270 26067
rect 20292 26047 20294 26067
rect 20388 26047 20390 26067
rect 20412 26047 20414 26067
rect 20508 26047 20510 26067
rect 20556 26047 20558 26067
rect 20604 26047 20606 26067
rect 20916 26047 20918 26067
rect 20964 26047 20966 26067
rect 21012 26047 21014 26067
rect 21060 26047 21062 26067
rect 21084 26047 21086 26067
rect 21108 26047 21110 26067
rect 21204 26047 21206 26067
rect 21300 26047 21302 26067
rect 21324 26047 21326 26067
rect 21444 26047 21446 26067
rect 21468 26047 21470 26067
rect 21564 26047 21566 26067
rect 21612 26047 21614 26067
rect 21684 26047 21686 26067
rect 21708 26047 21710 26067
rect 21828 26047 21830 26067
rect 21924 26047 21926 26067
rect 22068 26047 22070 26067
rect 22188 26047 22190 26067
rect 22212 26047 22214 26067
rect 22884 26047 22886 26067
rect 22980 26047 22982 26067
rect 23076 26047 23078 26067
rect 23100 26047 23102 26067
rect 23124 26047 23126 26067
rect 23244 26047 23246 26067
rect 23340 26047 23342 26067
rect 23412 26047 23414 26067
rect 23556 26047 23558 26067
rect 23628 26047 23630 26067
rect 23652 26047 23654 26067
rect 23676 26047 23678 26067
rect 23724 26047 23726 26067
rect 23772 26047 23774 26067
rect 23820 26047 23822 26067
rect 23868 26047 23870 26067
rect 23916 26047 23918 26067
rect 24012 26047 24014 26067
rect 24084 26047 24086 26067
rect 24303 26064 24317 26067
rect 24396 26047 24398 26067
rect 24492 26047 24494 26067
rect 24516 26047 24518 26067
rect 24588 26047 24590 26067
rect 24612 26047 24614 26067
rect 24708 26048 24710 26067
rect 24673 26047 24731 26048
rect 24732 26047 24734 26067
rect 24756 26047 24758 26067
rect 24852 26047 24854 26067
rect 24876 26047 24878 26067
rect 24972 26047 24974 26067
rect 24996 26047 24998 26067
rect 25068 26047 25070 26067
rect 25164 26047 25166 26067
rect 25260 26047 25262 26067
rect 25308 26047 25310 26067
rect 25356 26047 25358 26067
rect 25380 26047 25382 26067
rect 25404 26047 25406 26067
rect 25452 26047 25454 26067
rect 25500 26047 25502 26067
rect 25596 26047 25598 26067
rect 26929 26047 26987 26048
rect 27108 26047 27110 26067
rect 27324 26047 27326 26067
rect 27396 26047 27398 26067
rect 27420 26047 27422 26067
rect 27540 26047 27542 26067
rect 27564 26047 27566 26067
rect 30564 26047 30566 26067
rect 30660 26048 30662 26067
rect 30649 26047 30683 26048
rect -17433 26043 -17059 26047
rect -17433 26040 -17419 26043
rect -17388 26040 -17386 26043
rect -17217 26040 -17203 26043
rect -17073 26040 -17059 26043
rect -17052 26043 -14107 26047
rect -17052 26040 -17035 26043
rect -17388 26023 -17385 26040
rect -17052 26023 -17050 26040
rect -16836 26023 -16834 26043
rect -16764 26023 -16762 26043
rect -16740 26023 -16738 26043
rect -16415 26023 -16381 26024
rect -17409 26019 -16381 26023
rect -17409 26016 -17395 26019
rect -17388 26016 -17385 26019
rect -17385 25999 -17365 26000
rect -17052 25999 -17050 26019
rect -16836 25999 -16834 26019
rect -16809 26016 -16795 26019
rect -16764 25999 -16762 26019
rect -16740 25999 -16738 26019
rect -16415 26014 -16412 26019
rect -16405 26000 -16402 26014
rect -16404 25999 -16402 26000
rect -16380 25999 -16378 26043
rect -16356 25999 -16354 26043
rect -16343 26023 -16309 26024
rect -16284 26023 -16282 26043
rect -16260 26023 -16258 26043
rect -16236 26023 -16234 26043
rect -15324 26023 -15322 26043
rect -15084 26023 -15082 26043
rect -14868 26023 -14866 26043
rect -14772 26023 -14770 26043
rect -14735 26038 -14732 26043
rect -14724 26038 -14722 26043
rect -14725 26024 -14722 26038
rect -14508 26023 -14506 26043
rect -14436 26023 -14434 26043
rect -14340 26023 -14338 26043
rect -14244 26023 -14242 26043
rect -14121 26040 -14107 26043
rect -14097 26043 -2779 26047
rect -14097 26040 -14083 26043
rect -14076 26040 -14073 26043
rect -13980 26023 -13978 26043
rect -13932 26023 -13930 26043
rect -13884 26023 -13882 26043
rect -13788 26023 -13786 26043
rect -13572 26023 -13570 26043
rect -13500 26023 -13498 26043
rect -13356 26023 -13354 26043
rect -13284 26023 -13282 26043
rect -13068 26023 -13066 26043
rect -12828 26023 -12826 26043
rect -12780 26023 -12778 26043
rect -12660 26023 -12658 26043
rect -12564 26023 -12562 26043
rect -12492 26023 -12490 26043
rect -12396 26023 -12394 26043
rect -12348 26023 -12346 26043
rect -12276 26040 -12274 26043
rect -12276 26023 -12273 26040
rect -12252 26023 -12250 26043
rect -12156 26023 -12154 26043
rect -12060 26023 -12058 26043
rect -11844 26023 -11842 26043
rect -11796 26023 -11794 26043
rect -11676 26023 -11674 26043
rect -11580 26023 -11578 26043
rect -11556 26023 -11554 26043
rect -11508 26023 -11506 26043
rect -11460 26023 -11458 26043
rect -11436 26023 -11434 26043
rect -11423 26023 -11365 26024
rect -11364 26023 -11362 26043
rect -11340 26023 -11338 26043
rect -11292 26023 -11290 26043
rect -11196 26023 -11194 26043
rect -11124 26023 -11122 26043
rect -11100 26023 -11098 26043
rect -11028 26023 -11026 26043
rect -11004 26023 -11002 26043
rect -10788 26023 -10786 26043
rect -10740 26023 -10738 26043
rect -10668 26023 -10666 26043
rect -10644 26023 -10642 26043
rect -9996 26023 -9994 26043
rect -9708 26023 -9706 26043
rect -9612 26023 -9610 26043
rect -9516 26023 -9514 26043
rect -9468 26023 -9466 26043
rect -9420 26023 -9418 26043
rect -9396 26023 -9394 26043
rect -9372 26023 -9370 26043
rect -9300 26023 -9298 26043
rect -9252 26023 -9250 26043
rect -9084 26023 -9082 26043
rect -8988 26023 -8986 26043
rect -8940 26023 -8938 26043
rect -8892 26023 -8890 26043
rect -8772 26023 -8770 26043
rect -8604 26023 -8602 26043
rect -8484 26023 -8482 26043
rect -8436 26023 -8434 26043
rect -8388 26023 -8386 26043
rect -8364 26023 -8362 26043
rect -8340 26023 -8338 26043
rect -8268 26023 -8266 26043
rect -8100 26023 -8098 26043
rect -8052 26023 -8050 26043
rect -7932 26023 -7930 26043
rect -7692 26023 -7690 26043
rect -7620 26023 -7618 26043
rect -7524 26023 -7522 26043
rect -7356 26023 -7354 26043
rect -7308 26023 -7306 26043
rect -7212 26023 -7210 26043
rect -7188 26023 -7186 26043
rect -7116 26023 -7114 26043
rect -7068 26023 -7066 26043
rect -6972 26023 -6970 26043
rect -6948 26023 -6946 26043
rect -6876 26023 -6874 26043
rect -6852 26023 -6850 26043
rect -6780 26023 -6778 26043
rect -6756 26023 -6754 26043
rect -6660 26023 -6658 26043
rect -6612 26023 -6610 26043
rect -6516 26023 -6514 26043
rect -6492 26023 -6490 26043
rect -6420 26023 -6418 26043
rect -6396 26023 -6394 26043
rect -6372 26023 -6370 26043
rect -6324 26023 -6322 26043
rect -6156 26023 -6154 26043
rect -6060 26023 -6058 26043
rect -6036 26023 -6033 26040
rect -5940 26023 -5938 26043
rect -5892 26023 -5890 26043
rect -5652 26023 -5650 26043
rect -5268 26023 -5266 26043
rect -5196 26023 -5194 26043
rect -5172 26023 -5170 26043
rect -5100 26023 -5098 26043
rect -5076 26023 -5074 26043
rect -4980 26023 -4978 26043
rect -4956 26023 -4954 26043
rect -4884 26023 -4882 26043
rect -4860 26023 -4858 26043
rect -4788 26023 -4786 26043
rect -4703 26038 -4700 26043
rect -4692 26038 -4690 26043
rect -4693 26024 -4690 26038
rect -4644 26023 -4642 26043
rect -4596 26040 -4594 26043
rect -4596 26023 -4593 26040
rect -4548 26023 -4546 26043
rect -4308 26023 -4306 26043
rect -4260 26023 -4258 26043
rect -4212 26023 -4210 26043
rect -4164 26023 -4162 26043
rect -4116 26023 -4114 26043
rect -4020 26023 -4018 26043
rect -3876 26023 -3874 26043
rect -3732 26023 -3730 26043
rect -3588 26023 -3586 26043
rect -3564 26023 -3562 26043
rect -3516 26023 -3514 26043
rect -3492 26023 -3490 26043
rect -3468 26023 -3466 26043
rect -3420 26023 -3418 26043
rect -3324 26023 -3322 26043
rect -3252 26023 -3250 26043
rect -3228 26023 -3226 26043
rect -3156 26023 -3154 26043
rect -3132 26023 -3130 26043
rect -3060 26023 -3058 26043
rect -3012 26023 -3010 26043
rect -2964 26023 -2962 26043
rect -2916 26023 -2914 26043
rect -2892 26023 -2890 26043
rect -2868 26023 -2866 26043
rect -2820 26023 -2818 26043
rect -2796 26023 -2794 26043
rect -2793 26040 -2779 26043
rect -2772 26043 1133 26047
rect -2772 26040 -2755 26043
rect -2772 26023 -2770 26040
rect -2700 26023 -2698 26043
rect -2676 26023 -2674 26043
rect -2604 26023 -2602 26043
rect -2580 26023 -2578 26043
rect -2364 26023 -2362 26043
rect -2268 26023 -2266 26043
rect -2244 26023 -2242 26043
rect -2172 26023 -2170 26043
rect -2148 26023 -2146 26043
rect -2076 26023 -2074 26043
rect -2052 26023 -2050 26043
rect -1980 26023 -1978 26043
rect -1884 26023 -1882 26043
rect -1836 26023 -1834 26043
rect -1716 26023 -1714 26043
rect -1596 26023 -1594 26043
rect -1572 26023 -1570 26043
rect -1476 26023 -1474 26043
rect -1380 26023 -1378 26043
rect -1356 26023 -1354 26043
rect -1308 26023 -1306 26043
rect -1260 26023 -1258 26043
rect -1140 26023 -1138 26043
rect -852 26023 -850 26043
rect -825 26040 -811 26043
rect -804 26040 -801 26043
rect -756 26023 -754 26043
rect -708 26023 -706 26043
rect -612 26023 -610 26043
rect -588 26023 -586 26043
rect -540 26023 -538 26043
rect -492 26023 -490 26043
rect -444 26023 -442 26043
rect -396 26023 -394 26043
rect -300 26023 -298 26043
rect -276 26023 -274 26043
rect -228 26023 -226 26043
rect -12 26023 -10 26043
rect 156 26023 158 26043
rect 204 26023 206 26043
rect 228 26023 230 26043
rect 252 26023 254 26043
rect 348 26023 350 26043
rect 468 26023 470 26043
rect 492 26023 494 26043
rect 564 26023 566 26043
rect 588 26023 590 26043
rect 636 26023 638 26043
rect 660 26023 662 26043
rect 732 26023 734 26043
rect 756 26023 758 26043
rect 852 26023 854 26043
rect 1020 26023 1022 26043
rect 1092 26023 1094 26043
rect 1116 26023 1118 26043
rect 1119 26040 1133 26043
rect 1143 26043 7901 26047
rect 1143 26040 1157 26043
rect 1164 26040 1167 26043
rect 1212 26023 1214 26043
rect 1308 26023 1310 26043
rect 1332 26023 1334 26043
rect 1380 26023 1382 26043
rect 1428 26023 1430 26043
rect 1476 26023 1478 26043
rect 1524 26023 1526 26043
rect 1548 26023 1550 26043
rect 1620 26023 1622 26043
rect 1644 26023 1646 26043
rect 1692 26023 1694 26043
rect 1716 26023 1718 26043
rect 1740 26023 1742 26043
rect 1788 26023 1790 26043
rect 1884 26023 1886 26043
rect 1980 26023 1982 26043
rect 2028 26023 2030 26043
rect 2076 26023 2078 26043
rect 2100 26023 2102 26043
rect 2124 26023 2126 26043
rect 2172 26023 2174 26043
rect 2196 26023 2198 26043
rect 2220 26023 2222 26043
rect 2268 26023 2270 26043
rect 2292 26023 2294 26043
rect 2316 26023 2318 26043
rect 2364 26023 2366 26043
rect 2412 26023 2414 26043
rect 2460 26023 2462 26043
rect 2508 26023 2510 26043
rect 2580 26023 2582 26043
rect 2604 26023 2606 26043
rect 2676 26023 2678 26043
rect 2700 26023 2702 26043
rect 2748 26023 2750 26043
rect 2772 26023 2774 26043
rect 2796 26023 2798 26043
rect 2844 26023 2846 26043
rect 2868 26023 2870 26043
rect 2892 26023 2894 26043
rect 2940 26023 2942 26043
rect 3012 26023 3014 26043
rect 3108 26023 3110 26043
rect 3156 26023 3158 26043
rect 3252 26023 3254 26043
rect 3348 26023 3350 26043
rect 3396 26023 3398 26043
rect 3468 26023 3470 26043
rect 3492 26023 3494 26043
rect 3564 26023 3566 26043
rect 3612 26023 3614 26043
rect 3636 26023 3638 26043
rect 3660 26023 3662 26043
rect 3708 26023 3710 26043
rect 3732 26023 3734 26043
rect 3804 26023 3806 26043
rect 3828 26023 3830 26043
rect 3924 26023 3926 26043
rect 4020 26023 4022 26043
rect 4044 26023 4046 26043
rect 4092 26023 4094 26043
rect 4116 26023 4118 26043
rect 4140 26023 4142 26043
rect 4188 26023 4190 26043
rect 4212 26023 4214 26043
rect 4236 26023 4238 26043
rect 4308 26023 4310 26043
rect 4332 26023 4334 26043
rect 4404 26023 4406 26043
rect 4500 26023 4502 26043
rect 4596 26023 4598 26043
rect 4860 26023 4862 26043
rect 4956 26023 4958 26043
rect 4980 26023 4982 26043
rect 5004 26023 5006 26043
rect 5076 26023 5078 26043
rect 5100 26023 5102 26043
rect 5124 26023 5126 26043
rect 5172 26023 5174 26043
rect 5220 26023 5222 26043
rect 5268 26023 5270 26043
rect 5388 26023 5390 26043
rect 5484 26023 5486 26043
rect 5508 26023 5510 26043
rect 5532 26023 5534 26043
rect 5628 26023 5630 26043
rect 5652 26023 5654 26043
rect 5748 26023 5750 26043
rect 5796 26023 5798 26043
rect 5844 26023 5846 26043
rect 5892 26023 5894 26043
rect 6132 26023 6134 26043
rect 6180 26023 6182 26043
rect 6228 26023 6230 26043
rect 6252 26023 6254 26043
rect 6276 26023 6278 26043
rect 6324 26023 6326 26043
rect 6372 26023 6374 26043
rect 6492 26023 6494 26043
rect 6588 26023 6590 26043
rect 6612 26023 6614 26043
rect 6660 26023 6662 26043
rect 6684 26023 6686 26043
rect 6708 26023 6710 26043
rect 6780 26023 6782 26043
rect 6804 26023 6806 26043
rect 6828 26023 6830 26043
rect 6900 26023 6902 26043
rect 6924 26023 6926 26043
rect 7020 26023 7022 26043
rect 7140 26023 7142 26043
rect 7236 26023 7238 26043
rect 7332 26023 7334 26043
rect 7380 26023 7382 26043
rect 7428 26023 7430 26043
rect 7452 26023 7454 26043
rect 7476 26023 7478 26043
rect 7524 26023 7526 26043
rect 7548 26023 7550 26043
rect 7572 26023 7574 26043
rect 7620 26023 7622 26043
rect 7644 26023 7646 26043
rect 7668 26023 7670 26043
rect 7740 26023 7742 26043
rect 7788 26023 7790 26043
rect 7884 26023 7886 26043
rect 7887 26040 7901 26043
rect 7911 26043 16157 26047
rect 7911 26040 7925 26043
rect 7932 26040 7935 26043
rect 7956 26023 7958 26043
rect 7980 26023 7982 26043
rect 8028 26023 8030 26043
rect 8196 26023 8198 26043
rect 8244 26023 8246 26043
rect 8268 26023 8270 26043
rect 8292 26023 8294 26043
rect 8340 26023 8342 26043
rect 8364 26023 8366 26043
rect 8388 26023 8390 26043
rect 8436 26023 8438 26043
rect 8460 26023 8462 26043
rect 8556 26023 8558 26043
rect 8604 26023 8606 26043
rect 8652 26023 8654 26043
rect 8700 26023 8702 26043
rect 8724 26023 8726 26043
rect 8748 26023 8750 26043
rect 8820 26023 8822 26043
rect 8844 26023 8846 26043
rect 8868 26023 8870 26043
rect 9516 26023 9518 26043
rect 9612 26023 9614 26043
rect 9660 26023 9662 26043
rect 9684 26023 9686 26043
rect 9708 26023 9710 26043
rect 9756 26023 9758 26043
rect 9780 26023 9782 26043
rect 9804 26023 9806 26043
rect 9852 26023 9854 26043
rect 9876 26023 9878 26043
rect 9900 26023 9902 26043
rect 9948 26023 9950 26043
rect 9972 26023 9974 26043
rect 9996 26023 9998 26043
rect 10068 26023 10070 26043
rect 10092 26023 10094 26043
rect 10116 26023 10118 26043
rect 10164 26023 10166 26043
rect 10188 26023 10190 26043
rect 10212 26023 10214 26043
rect 10284 26023 10286 26043
rect 10308 26023 10310 26043
rect 10332 26023 10334 26043
rect 10380 26023 10382 26043
rect 10404 26023 10406 26043
rect 10428 26023 10430 26043
rect 10476 26023 10478 26043
rect 10500 26023 10502 26043
rect 10524 26023 10526 26043
rect 10572 26023 10574 26043
rect 10596 26023 10598 26043
rect 10620 26023 10622 26043
rect 10668 26023 10670 26043
rect 10692 26023 10694 26043
rect 10716 26023 10718 26043
rect 10788 26023 10790 26043
rect 10836 26023 10838 26043
rect 10956 26023 10958 26043
rect 11052 26023 11054 26043
rect 11076 26023 11078 26043
rect 11124 26023 11126 26043
rect 11172 26023 11174 26043
rect 11220 26023 11222 26043
rect 11340 26023 11342 26043
rect 11436 26023 11438 26043
rect 11532 26023 11534 26043
rect 11580 26023 11582 26043
rect 11628 26023 11630 26043
rect 11676 26023 11678 26043
rect 11724 26023 11726 26043
rect 11772 26023 11774 26043
rect 11796 26023 11798 26043
rect 11892 26023 11894 26043
rect 11988 26023 11990 26043
rect 12060 26023 12062 26043
rect 12132 26023 12134 26043
rect 12228 26023 12230 26043
rect 12276 26023 12278 26043
rect 12324 26023 12326 26043
rect 12420 26023 12422 26043
rect 12444 26023 12446 26043
rect 12492 26023 12494 26043
rect 12516 26023 12518 26043
rect 12540 26023 12542 26043
rect 12588 26023 12590 26043
rect 12636 26023 12638 26043
rect 12732 26023 12734 26043
rect 12756 26023 12758 26043
rect 12804 26023 12806 26043
rect 12828 26023 12830 26043
rect 12852 26023 12854 26043
rect 12900 26023 12902 26043
rect 12948 26023 12950 26043
rect 13044 26023 13046 26043
rect 13068 26023 13070 26043
rect 13116 26023 13118 26043
rect 13284 26023 13286 26043
rect 13332 26023 13334 26043
rect 13428 26023 13430 26043
rect 13524 26023 13526 26043
rect 13572 26023 13574 26043
rect 13644 26023 13646 26043
rect 13668 26023 13670 26043
rect 13764 26023 13766 26043
rect 13812 26023 13814 26043
rect 13860 26023 13862 26043
rect 13908 26023 13910 26043
rect 13956 26023 13958 26043
rect 14004 26023 14006 26043
rect 14100 26023 14102 26043
rect 14196 26023 14198 26043
rect 14292 26023 14294 26043
rect 15132 26023 15134 26043
rect 15180 26023 15182 26043
rect 15228 26023 15230 26043
rect 15252 26023 15254 26043
rect 15324 26023 15326 26043
rect 15396 26023 15398 26043
rect 15420 26023 15422 26043
rect 15492 26023 15494 26043
rect 15540 26023 15542 26043
rect 15636 26023 15638 26043
rect 15660 26023 15662 26043
rect 15708 26023 15710 26043
rect 15732 26023 15734 26043
rect 15756 26023 15758 26043
rect 15804 26023 15806 26043
rect 15828 26023 15830 26043
rect 15852 26023 15854 26043
rect 15900 26023 15902 26043
rect 15948 26023 15950 26043
rect 15996 26023 15998 26043
rect 16044 26023 16046 26043
rect 16143 26040 16157 26043
rect 16164 26043 30683 26047
rect 16164 26040 16181 26043
rect 16164 26023 16166 26040
rect 16260 26023 16262 26043
rect 16308 26023 16310 26043
rect 16332 26023 16334 26043
rect 16356 26023 16358 26043
rect 16404 26023 16406 26043
rect 16452 26023 16454 26043
rect 16548 26023 16550 26043
rect 16572 26023 16574 26043
rect 16620 26023 16622 26043
rect 16668 26023 16670 26043
rect 16716 26023 16718 26043
rect 16764 26023 16766 26043
rect 16812 26023 16814 26043
rect 16884 26023 16886 26043
rect 16908 26023 16910 26043
rect 16980 26023 16982 26043
rect 17052 26023 17054 26043
rect 17196 26023 17198 26043
rect 17220 26023 17222 26043
rect 17292 26023 17294 26043
rect 17316 26023 17318 26043
rect 18084 26023 18086 26043
rect 18132 26023 18134 26043
rect 18396 26023 18398 26043
rect 18492 26023 18494 26043
rect 18516 26023 18518 26043
rect 18564 26023 18566 26043
rect 18612 26023 18614 26043
rect 18660 26023 18662 26043
rect 18708 26023 18710 26043
rect 18756 26023 18758 26043
rect 18804 26023 18806 26043
rect 18852 26023 18854 26043
rect 18900 26023 18902 26043
rect 18996 26023 18998 26043
rect 19020 26023 19022 26043
rect 19092 26023 19094 26043
rect 19116 26023 19118 26043
rect 19140 26023 19142 26043
rect 19188 26023 19190 26043
rect 19236 26023 19238 26043
rect 19332 26023 19334 26043
rect 19476 26023 19478 26043
rect 19695 26040 19709 26043
rect 19716 26040 19719 26043
rect 19788 26023 19790 26043
rect 19836 26023 19838 26043
rect 19860 26023 19862 26043
rect 19884 26023 19886 26043
rect 19932 26023 19934 26043
rect 19956 26023 19958 26043
rect 19980 26023 19982 26043
rect 20028 26023 20030 26043
rect 20052 26023 20054 26043
rect 20076 26023 20078 26043
rect 20148 26023 20150 26043
rect 20172 26023 20174 26043
rect 20196 26023 20198 26043
rect 20268 26023 20270 26043
rect 20292 26023 20294 26043
rect 20388 26023 20390 26043
rect 20412 26023 20414 26043
rect 20508 26023 20510 26043
rect 20556 26023 20558 26043
rect 20604 26023 20606 26043
rect 20916 26023 20918 26043
rect 20964 26023 20966 26043
rect 21012 26023 21014 26043
rect 21060 26023 21062 26043
rect 21084 26023 21086 26043
rect 21108 26023 21110 26043
rect 21204 26023 21206 26043
rect 21300 26023 21302 26043
rect 21324 26023 21326 26043
rect 21444 26023 21446 26043
rect 21468 26023 21470 26043
rect 21564 26023 21566 26043
rect 21612 26023 21614 26043
rect 21684 26023 21686 26043
rect 21708 26023 21710 26043
rect 21828 26023 21830 26043
rect 21924 26023 21926 26043
rect 22068 26023 22070 26043
rect 22188 26023 22190 26043
rect 22212 26023 22214 26043
rect 22884 26023 22886 26043
rect 22980 26023 22982 26043
rect 23076 26023 23078 26043
rect 23100 26023 23102 26043
rect 23124 26023 23126 26043
rect 23244 26023 23246 26043
rect 23340 26023 23342 26043
rect 23412 26023 23414 26043
rect 23556 26023 23558 26043
rect 23628 26023 23630 26043
rect 23652 26023 23654 26043
rect 23676 26023 23678 26043
rect 23724 26023 23726 26043
rect 23772 26023 23774 26043
rect 23820 26023 23822 26043
rect 23868 26023 23870 26043
rect 23916 26023 23918 26043
rect 24012 26023 24014 26043
rect 24084 26023 24086 26043
rect 24396 26023 24398 26043
rect 24492 26023 24494 26043
rect 24516 26023 24518 26043
rect 24588 26023 24590 26043
rect 24612 26023 24614 26043
rect 24673 26038 24676 26043
rect 24697 26038 24700 26043
rect 24708 26038 24710 26043
rect 24683 26024 24686 26038
rect 24707 26024 24710 26038
rect 24684 26023 24686 26024
rect 24732 26023 24734 26043
rect 24756 26023 24758 26043
rect 24780 26023 24783 26040
rect 24852 26023 24854 26043
rect 24876 26023 24878 26043
rect 24972 26023 24974 26043
rect 24996 26023 24998 26043
rect 25068 26023 25070 26043
rect 25164 26023 25166 26043
rect 25260 26023 25262 26043
rect 25308 26023 25310 26043
rect 25356 26023 25358 26043
rect 25380 26023 25382 26043
rect 25404 26023 25406 26043
rect 25452 26023 25454 26043
rect 25500 26023 25502 26043
rect 25596 26023 25598 26043
rect 27036 26023 27039 26040
rect 27108 26023 27110 26043
rect 27324 26023 27326 26043
rect 27396 26023 27398 26043
rect 27420 26023 27422 26043
rect 27540 26023 27542 26043
rect 27564 26023 27566 26043
rect 30564 26024 30566 26043
rect 30649 26038 30652 26043
rect 30660 26038 30662 26043
rect 30659 26024 30662 26038
rect 30553 26023 30587 26024
rect -16343 26019 -6043 26023
rect -16319 26006 -16315 26014
rect -16329 26000 -16319 26006
rect -17385 25995 -16315 25999
rect -17385 25992 -17371 25995
rect -17279 25975 -17245 25976
rect -17052 25975 -17050 25995
rect -16871 25975 -16837 25976
rect -16836 25975 -16834 25995
rect -16764 25975 -16762 25995
rect -16740 25975 -16738 25995
rect -16404 25975 -16402 25995
rect -16380 25975 -16378 25995
rect -16356 25975 -16354 25995
rect -16329 25992 -16315 25995
rect -16284 25975 -16282 26019
rect -16260 25975 -16258 26019
rect -16236 26016 -16234 26019
rect -16236 25999 -16233 26016
rect -15407 25999 -15373 26000
rect -15324 25999 -15322 26019
rect -15084 25999 -15082 26019
rect -14868 25999 -14866 26019
rect -14772 25999 -14770 26019
rect -14649 26016 -14635 26019
rect -14508 25999 -14506 26019
rect -14436 25999 -14434 26019
rect -14340 25999 -14338 26019
rect -14244 26000 -14242 26019
rect -14255 25999 -14221 26000
rect -13980 25999 -13978 26019
rect -13932 25999 -13930 26019
rect -13884 25999 -13882 26019
rect -13788 25999 -13786 26019
rect -13572 25999 -13570 26019
rect -13500 25999 -13498 26019
rect -13356 25999 -13354 26019
rect -13284 25999 -13282 26019
rect -13068 25999 -13066 26019
rect -12828 25999 -12826 26019
rect -12780 25999 -12778 26019
rect -12660 25999 -12658 26019
rect -12564 25999 -12562 26019
rect -12492 25999 -12490 26019
rect -12396 25999 -12394 26019
rect -12348 25999 -12346 26019
rect -12297 26016 -12283 26019
rect -12276 26016 -12273 26019
rect -12252 25999 -12250 26019
rect -12156 25999 -12154 26019
rect -12060 25999 -12058 26019
rect -11844 25999 -11842 26019
rect -11796 25999 -11794 26019
rect -11676 25999 -11674 26019
rect -11580 25999 -11578 26019
rect -11556 25999 -11554 26019
rect -11508 25999 -11506 26019
rect -11460 25999 -11458 26019
rect -11436 25999 -11434 26019
rect -11423 26014 -11420 26019
rect -11413 26000 -11410 26014
rect -11412 25999 -11410 26000
rect -11364 25999 -11362 26019
rect -11340 25999 -11338 26019
rect -11292 26016 -11290 26019
rect -11292 25999 -11289 26016
rect -11196 25999 -11194 26019
rect -11124 25999 -11122 26019
rect -11100 25999 -11098 26019
rect -11028 25999 -11026 26019
rect -11004 26000 -11002 26019
rect -10788 26000 -10786 26019
rect -11015 25999 -10981 26000
rect -10799 25999 -10765 26000
rect -10740 25999 -10738 26019
rect -10668 25999 -10666 26019
rect -10644 25999 -10642 26019
rect -9996 25999 -9994 26019
rect -9708 25999 -9706 26019
rect -9612 25999 -9610 26019
rect -9516 25999 -9514 26019
rect -9468 25999 -9466 26019
rect -9420 25999 -9418 26019
rect -9396 25999 -9394 26019
rect -9372 26000 -9370 26019
rect -9383 25999 -9349 26000
rect -9300 25999 -9298 26019
rect -9252 25999 -9250 26019
rect -9084 25999 -9082 26019
rect -8988 25999 -8986 26019
rect -8940 26000 -8938 26019
rect -8951 25999 -8917 26000
rect -8892 25999 -8890 26019
rect -8772 25999 -8770 26019
rect -8604 25999 -8602 26019
rect -8484 25999 -8482 26019
rect -8436 25999 -8434 26019
rect -8388 25999 -8386 26019
rect -8364 25999 -8362 26019
rect -8340 25999 -8338 26019
rect -8268 25999 -8266 26019
rect -8100 25999 -8098 26019
rect -8052 25999 -8050 26019
rect -7932 25999 -7930 26019
rect -7692 25999 -7690 26019
rect -7620 25999 -7618 26019
rect -7524 25999 -7522 26019
rect -7356 25999 -7354 26019
rect -7308 25999 -7306 26019
rect -7212 25999 -7210 26019
rect -7188 25999 -7186 26019
rect -7116 25999 -7114 26019
rect -7068 25999 -7066 26019
rect -6972 25999 -6970 26019
rect -6948 25999 -6946 26019
rect -6876 25999 -6874 26019
rect -6852 25999 -6850 26019
rect -6780 25999 -6778 26019
rect -6756 25999 -6754 26019
rect -6660 25999 -6658 26019
rect -6612 25999 -6610 26019
rect -6516 25999 -6514 26019
rect -6492 25999 -6490 26019
rect -6420 25999 -6418 26019
rect -6396 25999 -6394 26019
rect -6372 25999 -6370 26019
rect -6324 25999 -6322 26019
rect -6156 25999 -6154 26019
rect -6060 25999 -6058 26019
rect -6057 26016 -6043 26019
rect -6036 26019 -4627 26023
rect -6036 26016 -6019 26019
rect -6036 25999 -6034 26016
rect -5940 25999 -5938 26019
rect -5892 25999 -5890 26019
rect -5652 25999 -5650 26019
rect -5268 25999 -5266 26019
rect -5196 25999 -5194 26019
rect -5172 25999 -5170 26019
rect -5100 25999 -5098 26019
rect -5076 25999 -5074 26019
rect -4980 25999 -4978 26019
rect -4956 25999 -4954 26019
rect -4884 25999 -4882 26019
rect -4860 25999 -4858 26019
rect -4788 25999 -4786 26019
rect -4644 25999 -4642 26019
rect -4641 26016 -4627 26019
rect -4617 26019 24773 26023
rect -4617 26016 -4603 26019
rect -4596 26016 -4593 26019
rect -4548 25999 -4546 26019
rect -4308 25999 -4306 26019
rect -4260 25999 -4258 26019
rect -4212 26000 -4210 26019
rect -4223 25999 -4189 26000
rect -4164 25999 -4162 26019
rect -4116 25999 -4114 26019
rect -4020 25999 -4018 26019
rect -3876 25999 -3874 26019
rect -3732 25999 -3730 26019
rect -3588 25999 -3586 26019
rect -3564 25999 -3562 26019
rect -3516 25999 -3514 26019
rect -3492 25999 -3490 26019
rect -3468 25999 -3466 26019
rect -3420 25999 -3418 26019
rect -3324 25999 -3322 26019
rect -3252 25999 -3250 26019
rect -3228 25999 -3226 26019
rect -3156 25999 -3154 26019
rect -3132 25999 -3130 26019
rect -3060 25999 -3058 26019
rect -3012 25999 -3010 26019
rect -2964 25999 -2962 26019
rect -2916 25999 -2914 26019
rect -2892 25999 -2890 26019
rect -2868 25999 -2866 26019
rect -2820 25999 -2818 26019
rect -2796 25999 -2794 26019
rect -2772 25999 -2770 26019
rect -2700 25999 -2698 26019
rect -2676 25999 -2674 26019
rect -2604 25999 -2602 26019
rect -2580 25999 -2578 26019
rect -2364 25999 -2362 26019
rect -2268 25999 -2266 26019
rect -2244 25999 -2242 26019
rect -2172 25999 -2170 26019
rect -2148 25999 -2146 26019
rect -2076 25999 -2074 26019
rect -2052 25999 -2050 26019
rect -1980 25999 -1978 26019
rect -1884 25999 -1882 26019
rect -1836 25999 -1834 26019
rect -1716 26000 -1714 26019
rect -1727 25999 -1693 26000
rect -1596 25999 -1594 26019
rect -1572 25999 -1570 26019
rect -1476 25999 -1474 26019
rect -1380 25999 -1378 26019
rect -1356 25999 -1354 26019
rect -1308 25999 -1306 26019
rect -1260 25999 -1258 26019
rect -1140 25999 -1138 26019
rect -852 25999 -850 26019
rect -756 25999 -754 26019
rect -708 25999 -706 26019
rect -612 25999 -610 26019
rect -588 25999 -586 26019
rect -540 25999 -538 26019
rect -492 25999 -490 26019
rect -444 25999 -442 26019
rect -396 25999 -394 26019
rect -300 25999 -298 26019
rect -276 25999 -274 26019
rect -228 25999 -226 26019
rect -71 25999 -37 26000
rect -12 25999 -10 26019
rect 156 25999 158 26019
rect 204 25999 206 26019
rect 228 25999 230 26019
rect 252 25999 254 26019
rect 348 25999 350 26019
rect 468 25999 470 26019
rect 492 25999 494 26019
rect 564 25999 566 26019
rect 588 25999 590 26019
rect 636 25999 638 26019
rect 660 25999 662 26019
rect 732 25999 734 26019
rect 756 25999 758 26019
rect 852 25999 854 26019
rect 1020 25999 1022 26019
rect 1092 25999 1094 26019
rect 1116 25999 1118 26019
rect 1212 25999 1214 26019
rect 1308 25999 1310 26019
rect 1332 25999 1334 26019
rect 1380 25999 1382 26019
rect 1428 25999 1430 26019
rect 1476 25999 1478 26019
rect 1524 25999 1526 26019
rect 1548 25999 1550 26019
rect 1620 25999 1622 26019
rect 1644 25999 1646 26019
rect 1692 25999 1694 26019
rect 1716 25999 1718 26019
rect 1740 25999 1742 26019
rect 1788 25999 1790 26019
rect 1884 25999 1886 26019
rect 1980 25999 1982 26019
rect 2028 25999 2030 26019
rect 2076 25999 2078 26019
rect 2100 25999 2102 26019
rect 2124 25999 2126 26019
rect 2172 25999 2174 26019
rect 2196 25999 2198 26019
rect 2220 25999 2222 26019
rect 2268 25999 2270 26019
rect 2292 25999 2294 26019
rect 2316 25999 2318 26019
rect 2364 25999 2366 26019
rect 2412 25999 2414 26019
rect 2460 25999 2462 26019
rect 2508 25999 2510 26019
rect 2580 25999 2582 26019
rect 2604 25999 2606 26019
rect 2676 25999 2678 26019
rect 2700 25999 2702 26019
rect 2748 25999 2750 26019
rect 2772 25999 2774 26019
rect 2796 25999 2798 26019
rect 2844 25999 2846 26019
rect 2868 25999 2870 26019
rect 2892 25999 2894 26019
rect 2940 25999 2942 26019
rect 3012 25999 3014 26019
rect 3108 25999 3110 26019
rect 3156 25999 3158 26019
rect 3252 25999 3254 26019
rect 3348 25999 3350 26019
rect 3396 25999 3398 26019
rect 3468 25999 3470 26019
rect 3492 25999 3494 26019
rect 3564 25999 3566 26019
rect 3612 25999 3614 26019
rect 3636 25999 3638 26019
rect 3660 25999 3662 26019
rect 3708 25999 3710 26019
rect 3732 25999 3734 26019
rect 3804 25999 3806 26019
rect 3828 25999 3830 26019
rect 3924 25999 3926 26019
rect 4020 25999 4022 26019
rect 4044 25999 4046 26019
rect 4092 25999 4094 26019
rect 4116 25999 4118 26019
rect 4140 25999 4142 26019
rect 4188 25999 4190 26019
rect 4212 25999 4214 26019
rect 4236 25999 4238 26019
rect 4308 25999 4310 26019
rect 4332 25999 4334 26019
rect 4404 25999 4406 26019
rect 4500 25999 4502 26019
rect 4596 25999 4598 26019
rect 4860 25999 4862 26019
rect 4956 25999 4958 26019
rect 4980 25999 4982 26019
rect 5004 25999 5006 26019
rect 5076 25999 5078 26019
rect 5100 25999 5102 26019
rect 5124 25999 5126 26019
rect 5172 25999 5174 26019
rect 5220 25999 5222 26019
rect 5268 25999 5270 26019
rect 5388 25999 5390 26019
rect 5484 25999 5486 26019
rect 5508 25999 5510 26019
rect 5532 25999 5534 26019
rect 5628 25999 5630 26019
rect 5652 25999 5654 26019
rect 5748 25999 5750 26019
rect 5796 25999 5798 26019
rect 5844 25999 5846 26019
rect 5892 25999 5894 26019
rect 6132 25999 6134 26019
rect 6180 25999 6182 26019
rect 6228 25999 6230 26019
rect 6252 25999 6254 26019
rect 6276 25999 6278 26019
rect 6324 25999 6326 26019
rect 6372 25999 6374 26019
rect 6492 25999 6494 26019
rect 6588 25999 6590 26019
rect 6612 25999 6614 26019
rect 6660 25999 6662 26019
rect 6684 25999 6686 26019
rect 6708 25999 6710 26019
rect 6780 25999 6782 26019
rect 6804 25999 6806 26019
rect 6828 25999 6830 26019
rect 6900 25999 6902 26019
rect 6924 25999 6926 26019
rect 7020 25999 7022 26019
rect 7140 25999 7142 26019
rect 7236 25999 7238 26019
rect 7332 25999 7334 26019
rect 7380 25999 7382 26019
rect 7428 25999 7430 26019
rect 7452 25999 7454 26019
rect 7476 25999 7478 26019
rect 7524 25999 7526 26019
rect 7548 25999 7550 26019
rect 7572 25999 7574 26019
rect 7620 25999 7622 26019
rect 7644 25999 7646 26019
rect 7668 25999 7670 26019
rect 7740 25999 7742 26019
rect 7788 25999 7790 26019
rect 7884 25999 7886 26019
rect 7956 25999 7958 26019
rect 7980 25999 7982 26019
rect 8028 25999 8030 26019
rect 8196 25999 8198 26019
rect 8244 25999 8246 26019
rect 8268 25999 8270 26019
rect 8292 25999 8294 26019
rect 8340 25999 8342 26019
rect 8364 25999 8366 26019
rect 8388 25999 8390 26019
rect 8436 25999 8438 26019
rect 8460 25999 8462 26019
rect 8556 25999 8558 26019
rect 8604 25999 8606 26019
rect 8652 25999 8654 26019
rect 8700 25999 8702 26019
rect 8724 25999 8726 26019
rect 8748 25999 8750 26019
rect 8820 25999 8822 26019
rect 8844 25999 8846 26019
rect 8868 25999 8870 26019
rect 9516 25999 9518 26019
rect 9612 25999 9614 26019
rect 9660 25999 9662 26019
rect 9684 25999 9686 26019
rect 9708 25999 9710 26019
rect 9756 25999 9758 26019
rect 9780 25999 9782 26019
rect 9804 25999 9806 26019
rect 9852 25999 9854 26019
rect 9876 25999 9878 26019
rect 9900 25999 9902 26019
rect 9948 25999 9950 26019
rect 9972 25999 9974 26019
rect 9996 25999 9998 26019
rect 10068 25999 10070 26019
rect 10092 25999 10094 26019
rect 10116 25999 10118 26019
rect 10164 25999 10166 26019
rect 10188 25999 10190 26019
rect 10212 25999 10214 26019
rect 10284 25999 10286 26019
rect 10308 25999 10310 26019
rect 10332 25999 10334 26019
rect 10380 25999 10382 26019
rect 10404 25999 10406 26019
rect 10428 25999 10430 26019
rect 10476 25999 10478 26019
rect 10500 25999 10502 26019
rect 10524 25999 10526 26019
rect 10572 25999 10574 26019
rect 10596 25999 10598 26019
rect 10620 25999 10622 26019
rect 10668 25999 10670 26019
rect 10692 25999 10694 26019
rect 10716 25999 10718 26019
rect 10788 25999 10790 26019
rect 10836 25999 10838 26019
rect 10956 25999 10958 26019
rect 11052 25999 11054 26019
rect 11076 25999 11078 26019
rect 11124 25999 11126 26019
rect 11172 25999 11174 26019
rect 11220 25999 11222 26019
rect 11340 25999 11342 26019
rect 11436 25999 11438 26019
rect 11532 25999 11534 26019
rect 11580 25999 11582 26019
rect 11628 25999 11630 26019
rect 11676 25999 11678 26019
rect 11724 25999 11726 26019
rect 11772 25999 11774 26019
rect 11796 25999 11798 26019
rect 11892 25999 11894 26019
rect 11988 25999 11990 26019
rect 12060 25999 12062 26019
rect 12132 25999 12134 26019
rect 12228 25999 12230 26019
rect 12276 25999 12278 26019
rect 12324 25999 12326 26019
rect 12420 25999 12422 26019
rect 12444 25999 12446 26019
rect 12492 25999 12494 26019
rect 12516 25999 12518 26019
rect 12540 25999 12542 26019
rect 12588 25999 12590 26019
rect 12636 25999 12638 26019
rect 12732 25999 12734 26019
rect 12756 25999 12758 26019
rect 12804 25999 12806 26019
rect 12828 25999 12830 26019
rect 12852 25999 12854 26019
rect 12900 25999 12902 26019
rect 12948 25999 12950 26019
rect 13044 25999 13046 26019
rect 13068 25999 13070 26019
rect 13116 25999 13118 26019
rect 13284 25999 13286 26019
rect 13332 25999 13334 26019
rect 13428 25999 13430 26019
rect 13524 25999 13526 26019
rect 13572 25999 13574 26019
rect 13644 25999 13646 26019
rect 13668 25999 13670 26019
rect 13764 25999 13766 26019
rect 13812 25999 13814 26019
rect 13860 25999 13862 26019
rect 13908 25999 13910 26019
rect 13956 25999 13958 26019
rect 14004 25999 14006 26019
rect 14100 25999 14102 26019
rect 14196 25999 14198 26019
rect 14257 25999 14291 26000
rect 14292 25999 14294 26019
rect 15132 25999 15134 26019
rect 15180 25999 15182 26019
rect 15228 25999 15230 26019
rect 15252 25999 15254 26019
rect 15324 25999 15326 26019
rect 15396 25999 15398 26019
rect 15420 25999 15422 26019
rect 15492 25999 15494 26019
rect 15540 25999 15542 26019
rect 15636 25999 15638 26019
rect 15660 25999 15662 26019
rect 15708 25999 15710 26019
rect 15732 25999 15734 26019
rect 15756 25999 15758 26019
rect 15804 25999 15806 26019
rect 15828 25999 15830 26019
rect 15852 25999 15854 26019
rect 15900 25999 15902 26019
rect 15948 25999 15950 26019
rect 15996 25999 15998 26019
rect 16044 25999 16046 26019
rect 16164 25999 16166 26019
rect 16260 25999 16262 26019
rect 16308 25999 16310 26019
rect 16332 25999 16334 26019
rect 16356 25999 16358 26019
rect 16404 25999 16406 26019
rect 16452 25999 16454 26019
rect 16548 25999 16550 26019
rect 16572 25999 16574 26019
rect 16620 25999 16622 26019
rect 16668 25999 16670 26019
rect 16716 25999 16718 26019
rect 16764 25999 16766 26019
rect 16812 25999 16814 26019
rect 16884 25999 16886 26019
rect 16908 25999 16910 26019
rect 16980 25999 16982 26019
rect 17052 25999 17054 26019
rect 17196 25999 17198 26019
rect 17220 25999 17222 26019
rect 17292 25999 17294 26019
rect 17316 25999 17318 26019
rect 18084 25999 18086 26019
rect 18132 25999 18134 26019
rect 18396 25999 18398 26019
rect 18492 25999 18494 26019
rect 18516 25999 18518 26019
rect 18564 25999 18566 26019
rect 18612 25999 18614 26019
rect 18660 25999 18662 26019
rect 18708 25999 18710 26019
rect 18756 25999 18758 26019
rect 18804 25999 18806 26019
rect 18852 25999 18854 26019
rect 18900 25999 18902 26019
rect 18996 25999 18998 26019
rect 19020 25999 19022 26019
rect 19092 25999 19094 26019
rect 19116 25999 19118 26019
rect 19140 25999 19142 26019
rect 19188 25999 19190 26019
rect 19236 25999 19238 26019
rect 19332 25999 19334 26019
rect 19476 25999 19478 26019
rect 19788 25999 19790 26019
rect 19836 25999 19838 26019
rect 19860 25999 19862 26019
rect 19884 25999 19886 26019
rect 19932 25999 19934 26019
rect 19956 25999 19958 26019
rect 19980 25999 19982 26019
rect 20028 25999 20030 26019
rect 20052 25999 20054 26019
rect 20076 25999 20078 26019
rect 20148 25999 20150 26019
rect 20172 25999 20174 26019
rect 20196 25999 20198 26019
rect 20268 25999 20270 26019
rect 20292 25999 20294 26019
rect 20388 25999 20390 26019
rect 20412 25999 20414 26019
rect 20508 25999 20510 26019
rect 20556 25999 20558 26019
rect 20604 25999 20606 26019
rect 20916 25999 20918 26019
rect 20964 25999 20966 26019
rect 21012 25999 21014 26019
rect 21060 25999 21062 26019
rect 21084 25999 21086 26019
rect 21108 25999 21110 26019
rect 21204 25999 21206 26019
rect 21300 25999 21302 26019
rect 21324 25999 21326 26019
rect 21444 25999 21446 26019
rect 21468 25999 21470 26019
rect 21564 25999 21566 26019
rect 21612 25999 21614 26019
rect 21684 25999 21686 26019
rect 21708 25999 21710 26019
rect 21828 25999 21830 26019
rect 21924 25999 21926 26019
rect 22068 25999 22070 26019
rect 22188 25999 22190 26019
rect 22212 25999 22214 26019
rect 22417 25999 22451 26000
rect 22884 25999 22886 26019
rect 22980 25999 22982 26019
rect 23076 25999 23078 26019
rect 23100 25999 23102 26019
rect 23124 25999 23126 26019
rect 23244 25999 23246 26019
rect 23340 25999 23342 26019
rect 23412 25999 23414 26019
rect 23497 25999 23555 26000
rect 23556 25999 23558 26019
rect 23628 25999 23630 26019
rect 23652 25999 23654 26019
rect 23676 25999 23678 26019
rect 23724 25999 23726 26019
rect 23772 25999 23774 26019
rect 23820 25999 23822 26019
rect 23868 25999 23870 26019
rect 23916 25999 23918 26019
rect 24012 25999 24014 26019
rect 24084 25999 24086 26019
rect 24396 25999 24398 26019
rect 24492 25999 24494 26019
rect 24516 25999 24518 26019
rect 24588 25999 24590 26019
rect 24612 25999 24614 26019
rect 24684 25999 24686 26019
rect 24732 25999 24734 26019
rect 24756 25999 24758 26019
rect 24759 26016 24773 26019
rect 24780 26019 27029 26023
rect 24780 26016 24797 26019
rect 24780 25999 24782 26016
rect 24852 25999 24854 26019
rect 24876 25999 24878 26019
rect 24972 25999 24974 26019
rect 24996 25999 24998 26019
rect 25068 25999 25070 26019
rect 25164 25999 25166 26019
rect 25260 25999 25262 26019
rect 25308 25999 25310 26019
rect 25356 25999 25358 26019
rect 25380 25999 25382 26019
rect 25404 25999 25406 26019
rect 25452 26000 25454 26019
rect 25417 25999 25475 26000
rect 25500 25999 25502 26019
rect 25596 25999 25598 26019
rect 27015 26016 27029 26019
rect 27036 26019 30587 26023
rect 27036 26016 27053 26019
rect 27036 25999 27038 26016
rect 27108 25999 27110 26019
rect 27324 25999 27326 26019
rect 27396 25999 27398 26019
rect 27420 25999 27422 26019
rect 27540 25999 27542 26019
rect 27564 25999 27566 26019
rect 30553 26014 30556 26019
rect 30564 26014 30566 26019
rect 30563 26000 30566 26014
rect 30529 25999 30563 26000
rect -16257 25995 -11323 25999
rect -16257 25992 -16243 25995
rect -16236 25992 -16233 25995
rect -15324 25975 -15322 25995
rect -15084 25976 -15082 25995
rect -15119 25975 -15061 25976
rect -14999 25975 -14941 25976
rect -14868 25975 -14866 25995
rect -14772 25975 -14770 25995
rect -14508 25975 -14506 25995
rect -14436 25975 -14434 25995
rect -14340 25975 -14338 25995
rect -14255 25990 -14252 25995
rect -14244 25990 -14242 25995
rect -14245 25976 -14242 25990
rect -13980 25975 -13978 25995
rect -13932 25975 -13930 25995
rect -13884 25975 -13882 25995
rect -13788 25975 -13786 25995
rect -13572 25975 -13570 25995
rect -13500 25975 -13498 25995
rect -13356 25975 -13354 25995
rect -13284 25975 -13282 25995
rect -13068 25975 -13066 25995
rect -12828 25975 -12826 25995
rect -12780 25975 -12778 25995
rect -12660 25975 -12658 25995
rect -12564 25975 -12562 25995
rect -12492 25975 -12490 25995
rect -12396 25975 -12394 25995
rect -12348 25975 -12346 25995
rect -12252 25975 -12250 25995
rect -12156 25975 -12154 25995
rect -12060 25975 -12058 25995
rect -11844 25975 -11842 25995
rect -11796 25975 -11794 25995
rect -11676 25975 -11674 25995
rect -11580 25975 -11578 25995
rect -11556 25975 -11554 25995
rect -11508 25975 -11506 25995
rect -11460 25975 -11458 25995
rect -11436 25975 -11434 25995
rect -11412 25975 -11410 25995
rect -11364 25975 -11362 25995
rect -11340 25975 -11338 25995
rect -11337 25992 -11323 25995
rect -11313 25995 30563 25999
rect -11313 25992 -11299 25995
rect -11292 25992 -11289 25995
rect -11196 25975 -11194 25995
rect -11124 25975 -11122 25995
rect -11100 25975 -11098 25995
rect -11028 25975 -11026 25995
rect -11015 25990 -11012 25995
rect -11004 25990 -11002 25995
rect -10799 25990 -10796 25995
rect -10788 25990 -10786 25995
rect -11005 25976 -11002 25990
rect -10789 25976 -10786 25990
rect -10740 25975 -10738 25995
rect -10668 25975 -10666 25995
rect -10644 25975 -10642 25995
rect -9996 25975 -9994 25995
rect -9839 25975 -9781 25976
rect -9708 25975 -9706 25995
rect -9612 25975 -9610 25995
rect -9516 25975 -9514 25995
rect -9468 25975 -9466 25995
rect -9420 25975 -9418 25995
rect -9396 25975 -9394 25995
rect -9383 25990 -9380 25995
rect -9372 25990 -9370 25995
rect -9373 25976 -9370 25990
rect -9300 25975 -9298 25995
rect -9252 25975 -9250 25995
rect -9084 25975 -9082 25995
rect -8988 25975 -8986 25995
rect -8951 25990 -8948 25995
rect -8940 25990 -8938 25995
rect -8941 25976 -8938 25990
rect -8892 25975 -8890 25995
rect -8772 25975 -8770 25995
rect -8604 25975 -8602 25995
rect -8484 25975 -8482 25995
rect -8436 25975 -8434 25995
rect -8388 25975 -8386 25995
rect -8364 25975 -8362 25995
rect -8340 25975 -8338 25995
rect -8268 25975 -8266 25995
rect -8100 25975 -8098 25995
rect -8052 25975 -8050 25995
rect -7932 25975 -7930 25995
rect -7692 25975 -7690 25995
rect -7620 25975 -7618 25995
rect -7524 25975 -7522 25995
rect -7356 25975 -7354 25995
rect -7308 25975 -7306 25995
rect -7212 25975 -7210 25995
rect -7188 25975 -7186 25995
rect -7116 25975 -7114 25995
rect -7068 25975 -7066 25995
rect -6972 25975 -6970 25995
rect -6948 25975 -6946 25995
rect -6876 25975 -6874 25995
rect -6852 25975 -6850 25995
rect -6780 25975 -6778 25995
rect -6756 25975 -6754 25995
rect -6660 25975 -6658 25995
rect -6612 25975 -6610 25995
rect -6516 25975 -6514 25995
rect -6492 25975 -6490 25995
rect -6420 25975 -6418 25995
rect -6396 25975 -6394 25995
rect -6372 25975 -6370 25995
rect -6324 25975 -6322 25995
rect -6156 25975 -6154 25995
rect -6060 25975 -6058 25995
rect -6036 25975 -6034 25995
rect -5940 25976 -5938 25995
rect -5951 25975 -5917 25976
rect -5892 25975 -5890 25995
rect -5652 25975 -5650 25995
rect -5268 25975 -5266 25995
rect -5196 25975 -5194 25995
rect -5172 25975 -5170 25995
rect -5100 25975 -5098 25995
rect -5076 25975 -5074 25995
rect -4980 25975 -4978 25995
rect -4956 25975 -4954 25995
rect -4884 25975 -4882 25995
rect -4860 25975 -4858 25995
rect -4788 25975 -4786 25995
rect -4644 25975 -4642 25995
rect -4548 25975 -4546 25995
rect -4308 25975 -4306 25995
rect -4260 25975 -4258 25995
rect -4223 25990 -4220 25995
rect -4212 25990 -4210 25995
rect -4213 25976 -4210 25990
rect -4164 25975 -4162 25995
rect -4116 25992 -4114 25995
rect -4116 25975 -4113 25992
rect -4020 25975 -4018 25995
rect -3876 25975 -3874 25995
rect -3732 25975 -3730 25995
rect -3588 25975 -3586 25995
rect -3564 25975 -3562 25995
rect -3516 25975 -3514 25995
rect -3492 25975 -3490 25995
rect -3468 25975 -3466 25995
rect -3420 25975 -3418 25995
rect -3324 25975 -3322 25995
rect -3252 25975 -3250 25995
rect -3228 25975 -3226 25995
rect -3156 25975 -3154 25995
rect -3132 25975 -3130 25995
rect -3060 25975 -3058 25995
rect -3012 25975 -3010 25995
rect -2964 25975 -2962 25995
rect -2916 25975 -2914 25995
rect -2892 25975 -2890 25995
rect -2868 25975 -2866 25995
rect -2820 25975 -2818 25995
rect -2796 25975 -2794 25995
rect -2772 25975 -2770 25995
rect -2700 25975 -2698 25995
rect -2676 25975 -2674 25995
rect -2604 25975 -2602 25995
rect -2580 25975 -2578 25995
rect -2364 25975 -2362 25995
rect -2268 25975 -2266 25995
rect -2244 25975 -2242 25995
rect -2172 25975 -2170 25995
rect -2148 25975 -2146 25995
rect -2076 25975 -2074 25995
rect -2052 25975 -2050 25995
rect -1980 25975 -1978 25995
rect -1884 25975 -1882 25995
rect -1836 25975 -1834 25995
rect -1727 25990 -1724 25995
rect -1716 25990 -1714 25995
rect -1717 25976 -1714 25990
rect -1596 25975 -1594 25995
rect -1572 25975 -1570 25995
rect -1476 25975 -1474 25995
rect -1380 25975 -1378 25995
rect -1356 25975 -1354 25995
rect -1308 25975 -1306 25995
rect -1260 25975 -1258 25995
rect -1140 25975 -1138 25995
rect -852 25975 -850 25995
rect -756 25975 -754 25995
rect -708 25975 -706 25995
rect -612 25975 -610 25995
rect -588 25975 -586 25995
rect -540 25975 -538 25995
rect -492 25975 -490 25995
rect -444 25975 -442 25995
rect -396 25975 -394 25995
rect -300 25975 -298 25995
rect -276 25975 -274 25995
rect -228 25975 -226 25995
rect -12 25975 -10 25995
rect 156 25975 158 25995
rect 204 25975 206 25995
rect 228 25975 230 25995
rect 252 25975 254 25995
rect 348 25975 350 25995
rect 468 25975 470 25995
rect 492 25975 494 25995
rect 564 25975 566 25995
rect 588 25975 590 25995
rect 636 25975 638 25995
rect 660 25975 662 25995
rect 732 25975 734 25995
rect 756 25975 758 25995
rect 852 25975 854 25995
rect 1020 25975 1022 25995
rect 1092 25975 1094 25995
rect 1116 25975 1118 25995
rect 1212 25975 1214 25995
rect 1308 25975 1310 25995
rect 1332 25975 1334 25995
rect 1380 25975 1382 25995
rect 1428 25975 1430 25995
rect 1476 25975 1478 25995
rect 1524 25975 1526 25995
rect 1548 25975 1550 25995
rect 1620 25975 1622 25995
rect 1644 25975 1646 25995
rect 1692 25975 1694 25995
rect 1716 25975 1718 25995
rect 1740 25975 1742 25995
rect 1788 25975 1790 25995
rect 1884 25975 1886 25995
rect 1980 25975 1982 25995
rect 2028 25975 2030 25995
rect 2076 25975 2078 25995
rect 2100 25975 2102 25995
rect 2124 25975 2126 25995
rect 2172 25975 2174 25995
rect 2196 25975 2198 25995
rect 2220 25975 2222 25995
rect 2268 25975 2270 25995
rect 2292 25975 2294 25995
rect 2316 25975 2318 25995
rect 2364 25975 2366 25995
rect 2412 25975 2414 25995
rect 2460 25975 2462 25995
rect 2508 25975 2510 25995
rect 2580 25975 2582 25995
rect 2604 25975 2606 25995
rect 2676 25975 2678 25995
rect 2700 25975 2702 25995
rect 2748 25975 2750 25995
rect 2772 25975 2774 25995
rect 2796 25975 2798 25995
rect 2844 25975 2846 25995
rect 2868 25975 2870 25995
rect 2892 25975 2894 25995
rect 2940 25975 2942 25995
rect 3012 25975 3014 25995
rect 3108 25975 3110 25995
rect 3156 25975 3158 25995
rect 3252 25975 3254 25995
rect 3348 25975 3350 25995
rect 3396 25975 3398 25995
rect 3468 25975 3470 25995
rect 3492 25975 3494 25995
rect 3564 25975 3566 25995
rect 3612 25975 3614 25995
rect 3636 25975 3638 25995
rect 3660 25975 3662 25995
rect 3708 25975 3710 25995
rect 3732 25975 3734 25995
rect 3804 25975 3806 25995
rect 3828 25975 3830 25995
rect 3924 25975 3926 25995
rect 4020 25975 4022 25995
rect 4044 25975 4046 25995
rect 4092 25975 4094 25995
rect 4116 25975 4118 25995
rect 4140 25975 4142 25995
rect 4188 25975 4190 25995
rect 4212 25975 4214 25995
rect 4236 25975 4238 25995
rect 4308 25975 4310 25995
rect 4332 25975 4334 25995
rect 4404 25975 4406 25995
rect 4500 25975 4502 25995
rect 4596 25975 4598 25995
rect 4860 25975 4862 25995
rect 4956 25975 4958 25995
rect 4980 25975 4982 25995
rect 5004 25975 5006 25995
rect 5076 25975 5078 25995
rect 5100 25975 5102 25995
rect 5124 25975 5126 25995
rect 5172 25975 5174 25995
rect 5220 25975 5222 25995
rect 5268 25975 5270 25995
rect 5388 25975 5390 25995
rect 5484 25975 5486 25995
rect 5508 25975 5510 25995
rect 5532 25975 5534 25995
rect 5628 25975 5630 25995
rect 5652 25975 5654 25995
rect 5748 25975 5750 25995
rect 5796 25975 5798 25995
rect 5844 25975 5846 25995
rect 5892 25975 5894 25995
rect 6132 25975 6134 25995
rect 6180 25975 6182 25995
rect 6228 25975 6230 25995
rect 6252 25975 6254 25995
rect 6276 25975 6278 25995
rect 6324 25975 6326 25995
rect 6372 25975 6374 25995
rect 6492 25975 6494 25995
rect 6588 25975 6590 25995
rect 6612 25975 6614 25995
rect 6660 25975 6662 25995
rect 6684 25975 6686 25995
rect 6708 25975 6710 25995
rect 6780 25975 6782 25995
rect 6804 25975 6806 25995
rect 6828 25975 6830 25995
rect 6900 25975 6902 25995
rect 6924 25975 6926 25995
rect 7020 25975 7022 25995
rect 7140 25975 7142 25995
rect 7236 25975 7238 25995
rect 7332 25975 7334 25995
rect 7380 25975 7382 25995
rect 7428 25975 7430 25995
rect 7452 25975 7454 25995
rect 7476 25975 7478 25995
rect 7524 25975 7526 25995
rect 7548 25975 7550 25995
rect 7572 25975 7574 25995
rect 7620 25975 7622 25995
rect 7644 25975 7646 25995
rect 7668 25975 7670 25995
rect 7740 25975 7742 25995
rect 7788 25975 7790 25995
rect 7884 25975 7886 25995
rect 7956 25975 7958 25995
rect 7980 25975 7982 25995
rect 8028 25975 8030 25995
rect 8196 25975 8198 25995
rect 8244 25975 8246 25995
rect 8268 25975 8270 25995
rect 8292 25975 8294 25995
rect 8340 25975 8342 25995
rect 8364 25975 8366 25995
rect 8388 25975 8390 25995
rect 8436 25975 8438 25995
rect 8460 25975 8462 25995
rect 8556 25975 8558 25995
rect 8604 25975 8606 25995
rect 8652 25975 8654 25995
rect 8700 25975 8702 25995
rect 8724 25975 8726 25995
rect 8748 25975 8750 25995
rect 8820 25975 8822 25995
rect 8844 25975 8846 25995
rect 8868 25975 8870 25995
rect 9516 25975 9518 25995
rect 9612 25975 9614 25995
rect 9660 25975 9662 25995
rect 9684 25975 9686 25995
rect 9708 25975 9710 25995
rect 9756 25975 9758 25995
rect 9780 25975 9782 25995
rect 9804 25975 9806 25995
rect 9852 25975 9854 25995
rect 9876 25975 9878 25995
rect 9900 25975 9902 25995
rect 9948 25975 9950 25995
rect 9972 25975 9974 25995
rect 9996 25975 9998 25995
rect 10068 25975 10070 25995
rect 10092 25975 10094 25995
rect 10116 25975 10118 25995
rect 10164 25975 10166 25995
rect 10188 25975 10190 25995
rect 10212 25975 10214 25995
rect 10284 25975 10286 25995
rect 10308 25975 10310 25995
rect 10332 25975 10334 25995
rect 10380 25975 10382 25995
rect 10404 25975 10406 25995
rect 10428 25975 10430 25995
rect 10476 25975 10478 25995
rect 10500 25975 10502 25995
rect 10524 25975 10526 25995
rect 10572 25975 10574 25995
rect 10596 25975 10598 25995
rect 10620 25975 10622 25995
rect 10668 25975 10670 25995
rect 10692 25975 10694 25995
rect 10716 25975 10718 25995
rect 10788 25975 10790 25995
rect 10836 25975 10838 25995
rect 10956 25975 10958 25995
rect 11052 25975 11054 25995
rect 11076 25975 11078 25995
rect 11124 25975 11126 25995
rect 11172 25975 11174 25995
rect 11220 25975 11222 25995
rect 11340 25975 11342 25995
rect 11436 25975 11438 25995
rect 11532 25975 11534 25995
rect 11580 25975 11582 25995
rect 11628 25975 11630 25995
rect 11676 25975 11678 25995
rect 11724 25975 11726 25995
rect 11772 25975 11774 25995
rect 11796 25975 11798 25995
rect 11892 25975 11894 25995
rect 11988 25975 11990 25995
rect 12060 25975 12062 25995
rect 12132 25975 12134 25995
rect 12228 25975 12230 25995
rect 12276 25975 12278 25995
rect 12324 25975 12326 25995
rect 12420 25975 12422 25995
rect 12444 25975 12446 25995
rect 12492 25975 12494 25995
rect 12516 25975 12518 25995
rect 12540 25975 12542 25995
rect 12588 25975 12590 25995
rect 12636 25975 12638 25995
rect 12732 25975 12734 25995
rect 12756 25975 12758 25995
rect 12804 25975 12806 25995
rect 12828 25975 12830 25995
rect 12852 25975 12854 25995
rect 12900 25975 12902 25995
rect 12948 25975 12950 25995
rect 13044 25975 13046 25995
rect 13068 25975 13070 25995
rect 13116 25975 13118 25995
rect 13284 25975 13286 25995
rect 13332 25975 13334 25995
rect 13428 25975 13430 25995
rect 13524 25975 13526 25995
rect 13572 25975 13574 25995
rect 13644 25975 13646 25995
rect 13668 25975 13670 25995
rect 13764 25975 13766 25995
rect 13812 25975 13814 25995
rect 13860 25975 13862 25995
rect 13908 25975 13910 25995
rect 13956 25975 13958 25995
rect 14004 25975 14006 25995
rect 14100 25975 14102 25995
rect 14196 25975 14198 25995
rect 14292 25975 14294 25995
rect 15132 25975 15134 25995
rect 15180 25975 15182 25995
rect 15228 25975 15230 25995
rect 15252 25975 15254 25995
rect 15324 25975 15326 25995
rect 15396 25975 15398 25995
rect 15420 25975 15422 25995
rect 15492 25975 15494 25995
rect 15540 25975 15542 25995
rect 15636 25975 15638 25995
rect 15660 25975 15662 25995
rect 15708 25975 15710 25995
rect 15732 25975 15734 25995
rect 15756 25975 15758 25995
rect 15804 25975 15806 25995
rect 15828 25975 15830 25995
rect 15852 25975 15854 25995
rect 15900 25975 15902 25995
rect 15948 25975 15950 25995
rect 15996 25975 15998 25995
rect 16044 25975 16046 25995
rect 16164 25975 16166 25995
rect 16260 25975 16262 25995
rect 16308 25975 16310 25995
rect 16332 25975 16334 25995
rect 16356 25975 16358 25995
rect 16404 25975 16406 25995
rect 16452 25975 16454 25995
rect 16548 25975 16550 25995
rect 16572 25975 16574 25995
rect 16620 25975 16622 25995
rect 16668 25975 16670 25995
rect 16716 25975 16718 25995
rect 16764 25975 16766 25995
rect 16812 25975 16814 25995
rect 16884 25975 16886 25995
rect 16908 25975 16910 25995
rect 16980 25975 16982 25995
rect 17052 25975 17054 25995
rect 17196 25975 17198 25995
rect 17220 25975 17222 25995
rect 17292 25975 17294 25995
rect 17316 25975 17318 25995
rect 18084 25975 18086 25995
rect 18132 25975 18134 25995
rect 18396 25975 18398 25995
rect 18492 25975 18494 25995
rect 18516 25975 18518 25995
rect 18564 25975 18566 25995
rect 18612 25975 18614 25995
rect 18660 25975 18662 25995
rect 18708 25975 18710 25995
rect 18756 25975 18758 25995
rect 18804 25975 18806 25995
rect 18852 25975 18854 25995
rect 18900 25975 18902 25995
rect 18996 25975 18998 25995
rect 19020 25975 19022 25995
rect 19092 25975 19094 25995
rect 19116 25975 19118 25995
rect 19140 25975 19142 25995
rect 19188 25975 19190 25995
rect 19236 25975 19238 25995
rect 19332 25975 19334 25995
rect 19476 25975 19478 25995
rect 19788 25975 19790 25995
rect 19836 25975 19838 25995
rect 19860 25975 19862 25995
rect 19884 25975 19886 25995
rect 19932 25975 19934 25995
rect 19956 25975 19958 25995
rect 19980 25975 19982 25995
rect 20028 25975 20030 25995
rect 20052 25975 20054 25995
rect 20076 25975 20078 25995
rect 20148 25975 20150 25995
rect 20172 25975 20174 25995
rect 20196 25975 20198 25995
rect 20268 25975 20270 25995
rect 20292 25975 20294 25995
rect 20388 25975 20390 25995
rect 20412 25975 20414 25995
rect 20508 25975 20510 25995
rect 20556 25975 20558 25995
rect 20604 25975 20606 25995
rect 20916 25975 20918 25995
rect 20964 25975 20966 25995
rect 21012 25975 21014 25995
rect 21060 25975 21062 25995
rect 21084 25975 21086 25995
rect 21108 25975 21110 25995
rect 21204 25975 21206 25995
rect 21300 25975 21302 25995
rect 21324 25975 21326 25995
rect 21444 25975 21446 25995
rect 21468 25975 21470 25995
rect 21564 25975 21566 25995
rect 21612 25975 21614 25995
rect 21684 25975 21686 25995
rect 21708 25975 21710 25995
rect 21828 25975 21830 25995
rect 21924 25975 21926 25995
rect 22068 25975 22070 25995
rect 22188 25975 22190 25995
rect 22212 25975 22214 25995
rect 22884 25975 22886 25995
rect 22980 25975 22982 25995
rect 23076 25975 23078 25995
rect 23100 25975 23102 25995
rect 23124 25975 23126 25995
rect 23244 25975 23246 25995
rect 23340 25975 23342 25995
rect 23412 25975 23414 25995
rect 23497 25990 23500 25995
rect 23507 25976 23510 25990
rect 23508 25975 23510 25976
rect 23556 25975 23558 25995
rect 23628 25992 23630 25995
rect 23628 25975 23631 25992
rect 23652 25975 23654 25995
rect 23676 25975 23678 25995
rect 23724 25975 23726 25995
rect 23772 25975 23774 25995
rect 23820 25975 23822 25995
rect 23868 25975 23870 25995
rect 23916 25975 23918 25995
rect 24012 25975 24014 25995
rect 24084 25975 24086 25995
rect 24396 25975 24398 25995
rect 24492 25975 24494 25995
rect 24516 25975 24518 25995
rect 24588 25975 24590 25995
rect 24612 25975 24614 25995
rect 24684 25975 24686 25995
rect 24732 25975 24734 25995
rect 24756 25975 24758 25995
rect 24780 25975 24782 25995
rect 24852 25975 24854 25995
rect 24876 25975 24878 25995
rect 24972 25975 24974 25995
rect 24996 25975 24998 25995
rect 25068 25975 25070 25995
rect 25164 25975 25166 25995
rect 25260 25975 25262 25995
rect 25308 25975 25310 25995
rect 25356 25975 25358 25995
rect 25380 25975 25382 25995
rect 25404 25975 25406 25995
rect 25441 25990 25444 25995
rect 25452 25990 25454 25995
rect 25451 25976 25454 25990
rect 25500 25975 25502 25995
rect 25596 25975 25598 25995
rect 27036 25975 27038 25995
rect 27108 25975 27110 25995
rect 27324 25975 27326 25995
rect 27396 25975 27398 25995
rect 27420 25975 27422 25995
rect 27540 25975 27542 25995
rect 27564 25975 27566 25995
rect 29857 25975 29891 25976
rect -17279 25971 23597 25975
rect -17159 25951 -17125 25952
rect -17052 25951 -17050 25971
rect -16836 25951 -16834 25971
rect -16764 25968 -16762 25971
rect -16764 25952 -16761 25968
rect -16799 25951 -16741 25952
rect -16740 25951 -16738 25971
rect -16404 25951 -16402 25971
rect -16380 25951 -16378 25971
rect -16356 25951 -16354 25971
rect -16284 25951 -16282 25971
rect -16260 25951 -16258 25971
rect -15479 25951 -15445 25952
rect -15324 25951 -15322 25971
rect -15321 25968 -15307 25971
rect -15095 25966 -15092 25971
rect -15084 25966 -15082 25971
rect -14999 25966 -14996 25971
rect -14868 25968 -14866 25971
rect -15085 25952 -15082 25966
rect -14989 25952 -14985 25966
rect -14988 25951 -14985 25952
rect -14868 25951 -14865 25968
rect -14772 25951 -14770 25971
rect -14508 25951 -14506 25971
rect -14436 25951 -14434 25971
rect -14340 25951 -14338 25971
rect -14169 25968 -14155 25971
rect -13980 25951 -13978 25971
rect -13932 25951 -13930 25971
rect -13884 25951 -13882 25971
rect -13788 25951 -13786 25971
rect -13607 25951 -13573 25952
rect -13572 25951 -13570 25971
rect -13500 25951 -13498 25971
rect -13356 25951 -13354 25971
rect -13284 25951 -13282 25971
rect -13068 25951 -13066 25971
rect -12828 25951 -12826 25971
rect -12780 25951 -12778 25971
rect -12660 25951 -12658 25971
rect -12564 25951 -12562 25971
rect -12492 25951 -12490 25971
rect -12396 25951 -12394 25971
rect -12348 25951 -12346 25971
rect -12252 25951 -12250 25971
rect -12156 25951 -12154 25971
rect -12060 25951 -12058 25971
rect -11844 25951 -11842 25971
rect -11796 25951 -11794 25971
rect -11676 25951 -11674 25971
rect -11580 25951 -11578 25971
rect -11556 25951 -11554 25971
rect -11508 25951 -11506 25971
rect -11460 25951 -11458 25971
rect -11436 25951 -11434 25971
rect -11412 25951 -11410 25971
rect -11364 25951 -11362 25971
rect -11340 25951 -11338 25971
rect -11196 25951 -11194 25971
rect -11124 25951 -11122 25971
rect -11100 25951 -11098 25971
rect -11028 25951 -11026 25971
rect -10929 25968 -10915 25971
rect -10740 25951 -10738 25971
rect -10713 25968 -10699 25971
rect -10668 25951 -10666 25971
rect -10644 25951 -10642 25971
rect -9996 25951 -9994 25971
rect -9839 25966 -9836 25971
rect -9708 25968 -9706 25971
rect -9829 25952 -9826 25966
rect -9828 25951 -9826 25952
rect -9732 25951 -9729 25968
rect -9708 25951 -9705 25968
rect -9612 25951 -9610 25971
rect -9516 25951 -9514 25971
rect -9468 25951 -9466 25971
rect -9420 25951 -9418 25971
rect -9396 25951 -9394 25971
rect -9300 25951 -9298 25971
rect -9297 25968 -9283 25971
rect -9252 25951 -9250 25971
rect -9084 25951 -9082 25971
rect -8988 25951 -8986 25971
rect -8892 25951 -8890 25971
rect -8865 25968 -8851 25971
rect -8772 25951 -8770 25971
rect -8604 25951 -8602 25971
rect -8484 25951 -8482 25971
rect -8436 25951 -8434 25971
rect -8388 25951 -8386 25971
rect -8364 25951 -8362 25971
rect -8340 25951 -8338 25971
rect -8268 25951 -8266 25971
rect -8100 25951 -8098 25971
rect -8052 25951 -8050 25971
rect -7932 25951 -7930 25971
rect -7692 25951 -7690 25971
rect -7620 25951 -7618 25971
rect -7524 25951 -7522 25971
rect -7356 25951 -7354 25971
rect -7308 25951 -7306 25971
rect -7295 25951 -7261 25952
rect -7212 25951 -7210 25971
rect -7188 25951 -7186 25971
rect -7116 25951 -7114 25971
rect -7068 25951 -7066 25971
rect -6972 25951 -6970 25971
rect -6948 25951 -6946 25971
rect -6876 25951 -6874 25971
rect -6852 25951 -6850 25971
rect -6780 25951 -6778 25971
rect -6756 25951 -6754 25971
rect -6660 25951 -6658 25971
rect -6612 25951 -6610 25971
rect -6516 25951 -6514 25971
rect -6492 25951 -6490 25971
rect -6420 25951 -6418 25971
rect -6396 25951 -6394 25971
rect -6372 25951 -6370 25971
rect -6324 25951 -6322 25971
rect -6156 25951 -6154 25971
rect -6060 25951 -6058 25971
rect -6036 25951 -6034 25971
rect -5951 25966 -5948 25971
rect -5940 25966 -5938 25971
rect -5941 25952 -5938 25966
rect -5892 25951 -5890 25971
rect -5652 25951 -5650 25971
rect -5268 25951 -5266 25971
rect -5196 25951 -5194 25971
rect -5172 25951 -5170 25971
rect -5100 25951 -5098 25971
rect -5076 25951 -5074 25971
rect -4980 25951 -4978 25971
rect -4956 25951 -4954 25971
rect -4884 25951 -4882 25971
rect -4860 25951 -4858 25971
rect -4788 25951 -4786 25971
rect -4644 25951 -4642 25971
rect -4548 25951 -4546 25971
rect -4511 25951 -4453 25952
rect -4308 25951 -4306 25971
rect -4260 25951 -4258 25971
rect -4164 25951 -4162 25971
rect -4137 25968 -4123 25971
rect -4116 25968 -4113 25971
rect -4020 25951 -4018 25971
rect -3876 25951 -3874 25971
rect -3732 25951 -3730 25971
rect -3588 25951 -3586 25971
rect -3564 25951 -3562 25971
rect -3516 25951 -3514 25971
rect -3492 25951 -3490 25971
rect -3468 25951 -3466 25971
rect -3420 25951 -3418 25971
rect -3324 25951 -3322 25971
rect -3252 25951 -3250 25971
rect -3228 25951 -3226 25971
rect -3156 25951 -3154 25971
rect -3132 25951 -3130 25971
rect -3060 25951 -3058 25971
rect -3012 25951 -3010 25971
rect -2964 25951 -2962 25971
rect -2916 25951 -2914 25971
rect -2892 25951 -2890 25971
rect -2868 25951 -2866 25971
rect -2820 25951 -2818 25971
rect -2796 25951 -2794 25971
rect -2772 25951 -2770 25971
rect -2700 25951 -2698 25971
rect -2676 25951 -2674 25971
rect -2604 25951 -2602 25971
rect -2580 25951 -2578 25971
rect -2364 25951 -2362 25971
rect -2268 25951 -2266 25971
rect -2244 25951 -2242 25971
rect -2172 25951 -2170 25971
rect -2148 25951 -2146 25971
rect -2076 25951 -2074 25971
rect -2052 25951 -2050 25971
rect -1980 25951 -1978 25971
rect -1884 25951 -1882 25971
rect -1836 25951 -1834 25971
rect -1641 25968 -1627 25971
rect -1596 25951 -1594 25971
rect -1572 25951 -1570 25971
rect -1476 25951 -1474 25971
rect -1380 25951 -1378 25971
rect -1356 25951 -1354 25971
rect -1308 25951 -1306 25971
rect -1260 25951 -1258 25971
rect -1140 25951 -1138 25971
rect -852 25951 -850 25971
rect -756 25951 -754 25971
rect -708 25951 -706 25971
rect -612 25951 -610 25971
rect -588 25951 -586 25971
rect -540 25951 -538 25971
rect -492 25951 -490 25971
rect -444 25951 -442 25971
rect -396 25951 -394 25971
rect -300 25951 -298 25971
rect -276 25951 -274 25971
rect -228 25951 -226 25971
rect -12 25951 -10 25971
rect 15 25968 29 25971
rect 156 25951 158 25971
rect 204 25951 206 25971
rect 228 25951 230 25971
rect 252 25951 254 25971
rect 348 25951 350 25971
rect 468 25951 470 25971
rect 492 25951 494 25971
rect 564 25951 566 25971
rect 588 25951 590 25971
rect 636 25951 638 25971
rect 660 25951 662 25971
rect 732 25951 734 25971
rect 756 25951 758 25971
rect 852 25951 854 25971
rect 1020 25951 1022 25971
rect 1092 25951 1094 25971
rect 1116 25951 1118 25971
rect 1212 25951 1214 25971
rect 1308 25951 1310 25971
rect 1332 25951 1334 25971
rect 1380 25951 1382 25971
rect 1428 25951 1430 25971
rect 1476 25951 1478 25971
rect 1524 25951 1526 25971
rect 1548 25951 1550 25971
rect 1620 25951 1622 25971
rect 1644 25951 1646 25971
rect 1692 25951 1694 25971
rect 1716 25951 1718 25971
rect 1740 25951 1742 25971
rect 1788 25951 1790 25971
rect 1884 25952 1886 25971
rect 1849 25951 1907 25952
rect 1980 25951 1982 25971
rect 2028 25951 2030 25971
rect 2076 25951 2078 25971
rect 2100 25951 2102 25971
rect 2124 25951 2126 25971
rect 2172 25951 2174 25971
rect 2196 25951 2198 25971
rect 2220 25951 2222 25971
rect 2268 25951 2270 25971
rect 2292 25951 2294 25971
rect 2316 25951 2318 25971
rect 2364 25951 2366 25971
rect 2412 25951 2414 25971
rect 2460 25951 2462 25971
rect 2508 25951 2510 25971
rect 2580 25951 2582 25971
rect 2604 25951 2606 25971
rect 2676 25951 2678 25971
rect 2700 25951 2702 25971
rect 2748 25951 2750 25971
rect 2772 25951 2774 25971
rect 2796 25951 2798 25971
rect 2844 25951 2846 25971
rect 2868 25951 2870 25971
rect 2892 25951 2894 25971
rect 2940 25951 2942 25971
rect 3012 25951 3014 25971
rect 3108 25951 3110 25971
rect 3156 25951 3158 25971
rect 3252 25951 3254 25971
rect 3348 25951 3350 25971
rect 3396 25951 3398 25971
rect 3468 25951 3470 25971
rect 3492 25951 3494 25971
rect 3564 25951 3566 25971
rect 3612 25951 3614 25971
rect 3636 25951 3638 25971
rect 3660 25951 3662 25971
rect 3708 25951 3710 25971
rect 3732 25951 3734 25971
rect 3804 25951 3806 25971
rect 3828 25951 3830 25971
rect 3924 25951 3926 25971
rect 4020 25951 4022 25971
rect 4044 25951 4046 25971
rect 4092 25951 4094 25971
rect 4116 25951 4118 25971
rect 4140 25951 4142 25971
rect 4188 25951 4190 25971
rect 4212 25951 4214 25971
rect 4236 25951 4238 25971
rect 4308 25951 4310 25971
rect 4332 25951 4334 25971
rect 4404 25951 4406 25971
rect 4500 25951 4502 25971
rect 4596 25951 4598 25971
rect 4860 25951 4862 25971
rect 4956 25951 4958 25971
rect 4980 25951 4982 25971
rect 5004 25951 5006 25971
rect 5076 25951 5078 25971
rect 5100 25951 5102 25971
rect 5124 25951 5126 25971
rect 5172 25951 5174 25971
rect 5220 25951 5222 25971
rect 5268 25951 5270 25971
rect 5388 25951 5390 25971
rect 5484 25951 5486 25971
rect 5508 25951 5510 25971
rect 5532 25951 5534 25971
rect 5628 25951 5630 25971
rect 5652 25951 5654 25971
rect 5748 25951 5750 25971
rect 5796 25951 5798 25971
rect 5844 25951 5846 25971
rect 5892 25951 5894 25971
rect 6132 25951 6134 25971
rect 6180 25951 6182 25971
rect 6228 25951 6230 25971
rect 6252 25951 6254 25971
rect 6276 25951 6278 25971
rect 6324 25951 6326 25971
rect 6372 25951 6374 25971
rect 6492 25951 6494 25971
rect 6588 25951 6590 25971
rect 6612 25951 6614 25971
rect 6660 25951 6662 25971
rect 6684 25951 6686 25971
rect 6708 25951 6710 25971
rect 6780 25951 6782 25971
rect 6804 25951 6806 25971
rect 6828 25951 6830 25971
rect 6900 25951 6902 25971
rect 6924 25951 6926 25971
rect 7020 25951 7022 25971
rect 7140 25951 7142 25971
rect 7236 25951 7238 25971
rect 7332 25951 7334 25971
rect 7380 25951 7382 25971
rect 7428 25951 7430 25971
rect 7452 25951 7454 25971
rect 7476 25951 7478 25971
rect 7524 25951 7526 25971
rect 7548 25951 7550 25971
rect 7572 25951 7574 25971
rect 7620 25951 7622 25971
rect 7644 25951 7646 25971
rect 7668 25951 7670 25971
rect 7740 25951 7742 25971
rect 7788 25951 7790 25971
rect 7884 25951 7886 25971
rect 7956 25951 7958 25971
rect 7980 25951 7982 25971
rect 8028 25951 8030 25971
rect 8196 25951 8198 25971
rect 8244 25951 8246 25971
rect 8268 25951 8270 25971
rect 8292 25951 8294 25971
rect 8340 25951 8342 25971
rect 8364 25951 8366 25971
rect 8388 25951 8390 25971
rect 8436 25951 8438 25971
rect 8460 25951 8462 25971
rect 8556 25951 8558 25971
rect 8604 25951 8606 25971
rect 8652 25951 8654 25971
rect 8700 25951 8702 25971
rect 8724 25951 8726 25971
rect 8748 25951 8750 25971
rect 8820 25951 8822 25971
rect 8844 25951 8846 25971
rect 8868 25951 8870 25971
rect 9516 25951 9518 25971
rect 9612 25951 9614 25971
rect 9660 25951 9662 25971
rect 9684 25951 9686 25971
rect 9708 25951 9710 25971
rect 9756 25951 9758 25971
rect 9780 25951 9782 25971
rect 9804 25951 9806 25971
rect 9852 25951 9854 25971
rect 9876 25951 9878 25971
rect 9900 25951 9902 25971
rect 9948 25951 9950 25971
rect 9972 25951 9974 25971
rect 9996 25951 9998 25971
rect 10068 25951 10070 25971
rect 10092 25951 10094 25971
rect 10116 25951 10118 25971
rect 10164 25951 10166 25971
rect 10188 25951 10190 25971
rect 10212 25951 10214 25971
rect 10284 25951 10286 25971
rect 10308 25951 10310 25971
rect 10332 25951 10334 25971
rect 10380 25951 10382 25971
rect 10404 25951 10406 25971
rect 10428 25951 10430 25971
rect 10476 25951 10478 25971
rect 10500 25951 10502 25971
rect 10524 25951 10526 25971
rect 10572 25951 10574 25971
rect 10596 25951 10598 25971
rect 10620 25951 10622 25971
rect 10668 25951 10670 25971
rect 10692 25951 10694 25971
rect 10716 25951 10718 25971
rect 10788 25951 10790 25971
rect 10836 25951 10838 25971
rect 10956 25951 10958 25971
rect 10993 25951 11051 25952
rect 11052 25951 11054 25971
rect 11076 25951 11078 25971
rect 11124 25951 11126 25971
rect 11172 25951 11174 25971
rect 11220 25951 11222 25971
rect 11340 25951 11342 25971
rect 11436 25951 11438 25971
rect 11532 25951 11534 25971
rect 11580 25951 11582 25971
rect 11628 25951 11630 25971
rect 11676 25951 11678 25971
rect 11724 25951 11726 25971
rect 11772 25951 11774 25971
rect 11796 25951 11798 25971
rect 11892 25951 11894 25971
rect 11988 25951 11990 25971
rect 12060 25951 12062 25971
rect 12132 25951 12134 25971
rect 12228 25951 12230 25971
rect 12276 25951 12278 25971
rect 12324 25951 12326 25971
rect 12420 25951 12422 25971
rect 12444 25951 12446 25971
rect 12492 25951 12494 25971
rect 12516 25951 12518 25971
rect 12540 25951 12542 25971
rect 12588 25951 12590 25971
rect 12636 25951 12638 25971
rect 12732 25951 12734 25971
rect 12756 25951 12758 25971
rect 12804 25951 12806 25971
rect 12828 25951 12830 25971
rect 12852 25951 12854 25971
rect 12900 25951 12902 25971
rect 12948 25951 12950 25971
rect 13044 25951 13046 25971
rect 13068 25951 13070 25971
rect 13116 25951 13118 25971
rect 13284 25951 13286 25971
rect 13332 25951 13334 25971
rect 13428 25952 13430 25971
rect 13393 25951 13451 25952
rect 13524 25951 13526 25971
rect 13572 25951 13574 25971
rect 13644 25951 13646 25971
rect 13668 25951 13670 25971
rect 13764 25951 13766 25971
rect 13812 25951 13814 25971
rect 13860 25951 13862 25971
rect 13908 25951 13910 25971
rect 13956 25951 13958 25971
rect 14004 25951 14006 25971
rect 14100 25951 14102 25971
rect 14196 25951 14198 25971
rect 14292 25951 14294 25971
rect 14343 25968 14357 25971
rect 15132 25951 15134 25971
rect 15180 25951 15182 25971
rect 15228 25951 15230 25971
rect 15252 25951 15254 25971
rect 15324 25951 15326 25971
rect 15396 25951 15398 25971
rect 15420 25951 15422 25971
rect 15492 25951 15494 25971
rect 15540 25951 15542 25971
rect 15636 25951 15638 25971
rect 15660 25951 15662 25971
rect 15708 25951 15710 25971
rect 15732 25951 15734 25971
rect 15756 25951 15758 25971
rect 15804 25951 15806 25971
rect 15828 25951 15830 25971
rect 15852 25951 15854 25971
rect 15900 25951 15902 25971
rect 15948 25951 15950 25971
rect 15996 25951 15998 25971
rect 16044 25951 16046 25971
rect 16164 25951 16166 25971
rect 16260 25951 16262 25971
rect 16308 25951 16310 25971
rect 16332 25951 16334 25971
rect 16356 25951 16358 25971
rect 16404 25951 16406 25971
rect 16452 25951 16454 25971
rect 16548 25951 16550 25971
rect 16572 25951 16574 25971
rect 16620 25951 16622 25971
rect 16668 25951 16670 25971
rect 16716 25951 16718 25971
rect 16764 25951 16766 25971
rect 16812 25951 16814 25971
rect 16884 25951 16886 25971
rect 16908 25951 16910 25971
rect 16980 25951 16982 25971
rect 17052 25951 17054 25971
rect 17196 25951 17198 25971
rect 17220 25951 17222 25971
rect 17292 25951 17294 25971
rect 17316 25951 17318 25971
rect 18084 25951 18086 25971
rect 18132 25951 18134 25971
rect 18396 25951 18398 25971
rect 18492 25951 18494 25971
rect 18516 25951 18518 25971
rect 18564 25951 18566 25971
rect 18612 25951 18614 25971
rect 18660 25951 18662 25971
rect 18708 25951 18710 25971
rect 18756 25951 18758 25971
rect 18804 25951 18806 25971
rect 18852 25951 18854 25971
rect 18900 25951 18902 25971
rect 18996 25951 18998 25971
rect 19020 25951 19022 25971
rect 19092 25951 19094 25971
rect 19116 25951 19118 25971
rect 19140 25951 19142 25971
rect 19188 25951 19190 25971
rect 19236 25951 19238 25971
rect 19332 25951 19334 25971
rect 19476 25951 19478 25971
rect 19788 25951 19790 25971
rect 19836 25951 19838 25971
rect 19860 25951 19862 25971
rect 19884 25951 19886 25971
rect 19932 25951 19934 25971
rect 19956 25951 19958 25971
rect 19980 25951 19982 25971
rect 20028 25951 20030 25971
rect 20052 25951 20054 25971
rect 20076 25951 20078 25971
rect 20148 25951 20150 25971
rect 20172 25951 20174 25971
rect 20196 25951 20198 25971
rect 20268 25951 20270 25971
rect 20292 25951 20294 25971
rect 20388 25951 20390 25971
rect 20412 25951 20414 25971
rect 20508 25951 20510 25971
rect 20556 25951 20558 25971
rect 20604 25951 20606 25971
rect 20916 25951 20918 25971
rect 20964 25951 20966 25971
rect 21012 25951 21014 25971
rect 21060 25951 21062 25971
rect 21084 25951 21086 25971
rect 21108 25951 21110 25971
rect 21204 25951 21206 25971
rect 21300 25951 21302 25971
rect 21324 25951 21326 25971
rect 21444 25951 21446 25971
rect 21468 25951 21470 25971
rect 21564 25951 21566 25971
rect 21612 25951 21614 25971
rect 21684 25951 21686 25971
rect 21708 25951 21710 25971
rect 21828 25951 21830 25971
rect 21924 25951 21926 25971
rect 22068 25951 22070 25971
rect 22188 25951 22190 25971
rect 22212 25951 22214 25971
rect 22503 25968 22517 25971
rect 22884 25951 22886 25971
rect 22980 25951 22982 25971
rect 23076 25951 23078 25971
rect 23100 25951 23102 25971
rect 23124 25951 23126 25971
rect 23244 25951 23246 25971
rect 23340 25951 23342 25971
rect 23412 25951 23414 25971
rect 23508 25951 23510 25971
rect 23556 25951 23558 25971
rect 23583 25968 23597 25971
rect 23607 25971 25517 25975
rect 23607 25968 23621 25971
rect 23628 25968 23631 25971
rect 23652 25951 23654 25971
rect 23676 25951 23678 25971
rect 23724 25951 23726 25971
rect 23772 25951 23774 25971
rect 23820 25951 23822 25971
rect 23868 25952 23870 25971
rect 23833 25951 23891 25952
rect 23916 25951 23918 25971
rect 24012 25951 24014 25971
rect 24084 25951 24086 25971
rect 24396 25951 24398 25971
rect 24492 25951 24494 25971
rect 24516 25951 24518 25971
rect 24588 25951 24590 25971
rect 24612 25951 24614 25971
rect 24684 25951 24686 25971
rect 24732 25951 24734 25971
rect 24756 25951 24758 25971
rect 24780 25951 24782 25971
rect 24852 25951 24854 25971
rect 24876 25951 24878 25971
rect 24972 25951 24974 25971
rect 24996 25951 24998 25971
rect 25068 25951 25070 25971
rect 25164 25951 25166 25971
rect 25260 25951 25262 25971
rect 25308 25951 25310 25971
rect 25356 25951 25358 25971
rect 25380 25951 25382 25971
rect 25404 25951 25406 25971
rect 25500 25951 25502 25971
rect 25503 25968 25517 25971
rect 25527 25971 29891 25975
rect 30457 25975 30491 25976
rect 30505 25975 30539 25976
rect 30457 25971 30539 25975
rect 25527 25968 25541 25971
rect 25596 25951 25598 25971
rect 27036 25951 27038 25971
rect 27108 25951 27110 25971
rect 27324 25951 27326 25971
rect 27396 25951 27398 25971
rect 27420 25951 27422 25971
rect 27540 25951 27542 25971
rect 27564 25951 27566 25971
rect 28225 25951 28259 25952
rect 28945 25951 28979 25952
rect -17159 25947 -15019 25951
rect -17052 25944 -17050 25947
rect -17052 25928 -17049 25944
rect -17063 25927 -17029 25928
rect -16836 25927 -16834 25947
rect -16785 25944 -16771 25947
rect -16764 25944 -16761 25947
rect -16740 25927 -16738 25947
rect -16692 25927 -16689 25944
rect -16535 25927 -16477 25928
rect -16404 25927 -16402 25947
rect -16380 25927 -16378 25947
rect -16356 25927 -16354 25947
rect -16284 25927 -16282 25947
rect -16260 25927 -16258 25947
rect -15324 25927 -15322 25947
rect -15033 25944 -15019 25947
rect -15009 25947 -14899 25951
rect -15009 25944 -14995 25947
rect -14988 25944 -14985 25947
rect -14913 25944 -14899 25947
rect -14889 25947 -9739 25951
rect -14889 25944 -14875 25947
rect -14868 25944 -14865 25947
rect -14772 25927 -14770 25947
rect -14508 25927 -14506 25947
rect -14436 25927 -14434 25947
rect -14340 25927 -14338 25947
rect -13980 25927 -13978 25947
rect -13932 25927 -13930 25947
rect -13884 25927 -13882 25947
rect -13788 25927 -13786 25947
rect -13572 25927 -13570 25947
rect -13500 25944 -13498 25947
rect -13500 25927 -13497 25944
rect -13356 25927 -13354 25947
rect -13284 25927 -13282 25947
rect -13068 25927 -13066 25947
rect -12828 25927 -12826 25947
rect -12780 25927 -12778 25947
rect -12660 25927 -12658 25947
rect -12564 25927 -12562 25947
rect -12492 25927 -12490 25947
rect -12396 25927 -12394 25947
rect -12348 25927 -12346 25947
rect -12252 25927 -12250 25947
rect -12156 25927 -12154 25947
rect -12060 25927 -12058 25947
rect -11844 25927 -11842 25947
rect -11796 25927 -11794 25947
rect -11676 25927 -11674 25947
rect -11580 25927 -11578 25947
rect -11556 25927 -11554 25947
rect -11508 25927 -11506 25947
rect -11460 25927 -11458 25947
rect -11436 25927 -11434 25947
rect -11412 25927 -11410 25947
rect -11364 25927 -11362 25947
rect -11340 25927 -11338 25947
rect -11196 25927 -11194 25947
rect -11124 25927 -11122 25947
rect -11100 25927 -11098 25947
rect -11028 25927 -11026 25947
rect -10740 25927 -10738 25947
rect -10668 25927 -10666 25947
rect -10644 25927 -10642 25947
rect -9996 25927 -9994 25947
rect -9828 25927 -9826 25947
rect -9753 25944 -9739 25947
rect -9732 25947 28979 25951
rect -9732 25944 -9715 25947
rect -9708 25944 -9705 25947
rect -9732 25927 -9730 25944
rect -9612 25927 -9610 25947
rect -9516 25927 -9514 25947
rect -9468 25927 -9466 25947
rect -9420 25927 -9418 25947
rect -9396 25927 -9394 25947
rect -9300 25927 -9298 25947
rect -9252 25927 -9250 25947
rect -9084 25927 -9082 25947
rect -8988 25927 -8986 25947
rect -8892 25927 -8890 25947
rect -8772 25927 -8770 25947
rect -8604 25927 -8602 25947
rect -8484 25927 -8482 25947
rect -8436 25927 -8434 25947
rect -8388 25927 -8386 25947
rect -8364 25927 -8362 25947
rect -8340 25927 -8338 25947
rect -8268 25927 -8266 25947
rect -8100 25927 -8098 25947
rect -8052 25927 -8050 25947
rect -7932 25927 -7930 25947
rect -7692 25927 -7690 25947
rect -7620 25927 -7618 25947
rect -7524 25927 -7522 25947
rect -7356 25927 -7354 25947
rect -7308 25927 -7306 25947
rect -7212 25927 -7210 25947
rect -7188 25944 -7186 25947
rect -7188 25927 -7185 25944
rect -7116 25927 -7114 25947
rect -7068 25927 -7066 25947
rect -6972 25927 -6970 25947
rect -6948 25927 -6946 25947
rect -6876 25927 -6874 25947
rect -6852 25927 -6850 25947
rect -6780 25927 -6778 25947
rect -6756 25927 -6754 25947
rect -6660 25927 -6658 25947
rect -6612 25927 -6610 25947
rect -6516 25927 -6514 25947
rect -6492 25927 -6490 25947
rect -6420 25927 -6418 25947
rect -6396 25927 -6394 25947
rect -6372 25927 -6370 25947
rect -6324 25927 -6322 25947
rect -6156 25927 -6154 25947
rect -6060 25927 -6058 25947
rect -6036 25927 -6034 25947
rect -5892 25927 -5890 25947
rect -5865 25944 -5851 25947
rect -5652 25927 -5650 25947
rect -5268 25927 -5266 25947
rect -5196 25927 -5194 25947
rect -5172 25927 -5170 25947
rect -5100 25927 -5098 25947
rect -5076 25927 -5074 25947
rect -4980 25927 -4978 25947
rect -4956 25927 -4954 25947
rect -4884 25927 -4882 25947
rect -4860 25927 -4858 25947
rect -4788 25927 -4786 25947
rect -4644 25927 -4642 25947
rect -4548 25927 -4546 25947
rect -4511 25942 -4508 25947
rect -4501 25928 -4498 25942
rect -4500 25927 -4498 25928
rect -4404 25927 -4401 25944
rect -4308 25927 -4306 25947
rect -4260 25927 -4258 25947
rect -4164 25927 -4162 25947
rect -4020 25927 -4018 25947
rect -3876 25927 -3874 25947
rect -3732 25927 -3730 25947
rect -3588 25927 -3586 25947
rect -3564 25927 -3562 25947
rect -3516 25927 -3514 25947
rect -3492 25927 -3490 25947
rect -3468 25927 -3466 25947
rect -3420 25927 -3418 25947
rect -3324 25927 -3322 25947
rect -3252 25927 -3250 25947
rect -3228 25927 -3226 25947
rect -3156 25927 -3154 25947
rect -3132 25927 -3130 25947
rect -3060 25927 -3058 25947
rect -3012 25927 -3010 25947
rect -2964 25927 -2962 25947
rect -2916 25927 -2914 25947
rect -2892 25927 -2890 25947
rect -2868 25927 -2866 25947
rect -2820 25927 -2818 25947
rect -2796 25927 -2794 25947
rect -2772 25927 -2770 25947
rect -2700 25927 -2698 25947
rect -2676 25927 -2674 25947
rect -2604 25927 -2602 25947
rect -2580 25927 -2578 25947
rect -2364 25927 -2362 25947
rect -2268 25927 -2266 25947
rect -2244 25927 -2242 25947
rect -2172 25927 -2170 25947
rect -2148 25927 -2146 25947
rect -2076 25927 -2074 25947
rect -2052 25927 -2050 25947
rect -1980 25927 -1978 25947
rect -1884 25927 -1882 25947
rect -1836 25927 -1834 25947
rect -1596 25927 -1594 25947
rect -1572 25927 -1570 25947
rect -1476 25927 -1474 25947
rect -1380 25927 -1378 25947
rect -1356 25927 -1354 25947
rect -1308 25927 -1306 25947
rect -1260 25927 -1258 25947
rect -1140 25927 -1138 25947
rect -852 25927 -850 25947
rect -756 25927 -754 25947
rect -708 25927 -706 25947
rect -612 25927 -610 25947
rect -588 25927 -586 25947
rect -540 25927 -538 25947
rect -492 25927 -490 25947
rect -444 25927 -442 25947
rect -396 25927 -394 25947
rect -300 25927 -298 25947
rect -276 25927 -274 25947
rect -228 25927 -226 25947
rect -12 25927 -10 25947
rect 156 25927 158 25947
rect 204 25927 206 25947
rect 228 25927 230 25947
rect 252 25927 254 25947
rect 348 25927 350 25947
rect 468 25927 470 25947
rect 492 25927 494 25947
rect 564 25927 566 25947
rect 588 25927 590 25947
rect 636 25927 638 25947
rect 660 25927 662 25947
rect 732 25927 734 25947
rect 756 25927 758 25947
rect 852 25927 854 25947
rect 1020 25927 1022 25947
rect 1092 25927 1094 25947
rect 1116 25927 1118 25947
rect 1212 25927 1214 25947
rect 1308 25927 1310 25947
rect 1332 25927 1334 25947
rect 1380 25927 1382 25947
rect 1428 25927 1430 25947
rect 1476 25927 1478 25947
rect 1524 25927 1526 25947
rect 1548 25927 1550 25947
rect 1620 25927 1622 25947
rect 1644 25927 1646 25947
rect 1692 25927 1694 25947
rect 1716 25927 1718 25947
rect 1740 25927 1742 25947
rect 1788 25927 1790 25947
rect 1873 25942 1876 25947
rect 1884 25942 1886 25947
rect 1883 25928 1886 25942
rect 1980 25944 1982 25947
rect 1980 25927 1983 25944
rect 2028 25927 2030 25947
rect 2076 25927 2078 25947
rect 2100 25927 2102 25947
rect 2124 25927 2126 25947
rect 2172 25927 2174 25947
rect 2196 25927 2198 25947
rect 2220 25927 2222 25947
rect 2268 25927 2270 25947
rect 2292 25927 2294 25947
rect 2316 25927 2318 25947
rect 2364 25927 2366 25947
rect 2412 25927 2414 25947
rect 2460 25927 2462 25947
rect 2508 25927 2510 25947
rect 2580 25927 2582 25947
rect 2604 25927 2606 25947
rect 2676 25927 2678 25947
rect 2700 25927 2702 25947
rect 2748 25927 2750 25947
rect 2772 25927 2774 25947
rect 2796 25927 2798 25947
rect 2844 25927 2846 25947
rect 2868 25927 2870 25947
rect 2892 25927 2894 25947
rect 2940 25927 2942 25947
rect 3012 25927 3014 25947
rect 3108 25927 3110 25947
rect 3156 25927 3158 25947
rect 3252 25927 3254 25947
rect 3348 25927 3350 25947
rect 3396 25927 3398 25947
rect 3468 25927 3470 25947
rect 3492 25927 3494 25947
rect 3564 25927 3566 25947
rect 3612 25927 3614 25947
rect 3636 25927 3638 25947
rect 3660 25927 3662 25947
rect 3708 25927 3710 25947
rect 3732 25927 3734 25947
rect 3804 25927 3806 25947
rect 3828 25927 3830 25947
rect 3924 25927 3926 25947
rect 4020 25927 4022 25947
rect 4044 25927 4046 25947
rect 4092 25927 4094 25947
rect 4116 25927 4118 25947
rect 4140 25927 4142 25947
rect 4188 25927 4190 25947
rect 4212 25927 4214 25947
rect 4236 25927 4238 25947
rect 4308 25927 4310 25947
rect 4332 25927 4334 25947
rect 4404 25927 4406 25947
rect 4500 25927 4502 25947
rect 4596 25927 4598 25947
rect 4860 25927 4862 25947
rect 4956 25927 4958 25947
rect 4980 25927 4982 25947
rect 5004 25927 5006 25947
rect 5076 25927 5078 25947
rect 5100 25927 5102 25947
rect 5124 25927 5126 25947
rect 5172 25927 5174 25947
rect 5220 25927 5222 25947
rect 5268 25927 5270 25947
rect 5388 25927 5390 25947
rect 5484 25927 5486 25947
rect 5508 25927 5510 25947
rect 5532 25927 5534 25947
rect 5628 25927 5630 25947
rect 5652 25927 5654 25947
rect 5748 25927 5750 25947
rect 5796 25927 5798 25947
rect 5844 25927 5846 25947
rect 5892 25927 5894 25947
rect 6132 25927 6134 25947
rect 6180 25927 6182 25947
rect 6228 25927 6230 25947
rect 6252 25927 6254 25947
rect 6276 25927 6278 25947
rect 6324 25927 6326 25947
rect 6372 25927 6374 25947
rect 6492 25927 6494 25947
rect 6588 25927 6590 25947
rect 6612 25927 6614 25947
rect 6660 25927 6662 25947
rect 6684 25927 6686 25947
rect 6708 25927 6710 25947
rect 6780 25927 6782 25947
rect 6804 25927 6806 25947
rect 6828 25927 6830 25947
rect 6900 25927 6902 25947
rect 6924 25927 6926 25947
rect 7020 25927 7022 25947
rect 7140 25927 7142 25947
rect 7236 25927 7238 25947
rect 7332 25927 7334 25947
rect 7380 25927 7382 25947
rect 7428 25927 7430 25947
rect 7452 25927 7454 25947
rect 7476 25927 7478 25947
rect 7524 25927 7526 25947
rect 7548 25927 7550 25947
rect 7572 25927 7574 25947
rect 7620 25927 7622 25947
rect 7644 25927 7646 25947
rect 7668 25927 7670 25947
rect 7740 25927 7742 25947
rect 7788 25927 7790 25947
rect 7884 25927 7886 25947
rect 7956 25927 7958 25947
rect 7980 25927 7982 25947
rect 8028 25927 8030 25947
rect 8196 25927 8198 25947
rect 8244 25927 8246 25947
rect 8268 25927 8270 25947
rect 8292 25927 8294 25947
rect 8340 25927 8342 25947
rect 8364 25927 8366 25947
rect 8388 25927 8390 25947
rect 8436 25927 8438 25947
rect 8460 25927 8462 25947
rect 8556 25927 8558 25947
rect 8604 25927 8606 25947
rect 8652 25927 8654 25947
rect 8700 25927 8702 25947
rect 8724 25927 8726 25947
rect 8748 25927 8750 25947
rect 8820 25927 8822 25947
rect 8844 25927 8846 25947
rect 8868 25927 8870 25947
rect 9516 25927 9518 25947
rect 9612 25927 9614 25947
rect 9660 25927 9662 25947
rect 9684 25927 9686 25947
rect 9708 25927 9710 25947
rect 9756 25927 9758 25947
rect 9780 25927 9782 25947
rect 9804 25927 9806 25947
rect 9852 25927 9854 25947
rect 9876 25927 9878 25947
rect 9900 25927 9902 25947
rect 9948 25927 9950 25947
rect 9972 25927 9974 25947
rect 9996 25927 9998 25947
rect 10068 25927 10070 25947
rect 10092 25927 10094 25947
rect 10116 25927 10118 25947
rect 10164 25927 10166 25947
rect 10188 25927 10190 25947
rect 10212 25927 10214 25947
rect 10284 25927 10286 25947
rect 10308 25927 10310 25947
rect 10332 25927 10334 25947
rect 10380 25927 10382 25947
rect 10404 25927 10406 25947
rect 10428 25927 10430 25947
rect 10476 25927 10478 25947
rect 10500 25927 10502 25947
rect 10524 25927 10526 25947
rect 10572 25927 10574 25947
rect 10596 25927 10598 25947
rect 10620 25927 10622 25947
rect 10668 25927 10670 25947
rect 10692 25927 10694 25947
rect 10716 25927 10718 25947
rect 10788 25927 10790 25947
rect 10836 25927 10838 25947
rect 10956 25927 10958 25947
rect 10993 25942 10996 25947
rect 11003 25928 11006 25942
rect 11004 25927 11006 25928
rect 11052 25927 11054 25947
rect 11076 25927 11078 25947
rect 11124 25944 11126 25947
rect 11100 25927 11103 25944
rect 11124 25927 11127 25944
rect 11172 25927 11174 25947
rect 11220 25927 11222 25947
rect 11340 25927 11342 25947
rect 11436 25927 11438 25947
rect 11532 25927 11534 25947
rect 11580 25927 11582 25947
rect 11628 25927 11630 25947
rect 11676 25927 11678 25947
rect 11724 25927 11726 25947
rect 11772 25927 11774 25947
rect 11796 25927 11798 25947
rect 11892 25927 11894 25947
rect 11988 25927 11990 25947
rect 12060 25927 12062 25947
rect 12132 25927 12134 25947
rect 12228 25927 12230 25947
rect 12276 25927 12278 25947
rect 12324 25927 12326 25947
rect 12420 25927 12422 25947
rect 12444 25927 12446 25947
rect 12492 25927 12494 25947
rect 12516 25927 12518 25947
rect 12540 25927 12542 25947
rect 12588 25927 12590 25947
rect 12636 25927 12638 25947
rect 12732 25927 12734 25947
rect 12756 25927 12758 25947
rect 12804 25927 12806 25947
rect 12828 25927 12830 25947
rect 12852 25927 12854 25947
rect 12900 25927 12902 25947
rect 12948 25927 12950 25947
rect 13044 25927 13046 25947
rect 13068 25927 13070 25947
rect 13116 25927 13118 25947
rect 13284 25927 13286 25947
rect 13332 25927 13334 25947
rect 13417 25942 13420 25947
rect 13428 25942 13430 25947
rect 13427 25928 13430 25942
rect 13524 25944 13526 25947
rect 13524 25927 13527 25944
rect 13572 25927 13574 25947
rect 13644 25927 13646 25947
rect 13668 25927 13670 25947
rect 13764 25927 13766 25947
rect 13812 25927 13814 25947
rect 13860 25927 13862 25947
rect 13908 25927 13910 25947
rect 13956 25927 13958 25947
rect 14004 25927 14006 25947
rect 14100 25927 14102 25947
rect 14196 25927 14198 25947
rect 14292 25927 14294 25947
rect 15132 25927 15134 25947
rect 15180 25927 15182 25947
rect 15228 25927 15230 25947
rect 15252 25927 15254 25947
rect 15324 25927 15326 25947
rect 15396 25927 15398 25947
rect 15420 25927 15422 25947
rect 15492 25927 15494 25947
rect 15540 25927 15542 25947
rect 15636 25927 15638 25947
rect 15660 25927 15662 25947
rect 15708 25927 15710 25947
rect 15732 25927 15734 25947
rect 15756 25927 15758 25947
rect 15804 25927 15806 25947
rect 15828 25927 15830 25947
rect 15852 25927 15854 25947
rect 15900 25927 15902 25947
rect 15948 25927 15950 25947
rect 15996 25927 15998 25947
rect 16044 25927 16046 25947
rect 16164 25927 16166 25947
rect 16260 25927 16262 25947
rect 16308 25927 16310 25947
rect 16332 25927 16334 25947
rect 16356 25927 16358 25947
rect 16404 25927 16406 25947
rect 16452 25927 16454 25947
rect 16548 25927 16550 25947
rect 16572 25927 16574 25947
rect 16620 25927 16622 25947
rect 16668 25927 16670 25947
rect 16716 25927 16718 25947
rect 16764 25927 16766 25947
rect 16812 25927 16814 25947
rect 16884 25927 16886 25947
rect 16908 25927 16910 25947
rect 16980 25927 16982 25947
rect 17052 25927 17054 25947
rect 17196 25927 17198 25947
rect 17220 25927 17222 25947
rect 17292 25927 17294 25947
rect 17316 25927 17318 25947
rect 18084 25927 18086 25947
rect 18132 25927 18134 25947
rect 18396 25927 18398 25947
rect 18492 25927 18494 25947
rect 18516 25927 18518 25947
rect 18564 25927 18566 25947
rect 18612 25927 18614 25947
rect 18660 25927 18662 25947
rect 18708 25927 18710 25947
rect 18756 25927 18758 25947
rect 18804 25927 18806 25947
rect 18852 25927 18854 25947
rect 18900 25927 18902 25947
rect 18996 25927 18998 25947
rect 19020 25927 19022 25947
rect 19092 25927 19094 25947
rect 19116 25927 19118 25947
rect 19140 25927 19142 25947
rect 19188 25927 19190 25947
rect 19236 25927 19238 25947
rect 19332 25927 19334 25947
rect 19476 25927 19478 25947
rect 19788 25927 19790 25947
rect 19836 25927 19838 25947
rect 19860 25927 19862 25947
rect 19884 25927 19886 25947
rect 19932 25927 19934 25947
rect 19956 25927 19958 25947
rect 19980 25927 19982 25947
rect 20028 25927 20030 25947
rect 20052 25927 20054 25947
rect 20076 25927 20078 25947
rect 20148 25927 20150 25947
rect 20172 25927 20174 25947
rect 20196 25927 20198 25947
rect 20268 25927 20270 25947
rect 20292 25927 20294 25947
rect 20388 25927 20390 25947
rect 20412 25927 20414 25947
rect 20508 25927 20510 25947
rect 20556 25927 20558 25947
rect 20604 25927 20606 25947
rect 20916 25927 20918 25947
rect 20964 25927 20966 25947
rect 21012 25927 21014 25947
rect 21060 25927 21062 25947
rect 21084 25927 21086 25947
rect 21108 25927 21110 25947
rect 21204 25927 21206 25947
rect 21300 25927 21302 25947
rect 21324 25927 21326 25947
rect 21444 25927 21446 25947
rect 21468 25927 21470 25947
rect 21564 25927 21566 25947
rect 21612 25927 21614 25947
rect 21684 25927 21686 25947
rect 21708 25927 21710 25947
rect 21828 25927 21830 25947
rect 21924 25927 21926 25947
rect 22068 25927 22070 25947
rect 22188 25927 22190 25947
rect 22212 25927 22214 25947
rect 22884 25927 22886 25947
rect 22980 25927 22982 25947
rect 23076 25927 23078 25947
rect 23100 25927 23102 25947
rect 23124 25927 23126 25947
rect 23244 25927 23246 25947
rect 23340 25927 23342 25947
rect 23412 25927 23414 25947
rect 23508 25927 23510 25947
rect 23556 25927 23558 25947
rect 23652 25927 23654 25947
rect 23676 25927 23678 25947
rect 23724 25927 23726 25947
rect 23772 25927 23774 25947
rect 23820 25927 23822 25947
rect 23857 25942 23860 25947
rect 23868 25942 23870 25947
rect 23867 25928 23870 25942
rect 23916 25927 23918 25947
rect 24012 25927 24014 25947
rect 24084 25927 24086 25947
rect 24396 25927 24398 25947
rect 24492 25927 24494 25947
rect 24516 25927 24518 25947
rect 24588 25927 24590 25947
rect 24612 25927 24614 25947
rect 24684 25927 24686 25947
rect 24732 25927 24734 25947
rect 24756 25927 24758 25947
rect 24780 25927 24782 25947
rect 24852 25927 24854 25947
rect 24876 25927 24878 25947
rect 24972 25927 24974 25947
rect 24996 25927 24998 25947
rect 25068 25927 25070 25947
rect 25164 25927 25166 25947
rect 25260 25927 25262 25947
rect 25308 25927 25310 25947
rect 25356 25927 25358 25947
rect 25380 25927 25382 25947
rect 25404 25927 25406 25947
rect 25500 25927 25502 25947
rect 25596 25927 25598 25947
rect 27036 25927 27038 25947
rect 27108 25927 27110 25947
rect 27324 25927 27326 25947
rect 27396 25927 27398 25947
rect 27420 25927 27422 25947
rect 27540 25927 27542 25947
rect 27564 25927 27566 25947
rect 28417 25927 28451 25928
rect -17063 25923 -16699 25927
rect -17063 25920 -17059 25923
rect -17052 25920 -17049 25923
rect -16943 25903 -16909 25904
rect -16836 25903 -16834 25923
rect -16740 25903 -16738 25923
rect -16713 25920 -16699 25923
rect -16692 25923 -4411 25927
rect -16692 25920 -16675 25923
rect -16692 25903 -16690 25920
rect -16535 25918 -16532 25923
rect -16404 25920 -16402 25923
rect -16525 25904 -16522 25918
rect -16524 25903 -16522 25904
rect -16511 25903 -16453 25904
rect -16404 25903 -16401 25920
rect -16380 25903 -16378 25923
rect -16356 25903 -16354 25923
rect -16284 25903 -16282 25923
rect -16260 25903 -16258 25923
rect -15393 25920 -15379 25923
rect -15324 25903 -15322 25923
rect -14772 25903 -14770 25923
rect -14508 25903 -14506 25923
rect -14436 25903 -14434 25923
rect -14340 25903 -14338 25923
rect -13980 25903 -13978 25923
rect -13932 25903 -13930 25923
rect -13884 25903 -13882 25923
rect -13788 25903 -13786 25923
rect -13572 25903 -13570 25923
rect -13521 25920 -13507 25923
rect -13500 25920 -13497 25923
rect -13356 25903 -13354 25923
rect -13284 25903 -13282 25923
rect -13068 25903 -13066 25923
rect -12828 25903 -12826 25923
rect -12780 25903 -12778 25923
rect -12660 25903 -12658 25923
rect -12564 25903 -12562 25923
rect -12492 25903 -12490 25923
rect -12396 25903 -12394 25923
rect -12348 25903 -12346 25923
rect -12252 25903 -12250 25923
rect -12156 25903 -12154 25923
rect -12060 25903 -12058 25923
rect -11844 25903 -11842 25923
rect -11796 25903 -11794 25923
rect -11676 25903 -11674 25923
rect -11580 25903 -11578 25923
rect -11556 25903 -11554 25923
rect -11508 25903 -11506 25923
rect -11460 25903 -11458 25923
rect -11436 25903 -11434 25923
rect -11412 25903 -11410 25923
rect -11364 25903 -11362 25923
rect -11340 25903 -11338 25923
rect -11196 25903 -11194 25923
rect -11124 25903 -11122 25923
rect -11100 25903 -11098 25923
rect -11028 25903 -11026 25923
rect -10740 25903 -10738 25923
rect -10668 25903 -10666 25923
rect -10644 25903 -10642 25923
rect -9996 25903 -9994 25923
rect -9828 25903 -9826 25923
rect -9732 25903 -9730 25923
rect -9612 25903 -9610 25923
rect -9516 25903 -9514 25923
rect -9468 25903 -9466 25923
rect -9420 25903 -9418 25923
rect -9396 25903 -9394 25923
rect -9300 25903 -9298 25923
rect -9252 25903 -9250 25923
rect -9084 25903 -9082 25923
rect -8988 25903 -8986 25923
rect -8892 25903 -8890 25923
rect -8772 25903 -8770 25923
rect -8604 25903 -8602 25923
rect -8484 25903 -8482 25923
rect -8436 25903 -8434 25923
rect -8388 25903 -8386 25923
rect -8364 25903 -8362 25923
rect -8340 25903 -8338 25923
rect -8268 25903 -8266 25923
rect -8100 25903 -8098 25923
rect -8052 25903 -8050 25923
rect -7932 25903 -7930 25923
rect -7692 25903 -7690 25923
rect -7620 25903 -7618 25923
rect -7524 25903 -7522 25923
rect -7356 25903 -7354 25923
rect -7308 25903 -7306 25923
rect -7212 25903 -7210 25923
rect -7209 25920 -7195 25923
rect -7188 25920 -7185 25923
rect -7116 25903 -7114 25923
rect -7068 25903 -7066 25923
rect -6972 25903 -6970 25923
rect -6948 25903 -6946 25923
rect -6876 25903 -6874 25923
rect -6852 25903 -6850 25923
rect -6780 25903 -6778 25923
rect -6756 25903 -6754 25923
rect -6660 25903 -6658 25923
rect -6612 25903 -6610 25923
rect -6516 25903 -6514 25923
rect -6492 25903 -6490 25923
rect -6420 25903 -6418 25923
rect -6396 25903 -6394 25923
rect -6372 25903 -6370 25923
rect -6324 25903 -6322 25923
rect -6156 25903 -6154 25923
rect -6060 25903 -6058 25923
rect -6036 25903 -6034 25923
rect -5892 25903 -5890 25923
rect -5652 25903 -5650 25923
rect -5268 25903 -5266 25923
rect -5196 25903 -5194 25923
rect -5172 25903 -5170 25923
rect -5100 25903 -5098 25923
rect -5076 25903 -5074 25923
rect -4980 25903 -4978 25923
rect -4956 25903 -4954 25923
rect -4884 25903 -4882 25923
rect -4860 25903 -4858 25923
rect -4788 25903 -4786 25923
rect -4644 25903 -4642 25923
rect -4548 25903 -4546 25923
rect -4500 25903 -4498 25923
rect -4425 25920 -4411 25923
rect -4404 25923 1949 25927
rect -4404 25920 -4387 25923
rect -4404 25903 -4402 25920
rect -4308 25903 -4306 25923
rect -4260 25903 -4258 25923
rect -4164 25903 -4162 25923
rect -4020 25903 -4018 25923
rect -3876 25903 -3874 25923
rect -3732 25903 -3730 25923
rect -3588 25903 -3586 25923
rect -3564 25903 -3562 25923
rect -3516 25903 -3514 25923
rect -3492 25903 -3490 25923
rect -3468 25903 -3466 25923
rect -3420 25903 -3418 25923
rect -3324 25903 -3322 25923
rect -3252 25903 -3250 25923
rect -3228 25903 -3226 25923
rect -3156 25903 -3154 25923
rect -3132 25903 -3130 25923
rect -3060 25903 -3058 25923
rect -3012 25903 -3010 25923
rect -2964 25903 -2962 25923
rect -2916 25903 -2914 25923
rect -2892 25903 -2890 25923
rect -2868 25903 -2866 25923
rect -2820 25903 -2818 25923
rect -2796 25903 -2794 25923
rect -2772 25903 -2770 25923
rect -2700 25903 -2698 25923
rect -2676 25903 -2674 25923
rect -2604 25903 -2602 25923
rect -2580 25903 -2578 25923
rect -2364 25903 -2362 25923
rect -2268 25903 -2266 25923
rect -2244 25903 -2242 25923
rect -2172 25903 -2170 25923
rect -2148 25903 -2146 25923
rect -2076 25903 -2074 25923
rect -2052 25903 -2050 25923
rect -1980 25903 -1978 25923
rect -1884 25903 -1882 25923
rect -1836 25903 -1834 25923
rect -1596 25903 -1594 25923
rect -1572 25903 -1570 25923
rect -1476 25903 -1474 25923
rect -1380 25903 -1378 25923
rect -1356 25903 -1354 25923
rect -1308 25903 -1306 25923
rect -1260 25903 -1258 25923
rect -1140 25903 -1138 25923
rect -852 25903 -850 25923
rect -756 25903 -754 25923
rect -708 25903 -706 25923
rect -612 25903 -610 25923
rect -588 25903 -586 25923
rect -540 25903 -538 25923
rect -492 25903 -490 25923
rect -444 25903 -442 25923
rect -396 25903 -394 25923
rect -300 25903 -298 25923
rect -276 25903 -274 25923
rect -228 25903 -226 25923
rect -12 25903 -10 25923
rect 156 25903 158 25923
rect 204 25903 206 25923
rect 228 25903 230 25923
rect 252 25903 254 25923
rect 348 25903 350 25923
rect 468 25903 470 25923
rect 492 25903 494 25923
rect 564 25903 566 25923
rect 588 25903 590 25923
rect 636 25903 638 25923
rect 660 25903 662 25923
rect 732 25903 734 25923
rect 756 25903 758 25923
rect 852 25903 854 25923
rect 1020 25903 1022 25923
rect 1092 25903 1094 25923
rect 1116 25903 1118 25923
rect 1212 25903 1214 25923
rect 1308 25903 1310 25923
rect 1332 25903 1334 25923
rect 1380 25903 1382 25923
rect 1428 25903 1430 25923
rect 1476 25903 1478 25923
rect 1524 25903 1526 25923
rect 1548 25903 1550 25923
rect 1620 25903 1622 25923
rect 1644 25903 1646 25923
rect 1692 25903 1694 25923
rect 1716 25903 1718 25923
rect 1740 25903 1742 25923
rect 1788 25903 1790 25923
rect 1935 25920 1949 25923
rect 1959 25923 11093 25927
rect 1959 25920 1973 25923
rect 1980 25920 1983 25923
rect 2028 25903 2030 25923
rect 2076 25903 2078 25923
rect 2100 25903 2102 25923
rect 2124 25903 2126 25923
rect 2172 25903 2174 25923
rect 2196 25903 2198 25923
rect 2220 25903 2222 25923
rect 2268 25903 2270 25923
rect 2292 25903 2294 25923
rect 2316 25903 2318 25923
rect 2364 25903 2366 25923
rect 2412 25903 2414 25923
rect 2460 25903 2462 25923
rect 2508 25903 2510 25923
rect 2580 25903 2582 25923
rect 2604 25903 2606 25923
rect 2676 25903 2678 25923
rect 2700 25903 2702 25923
rect 2748 25903 2750 25923
rect 2772 25903 2774 25923
rect 2796 25903 2798 25923
rect 2844 25903 2846 25923
rect 2868 25903 2870 25923
rect 2892 25903 2894 25923
rect 2940 25903 2942 25923
rect 3012 25903 3014 25923
rect 3108 25903 3110 25923
rect 3156 25903 3158 25923
rect 3252 25903 3254 25923
rect 3348 25903 3350 25923
rect 3396 25903 3398 25923
rect 3468 25903 3470 25923
rect 3492 25903 3494 25923
rect 3564 25903 3566 25923
rect 3612 25903 3614 25923
rect 3636 25903 3638 25923
rect 3660 25903 3662 25923
rect 3708 25903 3710 25923
rect 3732 25903 3734 25923
rect 3804 25903 3806 25923
rect 3828 25903 3830 25923
rect 3924 25903 3926 25923
rect 4020 25903 4022 25923
rect 4044 25903 4046 25923
rect 4092 25903 4094 25923
rect 4116 25903 4118 25923
rect 4140 25903 4142 25923
rect 4188 25903 4190 25923
rect 4212 25903 4214 25923
rect 4236 25903 4238 25923
rect 4308 25903 4310 25923
rect 4332 25903 4334 25923
rect 4404 25903 4406 25923
rect 4500 25903 4502 25923
rect 4596 25903 4598 25923
rect 4860 25903 4862 25923
rect 4956 25903 4958 25923
rect 4980 25903 4982 25923
rect 5004 25903 5006 25923
rect 5076 25903 5078 25923
rect 5100 25903 5102 25923
rect 5124 25903 5126 25923
rect 5172 25903 5174 25923
rect 5220 25903 5222 25923
rect 5268 25903 5270 25923
rect 5388 25903 5390 25923
rect 5484 25903 5486 25923
rect 5508 25903 5510 25923
rect 5532 25903 5534 25923
rect 5628 25903 5630 25923
rect 5652 25903 5654 25923
rect 5748 25903 5750 25923
rect 5796 25903 5798 25923
rect 5844 25903 5846 25923
rect 5892 25903 5894 25923
rect 6132 25903 6134 25923
rect 6180 25903 6182 25923
rect 6228 25903 6230 25923
rect 6252 25903 6254 25923
rect 6276 25903 6278 25923
rect 6324 25903 6326 25923
rect 6372 25903 6374 25923
rect 6492 25903 6494 25923
rect 6588 25903 6590 25923
rect 6612 25903 6614 25923
rect 6660 25903 6662 25923
rect 6684 25903 6686 25923
rect 6708 25903 6710 25923
rect 6780 25903 6782 25923
rect 6804 25903 6806 25923
rect 6828 25903 6830 25923
rect 6900 25903 6902 25923
rect 6924 25903 6926 25923
rect 7020 25903 7022 25923
rect 7140 25903 7142 25923
rect 7236 25903 7238 25923
rect 7332 25903 7334 25923
rect 7380 25903 7382 25923
rect 7428 25903 7430 25923
rect 7452 25903 7454 25923
rect 7476 25903 7478 25923
rect 7524 25903 7526 25923
rect 7548 25903 7550 25923
rect 7572 25903 7574 25923
rect 7620 25903 7622 25923
rect 7644 25903 7646 25923
rect 7668 25903 7670 25923
rect 7740 25903 7742 25923
rect 7788 25903 7790 25923
rect 7884 25903 7886 25923
rect 7956 25903 7958 25923
rect 7980 25903 7982 25923
rect 8028 25903 8030 25923
rect 8196 25903 8198 25923
rect 8244 25903 8246 25923
rect 8268 25903 8270 25923
rect 8292 25903 8294 25923
rect 8340 25903 8342 25923
rect 8364 25903 8366 25923
rect 8388 25903 8390 25923
rect 8436 25903 8438 25923
rect 8460 25903 8462 25923
rect 8556 25903 8558 25923
rect 8604 25903 8606 25923
rect 8652 25903 8654 25923
rect 8700 25903 8702 25923
rect 8724 25903 8726 25923
rect 8748 25903 8750 25923
rect 8820 25903 8822 25923
rect 8844 25903 8846 25923
rect 8868 25903 8870 25923
rect 9516 25903 9518 25923
rect 9612 25903 9614 25923
rect 9660 25903 9662 25923
rect 9684 25903 9686 25923
rect 9708 25903 9710 25923
rect 9756 25903 9758 25923
rect 9780 25903 9782 25923
rect 9804 25903 9806 25923
rect 9852 25903 9854 25923
rect 9876 25903 9878 25923
rect 9900 25903 9902 25923
rect 9948 25903 9950 25923
rect 9972 25903 9974 25923
rect 9996 25903 9998 25923
rect 10068 25903 10070 25923
rect 10092 25903 10094 25923
rect 10116 25903 10118 25923
rect 10164 25903 10166 25923
rect 10188 25903 10190 25923
rect 10212 25903 10214 25923
rect 10284 25903 10286 25923
rect 10308 25903 10310 25923
rect 10332 25903 10334 25923
rect 10380 25903 10382 25923
rect 10404 25903 10406 25923
rect 10428 25903 10430 25923
rect 10476 25903 10478 25923
rect 10500 25903 10502 25923
rect 10524 25903 10526 25923
rect 10572 25903 10574 25923
rect 10596 25903 10598 25923
rect 10620 25903 10622 25923
rect 10668 25903 10670 25923
rect 10692 25903 10694 25923
rect 10716 25903 10718 25923
rect 10788 25903 10790 25923
rect 10836 25903 10838 25923
rect 10956 25903 10958 25923
rect 11004 25903 11006 25923
rect 11052 25903 11054 25923
rect 11076 25903 11078 25923
rect 11079 25920 11093 25923
rect 11100 25923 13493 25927
rect 11100 25920 11117 25923
rect 11124 25920 11127 25923
rect 11100 25903 11102 25920
rect 11172 25903 11174 25923
rect 11220 25903 11222 25923
rect 11340 25903 11342 25923
rect 11436 25903 11438 25923
rect 11532 25903 11534 25923
rect 11580 25903 11582 25923
rect 11628 25903 11630 25923
rect 11676 25903 11678 25923
rect 11724 25903 11726 25923
rect 11772 25903 11774 25923
rect 11796 25903 11798 25923
rect 11892 25903 11894 25923
rect 11988 25903 11990 25923
rect 12060 25903 12062 25923
rect 12132 25903 12134 25923
rect 12228 25903 12230 25923
rect 12276 25903 12278 25923
rect 12324 25903 12326 25923
rect 12420 25903 12422 25923
rect 12444 25903 12446 25923
rect 12492 25903 12494 25923
rect 12516 25903 12518 25923
rect 12540 25903 12542 25923
rect 12588 25903 12590 25923
rect 12636 25903 12638 25923
rect 12732 25903 12734 25923
rect 12756 25903 12758 25923
rect 12804 25903 12806 25923
rect 12828 25903 12830 25923
rect 12852 25903 12854 25923
rect 12900 25903 12902 25923
rect 12948 25903 12950 25923
rect 13044 25903 13046 25923
rect 13068 25903 13070 25923
rect 13116 25903 13118 25923
rect 13284 25903 13286 25923
rect 13332 25903 13334 25923
rect 13479 25920 13493 25923
rect 13503 25923 23933 25927
rect 13503 25920 13517 25923
rect 13524 25920 13527 25923
rect 13572 25903 13574 25923
rect 13644 25903 13646 25923
rect 13668 25903 13670 25923
rect 13764 25903 13766 25923
rect 13812 25903 13814 25923
rect 13860 25903 13862 25923
rect 13908 25903 13910 25923
rect 13956 25903 13958 25923
rect 14004 25903 14006 25923
rect 14100 25903 14102 25923
rect 14196 25903 14198 25923
rect 14292 25903 14294 25923
rect 15132 25903 15134 25923
rect 15180 25903 15182 25923
rect 15228 25903 15230 25923
rect 15252 25903 15254 25923
rect 15324 25903 15326 25923
rect 15396 25903 15398 25923
rect 15420 25903 15422 25923
rect 15492 25903 15494 25923
rect 15540 25903 15542 25923
rect 15636 25903 15638 25923
rect 15660 25903 15662 25923
rect 15708 25903 15710 25923
rect 15732 25903 15734 25923
rect 15756 25903 15758 25923
rect 15804 25903 15806 25923
rect 15828 25903 15830 25923
rect 15852 25903 15854 25923
rect 15900 25903 15902 25923
rect 15948 25903 15950 25923
rect 15996 25903 15998 25923
rect 16044 25903 16046 25923
rect 16164 25903 16166 25923
rect 16260 25903 16262 25923
rect 16308 25903 16310 25923
rect 16332 25903 16334 25923
rect 16356 25903 16358 25923
rect 16404 25903 16406 25923
rect 16452 25903 16454 25923
rect 16548 25903 16550 25923
rect 16572 25903 16574 25923
rect 16620 25903 16622 25923
rect 16668 25903 16670 25923
rect 16716 25903 16718 25923
rect 16764 25903 16766 25923
rect 16812 25903 16814 25923
rect 16884 25903 16886 25923
rect 16908 25903 16910 25923
rect 16980 25903 16982 25923
rect 17052 25903 17054 25923
rect 17196 25903 17198 25923
rect 17220 25903 17222 25923
rect 17292 25903 17294 25923
rect 17316 25903 17318 25923
rect 18084 25903 18086 25923
rect 18132 25903 18134 25923
rect 18396 25903 18398 25923
rect 18492 25903 18494 25923
rect 18516 25903 18518 25923
rect 18564 25903 18566 25923
rect 18612 25903 18614 25923
rect 18660 25903 18662 25923
rect 18708 25903 18710 25923
rect 18756 25903 18758 25923
rect 18804 25903 18806 25923
rect 18852 25903 18854 25923
rect 18900 25903 18902 25923
rect 18996 25903 18998 25923
rect 19020 25903 19022 25923
rect 19092 25903 19094 25923
rect 19116 25903 19118 25923
rect 19140 25903 19142 25923
rect 19188 25903 19190 25923
rect 19236 25903 19238 25923
rect 19332 25903 19334 25923
rect 19476 25903 19478 25923
rect 19788 25903 19790 25923
rect 19836 25903 19838 25923
rect 19860 25903 19862 25923
rect 19884 25903 19886 25923
rect 19932 25903 19934 25923
rect 19956 25903 19958 25923
rect 19980 25903 19982 25923
rect 20028 25903 20030 25923
rect 20052 25903 20054 25923
rect 20076 25903 20078 25923
rect 20148 25903 20150 25923
rect 20172 25903 20174 25923
rect 20196 25903 20198 25923
rect 20268 25903 20270 25923
rect 20292 25903 20294 25923
rect 20388 25903 20390 25923
rect 20412 25903 20414 25923
rect 20508 25903 20510 25923
rect 20556 25903 20558 25923
rect 20604 25903 20606 25923
rect 20916 25903 20918 25923
rect 20964 25903 20966 25923
rect 21012 25903 21014 25923
rect 21060 25903 21062 25923
rect 21084 25903 21086 25923
rect 21108 25903 21110 25923
rect 21204 25903 21206 25923
rect 21300 25903 21302 25923
rect 21324 25903 21326 25923
rect 21444 25903 21446 25923
rect 21468 25903 21470 25923
rect 21564 25903 21566 25923
rect 21612 25903 21614 25923
rect 21684 25903 21686 25923
rect 21708 25903 21710 25923
rect 21828 25903 21830 25923
rect 21924 25903 21926 25923
rect 22068 25903 22070 25923
rect 22188 25903 22190 25923
rect 22212 25903 22214 25923
rect 22884 25903 22886 25923
rect 22980 25903 22982 25923
rect 23076 25903 23078 25923
rect 23100 25903 23102 25923
rect 23124 25903 23126 25923
rect 23244 25903 23246 25923
rect 23340 25903 23342 25923
rect 23412 25903 23414 25923
rect 23508 25903 23510 25923
rect 23556 25903 23558 25923
rect 23652 25903 23654 25923
rect 23676 25903 23678 25923
rect 23724 25903 23726 25923
rect 23772 25903 23774 25923
rect 23820 25903 23822 25923
rect 23916 25903 23918 25923
rect 23919 25920 23933 25923
rect 23943 25923 28451 25927
rect 23943 25920 23957 25923
rect 24012 25903 24014 25923
rect 24084 25903 24086 25923
rect 24396 25903 24398 25923
rect 24492 25903 24494 25923
rect 24516 25903 24518 25923
rect 24588 25903 24590 25923
rect 24612 25903 24614 25923
rect 24684 25903 24686 25923
rect 24732 25903 24734 25923
rect 24756 25903 24758 25923
rect 24780 25903 24782 25923
rect 24852 25903 24854 25923
rect 24876 25903 24878 25923
rect 24972 25903 24974 25923
rect 24996 25903 24998 25923
rect 25068 25903 25070 25923
rect 25164 25903 25166 25923
rect 25260 25903 25262 25923
rect 25308 25903 25310 25923
rect 25356 25903 25358 25923
rect 25380 25903 25382 25923
rect 25404 25903 25406 25923
rect 25500 25903 25502 25923
rect 25596 25903 25598 25923
rect 27036 25903 27038 25923
rect 27108 25903 27110 25923
rect 27324 25903 27326 25923
rect 27396 25903 27398 25923
rect 27420 25903 27422 25923
rect 27540 25903 27542 25923
rect 27564 25903 27566 25923
rect 28311 25920 28325 25923
rect 27697 25903 27731 25904
rect -16943 25899 -16435 25903
rect -16836 25896 -16834 25899
rect -16836 25880 -16833 25896
rect -16847 25879 -16813 25880
rect -16740 25879 -16738 25899
rect -16692 25879 -16690 25899
rect -16524 25879 -16522 25899
rect -16449 25896 -16435 25899
rect -16425 25899 27731 25903
rect -16425 25896 -16411 25899
rect -16404 25879 -16401 25899
rect -16380 25896 -16378 25899
rect -16380 25879 -16377 25896
rect -16356 25879 -16354 25899
rect -16284 25879 -16282 25899
rect -16260 25879 -16258 25899
rect -15324 25879 -15322 25899
rect -14772 25879 -14770 25899
rect -14508 25879 -14506 25899
rect -14436 25879 -14434 25899
rect -14340 25879 -14338 25899
rect -13980 25879 -13978 25899
rect -13932 25879 -13930 25899
rect -13884 25879 -13882 25899
rect -13788 25879 -13786 25899
rect -13572 25879 -13570 25899
rect -13356 25879 -13354 25899
rect -13284 25879 -13282 25899
rect -13068 25879 -13066 25899
rect -12828 25880 -12826 25899
rect -12863 25879 -12805 25880
rect -12780 25879 -12778 25899
rect -12660 25879 -12658 25899
rect -12564 25879 -12562 25899
rect -12492 25879 -12490 25899
rect -12396 25879 -12394 25899
rect -12348 25879 -12346 25899
rect -12252 25879 -12250 25899
rect -12156 25879 -12154 25899
rect -12060 25879 -12058 25899
rect -11844 25879 -11842 25899
rect -11796 25879 -11794 25899
rect -11676 25879 -11674 25899
rect -11580 25879 -11578 25899
rect -11556 25879 -11554 25899
rect -11508 25879 -11506 25899
rect -11460 25879 -11458 25899
rect -11436 25879 -11434 25899
rect -11412 25879 -11410 25899
rect -11364 25879 -11362 25899
rect -11340 25879 -11338 25899
rect -11196 25879 -11194 25899
rect -11124 25879 -11122 25899
rect -11100 25879 -11098 25899
rect -11028 25879 -11026 25899
rect -10740 25879 -10738 25899
rect -10668 25879 -10666 25899
rect -10644 25879 -10642 25899
rect -9996 25879 -9994 25899
rect -9828 25879 -9826 25899
rect -9732 25879 -9730 25899
rect -9612 25879 -9610 25899
rect -9516 25879 -9514 25899
rect -9468 25879 -9466 25899
rect -9420 25879 -9418 25899
rect -9396 25879 -9394 25899
rect -9300 25879 -9298 25899
rect -9252 25879 -9250 25899
rect -9084 25880 -9082 25899
rect -9119 25879 -9061 25880
rect -8988 25879 -8986 25899
rect -8892 25879 -8890 25899
rect -8772 25879 -8770 25899
rect -8604 25879 -8602 25899
rect -8484 25879 -8482 25899
rect -8436 25879 -8434 25899
rect -8388 25879 -8386 25899
rect -8364 25879 -8362 25899
rect -8340 25879 -8338 25899
rect -8268 25879 -8266 25899
rect -8100 25879 -8098 25899
rect -8052 25879 -8050 25899
rect -7932 25879 -7930 25899
rect -7692 25879 -7690 25899
rect -7620 25879 -7618 25899
rect -7524 25879 -7522 25899
rect -7356 25879 -7354 25899
rect -7308 25879 -7306 25899
rect -7212 25879 -7210 25899
rect -7116 25879 -7114 25899
rect -7068 25879 -7066 25899
rect -6972 25879 -6970 25899
rect -6948 25879 -6946 25899
rect -6876 25879 -6874 25899
rect -6852 25879 -6850 25899
rect -6780 25879 -6778 25899
rect -6756 25879 -6754 25899
rect -6660 25879 -6658 25899
rect -6612 25879 -6610 25899
rect -6516 25879 -6514 25899
rect -6492 25879 -6490 25899
rect -6420 25879 -6418 25899
rect -6396 25879 -6394 25899
rect -6372 25879 -6370 25899
rect -6324 25879 -6322 25899
rect -6156 25879 -6154 25899
rect -6060 25879 -6058 25899
rect -6036 25879 -6034 25899
rect -5892 25879 -5890 25899
rect -5652 25879 -5650 25899
rect -5268 25879 -5266 25899
rect -5196 25879 -5194 25899
rect -5172 25879 -5170 25899
rect -5100 25879 -5098 25899
rect -5076 25879 -5074 25899
rect -4980 25879 -4978 25899
rect -4956 25879 -4954 25899
rect -4884 25879 -4882 25899
rect -4860 25879 -4858 25899
rect -4788 25879 -4786 25899
rect -4644 25879 -4642 25899
rect -4548 25879 -4546 25899
rect -4500 25879 -4498 25899
rect -4404 25879 -4402 25899
rect -4308 25879 -4306 25899
rect -4260 25879 -4258 25899
rect -4164 25879 -4162 25899
rect -4020 25879 -4018 25899
rect -3876 25879 -3874 25899
rect -3732 25879 -3730 25899
rect -3588 25879 -3586 25899
rect -3564 25879 -3562 25899
rect -3516 25879 -3514 25899
rect -3492 25879 -3490 25899
rect -3468 25879 -3466 25899
rect -3420 25879 -3418 25899
rect -3359 25879 -3325 25880
rect -3324 25879 -3322 25899
rect -3252 25879 -3250 25899
rect -3228 25879 -3226 25899
rect -3156 25879 -3154 25899
rect -3132 25879 -3130 25899
rect -3060 25879 -3058 25899
rect -3012 25879 -3010 25899
rect -2964 25879 -2962 25899
rect -2916 25879 -2914 25899
rect -2892 25879 -2890 25899
rect -2868 25879 -2866 25899
rect -2820 25879 -2818 25899
rect -2796 25879 -2794 25899
rect -2772 25879 -2770 25899
rect -2700 25879 -2698 25899
rect -2676 25879 -2674 25899
rect -2604 25879 -2602 25899
rect -2580 25879 -2578 25899
rect -2364 25879 -2362 25899
rect -2268 25879 -2266 25899
rect -2244 25879 -2242 25899
rect -2172 25879 -2170 25899
rect -2148 25879 -2146 25899
rect -2076 25879 -2074 25899
rect -2052 25879 -2050 25899
rect -1980 25879 -1978 25899
rect -1884 25879 -1882 25899
rect -1836 25879 -1834 25899
rect -1596 25879 -1594 25899
rect -1572 25879 -1570 25899
rect -1476 25879 -1474 25899
rect -1380 25879 -1378 25899
rect -1356 25879 -1354 25899
rect -1308 25879 -1306 25899
rect -1260 25879 -1258 25899
rect -1140 25879 -1138 25899
rect -852 25879 -850 25899
rect -756 25879 -754 25899
rect -708 25879 -706 25899
rect -612 25879 -610 25899
rect -588 25879 -586 25899
rect -540 25879 -538 25899
rect -492 25879 -490 25899
rect -444 25879 -442 25899
rect -396 25879 -394 25899
rect -300 25879 -298 25899
rect -276 25879 -274 25899
rect -228 25879 -226 25899
rect -12 25879 -10 25899
rect 156 25879 158 25899
rect 204 25879 206 25899
rect 228 25879 230 25899
rect 252 25879 254 25899
rect 348 25879 350 25899
rect 468 25879 470 25899
rect 492 25879 494 25899
rect 564 25879 566 25899
rect 588 25879 590 25899
rect 636 25879 638 25899
rect 660 25879 662 25899
rect 732 25879 734 25899
rect 756 25879 758 25899
rect 852 25879 854 25899
rect 1020 25879 1022 25899
rect 1092 25879 1094 25899
rect 1116 25879 1118 25899
rect 1212 25879 1214 25899
rect 1308 25879 1310 25899
rect 1332 25879 1334 25899
rect 1380 25879 1382 25899
rect 1428 25879 1430 25899
rect 1476 25879 1478 25899
rect 1524 25879 1526 25899
rect 1548 25879 1550 25899
rect 1620 25879 1622 25899
rect 1644 25879 1646 25899
rect 1692 25879 1694 25899
rect 1716 25879 1718 25899
rect 1740 25879 1742 25899
rect 1788 25879 1790 25899
rect 2028 25879 2030 25899
rect 2076 25879 2078 25899
rect 2100 25879 2102 25899
rect 2124 25879 2126 25899
rect 2172 25879 2174 25899
rect 2196 25879 2198 25899
rect 2220 25879 2222 25899
rect 2268 25879 2270 25899
rect 2292 25879 2294 25899
rect 2316 25879 2318 25899
rect 2364 25879 2366 25899
rect 2412 25879 2414 25899
rect 2460 25879 2462 25899
rect 2508 25879 2510 25899
rect 2580 25879 2582 25899
rect 2604 25879 2606 25899
rect 2676 25879 2678 25899
rect 2700 25879 2702 25899
rect 2748 25879 2750 25899
rect 2772 25879 2774 25899
rect 2796 25879 2798 25899
rect 2844 25879 2846 25899
rect 2868 25879 2870 25899
rect 2892 25879 2894 25899
rect 2940 25879 2942 25899
rect 3012 25879 3014 25899
rect 3108 25879 3110 25899
rect 3156 25879 3158 25899
rect 3252 25879 3254 25899
rect 3348 25879 3350 25899
rect 3396 25879 3398 25899
rect 3468 25879 3470 25899
rect 3492 25879 3494 25899
rect 3564 25879 3566 25899
rect 3612 25879 3614 25899
rect 3636 25879 3638 25899
rect 3660 25879 3662 25899
rect 3708 25879 3710 25899
rect 3732 25879 3734 25899
rect 3804 25879 3806 25899
rect 3828 25879 3830 25899
rect 3924 25879 3926 25899
rect 4020 25879 4022 25899
rect 4044 25879 4046 25899
rect 4092 25879 4094 25899
rect 4116 25879 4118 25899
rect 4140 25879 4142 25899
rect 4188 25879 4190 25899
rect 4212 25879 4214 25899
rect 4236 25879 4238 25899
rect 4308 25879 4310 25899
rect 4332 25879 4334 25899
rect 4404 25879 4406 25899
rect 4500 25879 4502 25899
rect 4596 25879 4598 25899
rect 4860 25879 4862 25899
rect 4956 25879 4958 25899
rect 4980 25879 4982 25899
rect 5004 25879 5006 25899
rect 5076 25879 5078 25899
rect 5100 25879 5102 25899
rect 5124 25879 5126 25899
rect 5172 25879 5174 25899
rect 5220 25879 5222 25899
rect 5268 25879 5270 25899
rect 5388 25879 5390 25899
rect 5484 25879 5486 25899
rect 5508 25879 5510 25899
rect 5532 25879 5534 25899
rect 5628 25879 5630 25899
rect 5652 25879 5654 25899
rect 5748 25879 5750 25899
rect 5796 25879 5798 25899
rect 5844 25879 5846 25899
rect 5892 25879 5894 25899
rect 6132 25879 6134 25899
rect 6180 25879 6182 25899
rect 6228 25879 6230 25899
rect 6252 25879 6254 25899
rect 6276 25879 6278 25899
rect 6324 25879 6326 25899
rect 6372 25879 6374 25899
rect 6492 25879 6494 25899
rect 6588 25879 6590 25899
rect 6612 25879 6614 25899
rect 6660 25879 6662 25899
rect 6684 25879 6686 25899
rect 6708 25879 6710 25899
rect 6780 25879 6782 25899
rect 6804 25879 6806 25899
rect 6828 25879 6830 25899
rect 6900 25879 6902 25899
rect 6924 25879 6926 25899
rect 7020 25879 7022 25899
rect 7140 25879 7142 25899
rect 7236 25879 7238 25899
rect 7332 25879 7334 25899
rect 7380 25879 7382 25899
rect 7428 25879 7430 25899
rect 7452 25879 7454 25899
rect 7476 25879 7478 25899
rect 7524 25879 7526 25899
rect 7548 25879 7550 25899
rect 7572 25879 7574 25899
rect 7620 25879 7622 25899
rect 7644 25879 7646 25899
rect 7668 25879 7670 25899
rect 7740 25879 7742 25899
rect 7788 25879 7790 25899
rect 7884 25879 7886 25899
rect 7956 25879 7958 25899
rect 7980 25879 7982 25899
rect 8028 25879 8030 25899
rect 8196 25879 8198 25899
rect 8244 25879 8246 25899
rect 8268 25879 8270 25899
rect 8292 25879 8294 25899
rect 8340 25879 8342 25899
rect 8364 25879 8366 25899
rect 8388 25879 8390 25899
rect 8436 25879 8438 25899
rect 8460 25879 8462 25899
rect 8556 25879 8558 25899
rect 8604 25879 8606 25899
rect 8652 25879 8654 25899
rect 8700 25879 8702 25899
rect 8724 25879 8726 25899
rect 8748 25879 8750 25899
rect 8820 25879 8822 25899
rect 8844 25879 8846 25899
rect 8868 25879 8870 25899
rect 9516 25879 9518 25899
rect 9612 25879 9614 25899
rect 9660 25879 9662 25899
rect 9684 25879 9686 25899
rect 9708 25879 9710 25899
rect 9756 25879 9758 25899
rect 9780 25879 9782 25899
rect 9804 25879 9806 25899
rect 9852 25879 9854 25899
rect 9876 25879 9878 25899
rect 9900 25879 9902 25899
rect 9948 25879 9950 25899
rect 9972 25879 9974 25899
rect 9996 25879 9998 25899
rect 10068 25879 10070 25899
rect 10092 25879 10094 25899
rect 10116 25879 10118 25899
rect 10164 25879 10166 25899
rect 10188 25879 10190 25899
rect 10212 25879 10214 25899
rect 10284 25879 10286 25899
rect 10308 25879 10310 25899
rect 10332 25879 10334 25899
rect 10380 25879 10382 25899
rect 10404 25879 10406 25899
rect 10428 25879 10430 25899
rect 10476 25879 10478 25899
rect 10500 25879 10502 25899
rect 10524 25879 10526 25899
rect 10572 25879 10574 25899
rect 10596 25879 10598 25899
rect 10620 25879 10622 25899
rect 10668 25879 10670 25899
rect 10692 25879 10694 25899
rect 10716 25879 10718 25899
rect 10788 25879 10790 25899
rect 10836 25879 10838 25899
rect 10956 25879 10958 25899
rect 11004 25879 11006 25899
rect 11052 25879 11054 25899
rect 11076 25879 11078 25899
rect 11100 25879 11102 25899
rect 11172 25879 11174 25899
rect 11220 25879 11222 25899
rect 11340 25879 11342 25899
rect 11436 25879 11438 25899
rect 11532 25879 11534 25899
rect 11580 25879 11582 25899
rect 11628 25879 11630 25899
rect 11676 25879 11678 25899
rect 11724 25879 11726 25899
rect 11772 25879 11774 25899
rect 11796 25879 11798 25899
rect 11892 25879 11894 25899
rect 11988 25879 11990 25899
rect 12060 25879 12062 25899
rect 12132 25879 12134 25899
rect 12228 25879 12230 25899
rect 12276 25879 12278 25899
rect 12324 25879 12326 25899
rect 12420 25879 12422 25899
rect 12444 25879 12446 25899
rect 12492 25879 12494 25899
rect 12516 25879 12518 25899
rect 12540 25879 12542 25899
rect 12588 25879 12590 25899
rect 12636 25879 12638 25899
rect 12732 25879 12734 25899
rect 12756 25879 12758 25899
rect 12804 25879 12806 25899
rect 12828 25879 12830 25899
rect 12852 25879 12854 25899
rect 12900 25879 12902 25899
rect 12948 25879 12950 25899
rect 13044 25879 13046 25899
rect 13068 25879 13070 25899
rect 13116 25879 13118 25899
rect 13284 25879 13286 25899
rect 13332 25879 13334 25899
rect 13572 25879 13574 25899
rect 13644 25879 13646 25899
rect 13668 25879 13670 25899
rect 13764 25879 13766 25899
rect 13812 25879 13814 25899
rect 13860 25879 13862 25899
rect 13908 25879 13910 25899
rect 13956 25879 13958 25899
rect 14004 25879 14006 25899
rect 14100 25879 14102 25899
rect 14196 25879 14198 25899
rect 14292 25879 14294 25899
rect 15132 25879 15134 25899
rect 15180 25879 15182 25899
rect 15228 25879 15230 25899
rect 15252 25879 15254 25899
rect 15324 25879 15326 25899
rect 15396 25879 15398 25899
rect 15420 25879 15422 25899
rect 15492 25879 15494 25899
rect 15540 25879 15542 25899
rect 15636 25879 15638 25899
rect 15660 25879 15662 25899
rect 15708 25879 15710 25899
rect 15732 25879 15734 25899
rect 15756 25879 15758 25899
rect 15804 25879 15806 25899
rect 15828 25879 15830 25899
rect 15852 25879 15854 25899
rect 15900 25879 15902 25899
rect 15948 25879 15950 25899
rect 15996 25879 15998 25899
rect 16044 25879 16046 25899
rect 16164 25879 16166 25899
rect 16260 25879 16262 25899
rect 16308 25879 16310 25899
rect 16332 25879 16334 25899
rect 16356 25879 16358 25899
rect 16404 25879 16406 25899
rect 16452 25879 16454 25899
rect 16548 25879 16550 25899
rect 16572 25879 16574 25899
rect 16620 25879 16622 25899
rect 16668 25879 16670 25899
rect 16716 25879 16718 25899
rect 16764 25879 16766 25899
rect 16812 25879 16814 25899
rect 16884 25879 16886 25899
rect 16908 25879 16910 25899
rect 16980 25879 16982 25899
rect 17052 25879 17054 25899
rect 17196 25879 17198 25899
rect 17220 25879 17222 25899
rect 17292 25879 17294 25899
rect 17316 25879 17318 25899
rect 18084 25879 18086 25899
rect 18132 25879 18134 25899
rect 18217 25879 18275 25880
rect 18396 25879 18398 25899
rect 18492 25879 18494 25899
rect 18516 25879 18518 25899
rect 18564 25879 18566 25899
rect 18612 25879 18614 25899
rect 18660 25879 18662 25899
rect 18708 25879 18710 25899
rect 18756 25879 18758 25899
rect 18804 25879 18806 25899
rect 18852 25879 18854 25899
rect 18900 25879 18902 25899
rect 18996 25879 18998 25899
rect 19020 25879 19022 25899
rect 19092 25879 19094 25899
rect 19116 25879 19118 25899
rect 19140 25879 19142 25899
rect 19188 25879 19190 25899
rect 19236 25879 19238 25899
rect 19332 25879 19334 25899
rect 19476 25879 19478 25899
rect 19788 25879 19790 25899
rect 19836 25879 19838 25899
rect 19860 25879 19862 25899
rect 19884 25879 19886 25899
rect 19932 25879 19934 25899
rect 19956 25879 19958 25899
rect 19980 25879 19982 25899
rect 20028 25879 20030 25899
rect 20052 25879 20054 25899
rect 20076 25879 20078 25899
rect 20148 25879 20150 25899
rect 20172 25879 20174 25899
rect 20196 25879 20198 25899
rect 20268 25879 20270 25899
rect 20292 25879 20294 25899
rect 20388 25879 20390 25899
rect 20412 25879 20414 25899
rect 20508 25879 20510 25899
rect 20556 25879 20558 25899
rect 20604 25879 20606 25899
rect 20916 25879 20918 25899
rect 20964 25879 20966 25899
rect 21012 25879 21014 25899
rect 21060 25879 21062 25899
rect 21084 25879 21086 25899
rect 21108 25879 21110 25899
rect 21204 25879 21206 25899
rect 21300 25879 21302 25899
rect 21324 25879 21326 25899
rect 21444 25879 21446 25899
rect 21468 25879 21470 25899
rect 21564 25879 21566 25899
rect 21612 25879 21614 25899
rect 21684 25879 21686 25899
rect 21708 25879 21710 25899
rect 21828 25879 21830 25899
rect 21924 25879 21926 25899
rect 22068 25879 22070 25899
rect 22188 25879 22190 25899
rect 22212 25879 22214 25899
rect 22884 25879 22886 25899
rect 22980 25879 22982 25899
rect 23076 25879 23078 25899
rect 23100 25879 23102 25899
rect 23124 25879 23126 25899
rect 23244 25879 23246 25899
rect 23340 25879 23342 25899
rect 23412 25879 23414 25899
rect 23508 25879 23510 25899
rect 23556 25879 23558 25899
rect 23652 25879 23654 25899
rect 23676 25879 23678 25899
rect 23724 25879 23726 25899
rect 23772 25879 23774 25899
rect 23820 25879 23822 25899
rect 23916 25879 23918 25899
rect 24012 25879 24014 25899
rect 24084 25879 24086 25899
rect 24396 25879 24398 25899
rect 24492 25879 24494 25899
rect 24516 25879 24518 25899
rect 24588 25879 24590 25899
rect 24612 25879 24614 25899
rect 24684 25879 24686 25899
rect 24732 25879 24734 25899
rect 24756 25879 24758 25899
rect 24780 25879 24782 25899
rect 24852 25879 24854 25899
rect 24876 25879 24878 25899
rect 24972 25879 24974 25899
rect 24996 25879 24998 25899
rect 25068 25879 25070 25899
rect 25164 25879 25166 25899
rect 25177 25879 25235 25880
rect 25260 25879 25262 25899
rect 25308 25879 25310 25899
rect 25356 25879 25358 25899
rect 25380 25879 25382 25899
rect 25404 25879 25406 25899
rect 25500 25879 25502 25899
rect 25596 25879 25598 25899
rect 27036 25879 27038 25899
rect 27108 25879 27110 25899
rect 27324 25879 27326 25899
rect 27396 25879 27398 25899
rect 27420 25879 27422 25899
rect 27540 25879 27542 25899
rect 27564 25880 27566 25899
rect 27553 25879 27587 25880
rect -16847 25875 -16411 25879
rect -16847 25872 -16843 25875
rect -16836 25872 -16833 25875
rect -16740 25872 -16738 25875
rect -16740 25855 -16737 25872
rect -16692 25855 -16690 25875
rect -16524 25855 -16522 25875
rect -16425 25872 -16411 25875
rect -16404 25875 27587 25879
rect -16404 25872 -16387 25875
rect -16380 25872 -16377 25875
rect -16404 25855 -16402 25872
rect -16356 25855 -16354 25875
rect -16284 25855 -16282 25875
rect -16260 25855 -16258 25875
rect -15324 25855 -15322 25875
rect -14772 25855 -14770 25875
rect -14615 25855 -14581 25856
rect -14508 25855 -14506 25875
rect -14436 25855 -14434 25875
rect -14340 25855 -14338 25875
rect -13980 25855 -13978 25875
rect -13932 25855 -13930 25875
rect -13884 25855 -13882 25875
rect -13788 25855 -13786 25875
rect -13572 25855 -13570 25875
rect -13356 25855 -13354 25875
rect -13284 25855 -13282 25875
rect -13068 25855 -13066 25875
rect -12839 25870 -12836 25875
rect -12828 25870 -12826 25875
rect -12829 25856 -12826 25870
rect -12780 25855 -12778 25875
rect -12756 25855 -12753 25872
rect -12660 25855 -12658 25875
rect -12564 25855 -12562 25875
rect -12492 25855 -12490 25875
rect -12396 25855 -12394 25875
rect -12348 25855 -12346 25875
rect -12252 25855 -12250 25875
rect -12156 25855 -12154 25875
rect -12060 25855 -12058 25875
rect -11844 25855 -11842 25875
rect -11796 25855 -11794 25875
rect -11676 25855 -11674 25875
rect -11580 25856 -11578 25875
rect -11591 25855 -11557 25856
rect -11556 25855 -11554 25875
rect -11508 25855 -11506 25875
rect -11460 25856 -11458 25875
rect -11471 25855 -11437 25856
rect -11436 25855 -11434 25875
rect -11412 25855 -11410 25875
rect -11364 25855 -11362 25875
rect -11340 25855 -11338 25875
rect -11196 25855 -11194 25875
rect -11124 25855 -11122 25875
rect -11100 25855 -11098 25875
rect -11028 25855 -11026 25875
rect -10740 25855 -10738 25875
rect -10668 25855 -10666 25875
rect -10644 25855 -10642 25875
rect -9996 25855 -9994 25875
rect -9828 25855 -9826 25875
rect -9732 25855 -9730 25875
rect -9612 25855 -9610 25875
rect -9516 25855 -9514 25875
rect -9468 25855 -9466 25875
rect -9420 25855 -9418 25875
rect -9396 25856 -9394 25875
rect -9407 25855 -9373 25856
rect -9300 25855 -9298 25875
rect -9252 25855 -9250 25875
rect -9095 25870 -9092 25875
rect -9084 25870 -9082 25875
rect -9085 25856 -9082 25870
rect -8988 25872 -8986 25875
rect -8988 25855 -8985 25872
rect -8892 25856 -8890 25875
rect -8903 25855 -8869 25856
rect -8772 25855 -8770 25875
rect -8604 25855 -8602 25875
rect -8484 25855 -8482 25875
rect -8436 25855 -8434 25875
rect -8388 25855 -8386 25875
rect -8364 25855 -8362 25875
rect -8340 25855 -8338 25875
rect -8268 25855 -8266 25875
rect -8100 25855 -8098 25875
rect -8052 25855 -8050 25875
rect -7932 25855 -7930 25875
rect -7692 25855 -7690 25875
rect -7620 25855 -7618 25875
rect -7524 25855 -7522 25875
rect -7356 25855 -7354 25875
rect -7308 25855 -7306 25875
rect -7212 25855 -7210 25875
rect -7116 25855 -7114 25875
rect -7068 25855 -7066 25875
rect -6972 25855 -6970 25875
rect -6948 25855 -6946 25875
rect -6876 25855 -6874 25875
rect -6852 25855 -6850 25875
rect -6780 25855 -6778 25875
rect -6756 25855 -6754 25875
rect -6660 25855 -6658 25875
rect -6612 25855 -6610 25875
rect -6516 25855 -6514 25875
rect -6492 25855 -6490 25875
rect -6420 25855 -6418 25875
rect -6396 25855 -6394 25875
rect -6372 25855 -6370 25875
rect -6324 25855 -6322 25875
rect -6156 25855 -6154 25875
rect -6060 25855 -6058 25875
rect -6036 25855 -6034 25875
rect -5892 25855 -5890 25875
rect -5652 25855 -5650 25875
rect -5268 25855 -5266 25875
rect -5196 25855 -5194 25875
rect -5172 25855 -5170 25875
rect -5100 25855 -5098 25875
rect -5076 25855 -5074 25875
rect -4980 25855 -4978 25875
rect -4956 25855 -4954 25875
rect -4884 25855 -4882 25875
rect -4860 25855 -4858 25875
rect -4788 25855 -4786 25875
rect -4644 25855 -4642 25875
rect -4548 25855 -4546 25875
rect -4500 25855 -4498 25875
rect -4404 25855 -4402 25875
rect -4308 25855 -4306 25875
rect -4260 25855 -4258 25875
rect -4164 25855 -4162 25875
rect -4020 25855 -4018 25875
rect -3876 25855 -3874 25875
rect -3732 25855 -3730 25875
rect -3588 25855 -3586 25875
rect -3564 25855 -3562 25875
rect -3516 25855 -3514 25875
rect -3492 25855 -3490 25875
rect -3468 25855 -3466 25875
rect -3420 25855 -3418 25875
rect -3324 25855 -3322 25875
rect -3252 25872 -3250 25875
rect -3252 25855 -3249 25872
rect -3228 25855 -3226 25875
rect -3156 25855 -3154 25875
rect -3132 25855 -3130 25875
rect -3060 25855 -3058 25875
rect -3012 25855 -3010 25875
rect -2964 25855 -2962 25875
rect -2916 25855 -2914 25875
rect -2892 25855 -2890 25875
rect -2868 25855 -2866 25875
rect -2820 25855 -2818 25875
rect -2796 25855 -2794 25875
rect -2772 25855 -2770 25875
rect -2700 25856 -2698 25875
rect -2711 25855 -2677 25856
rect -2676 25855 -2674 25875
rect -2604 25855 -2602 25875
rect -2580 25855 -2578 25875
rect -2364 25855 -2362 25875
rect -2268 25855 -2266 25875
rect -2244 25855 -2242 25875
rect -2172 25855 -2170 25875
rect -2148 25855 -2146 25875
rect -2076 25855 -2074 25875
rect -2052 25855 -2050 25875
rect -1980 25855 -1978 25875
rect -1884 25855 -1882 25875
rect -1836 25855 -1834 25875
rect -1596 25856 -1594 25875
rect -1607 25855 -1573 25856
rect -1572 25855 -1570 25875
rect -1476 25855 -1474 25875
rect -1380 25855 -1378 25875
rect -1356 25855 -1354 25875
rect -1308 25855 -1306 25875
rect -1260 25855 -1258 25875
rect -1140 25855 -1138 25875
rect -852 25855 -850 25875
rect -756 25855 -754 25875
rect -708 25855 -706 25875
rect -612 25855 -610 25875
rect -588 25855 -586 25875
rect -540 25855 -538 25875
rect -492 25855 -490 25875
rect -444 25855 -442 25875
rect -396 25855 -394 25875
rect -300 25855 -298 25875
rect -276 25855 -274 25875
rect -228 25855 -226 25875
rect -12 25855 -10 25875
rect 156 25855 158 25875
rect 204 25855 206 25875
rect 228 25856 230 25875
rect 217 25855 251 25856
rect 252 25855 254 25875
rect 348 25855 350 25875
rect 468 25855 470 25875
rect 492 25855 494 25875
rect 564 25855 566 25875
rect 588 25855 590 25875
rect 636 25855 638 25875
rect 660 25855 662 25875
rect 732 25855 734 25875
rect 756 25856 758 25875
rect 745 25855 779 25856
rect 852 25855 854 25875
rect 1020 25855 1022 25875
rect 1092 25855 1094 25875
rect 1116 25855 1118 25875
rect 1212 25855 1214 25875
rect 1308 25855 1310 25875
rect 1332 25855 1334 25875
rect 1380 25855 1382 25875
rect 1428 25855 1430 25875
rect 1476 25855 1478 25875
rect 1524 25856 1526 25875
rect 1513 25855 1547 25856
rect 1548 25855 1550 25875
rect 1620 25856 1622 25875
rect 1609 25855 1643 25856
rect 1644 25855 1646 25875
rect 1692 25855 1694 25875
rect 1716 25855 1718 25875
rect 1740 25855 1742 25875
rect 1788 25855 1790 25875
rect 2028 25855 2030 25875
rect 2076 25855 2078 25875
rect 2100 25855 2102 25875
rect 2124 25855 2126 25875
rect 2172 25855 2174 25875
rect 2196 25855 2198 25875
rect 2220 25855 2222 25875
rect 2268 25855 2270 25875
rect 2292 25856 2294 25875
rect 2281 25855 2315 25856
rect 2316 25855 2318 25875
rect 2364 25855 2366 25875
rect 2412 25855 2414 25875
rect 2460 25855 2462 25875
rect 2508 25855 2510 25875
rect 2580 25855 2582 25875
rect 2604 25855 2606 25875
rect 2676 25855 2678 25875
rect 2700 25855 2702 25875
rect 2748 25855 2750 25875
rect 2772 25855 2774 25875
rect 2796 25855 2798 25875
rect 2844 25855 2846 25875
rect 2868 25855 2870 25875
rect 2892 25855 2894 25875
rect 2940 25855 2942 25875
rect 3012 25855 3014 25875
rect 3108 25855 3110 25875
rect 3121 25855 3155 25856
rect 3156 25855 3158 25875
rect 3252 25855 3254 25875
rect 3348 25855 3350 25875
rect 3361 25855 3395 25856
rect 3396 25855 3398 25875
rect 3468 25855 3470 25875
rect 3492 25856 3494 25875
rect 3481 25855 3515 25856
rect 3564 25855 3566 25875
rect 3612 25855 3614 25875
rect 3636 25855 3638 25875
rect 3660 25855 3662 25875
rect 3708 25855 3710 25875
rect 3732 25855 3734 25875
rect 3804 25855 3806 25875
rect 3828 25855 3830 25875
rect 3924 25855 3926 25875
rect 4020 25855 4022 25875
rect 4044 25855 4046 25875
rect 4092 25855 4094 25875
rect 4116 25855 4118 25875
rect 4140 25855 4142 25875
rect 4188 25855 4190 25875
rect 4212 25855 4214 25875
rect 4236 25855 4238 25875
rect 4308 25855 4310 25875
rect 4332 25855 4334 25875
rect 4404 25855 4406 25875
rect 4500 25855 4502 25875
rect 4596 25855 4598 25875
rect 4681 25855 4739 25856
rect 4860 25855 4862 25875
rect 4956 25855 4958 25875
rect 4980 25855 4982 25875
rect 5004 25855 5006 25875
rect 5076 25855 5078 25875
rect 5100 25855 5102 25875
rect 5124 25855 5126 25875
rect 5172 25855 5174 25875
rect 5220 25855 5222 25875
rect 5268 25855 5270 25875
rect 5388 25855 5390 25875
rect 5484 25855 5486 25875
rect 5508 25855 5510 25875
rect 5532 25855 5534 25875
rect 5628 25855 5630 25875
rect 5652 25855 5654 25875
rect 5748 25855 5750 25875
rect 5796 25855 5798 25875
rect 5844 25855 5846 25875
rect 5892 25855 5894 25875
rect 6132 25855 6134 25875
rect 6180 25855 6182 25875
rect 6228 25855 6230 25875
rect 6252 25855 6254 25875
rect 6276 25855 6278 25875
rect 6324 25855 6326 25875
rect 6372 25855 6374 25875
rect 6492 25855 6494 25875
rect 6588 25855 6590 25875
rect 6612 25855 6614 25875
rect 6660 25855 6662 25875
rect 6684 25855 6686 25875
rect 6708 25855 6710 25875
rect 6780 25855 6782 25875
rect 6804 25855 6806 25875
rect 6828 25855 6830 25875
rect 6900 25855 6902 25875
rect 6924 25855 6926 25875
rect 7020 25855 7022 25875
rect 7140 25855 7142 25875
rect 7236 25855 7238 25875
rect 7332 25855 7334 25875
rect 7380 25855 7382 25875
rect 7428 25855 7430 25875
rect 7452 25855 7454 25875
rect 7476 25855 7478 25875
rect 7524 25855 7526 25875
rect 7548 25855 7550 25875
rect 7572 25855 7574 25875
rect 7620 25855 7622 25875
rect 7644 25855 7646 25875
rect 7668 25855 7670 25875
rect 7740 25855 7742 25875
rect 7788 25855 7790 25875
rect 7884 25855 7886 25875
rect 7956 25855 7958 25875
rect 7980 25855 7982 25875
rect 8028 25855 8030 25875
rect 8196 25855 8198 25875
rect 8244 25855 8246 25875
rect 8268 25855 8270 25875
rect 8292 25855 8294 25875
rect 8340 25855 8342 25875
rect 8364 25855 8366 25875
rect 8388 25855 8390 25875
rect 8436 25855 8438 25875
rect 8460 25855 8462 25875
rect 8556 25855 8558 25875
rect 8604 25855 8606 25875
rect 8652 25855 8654 25875
rect 8700 25855 8702 25875
rect 8724 25855 8726 25875
rect 8748 25855 8750 25875
rect 8820 25855 8822 25875
rect 8844 25855 8846 25875
rect 8868 25855 8870 25875
rect 9516 25855 9518 25875
rect 9612 25855 9614 25875
rect 9660 25855 9662 25875
rect 9684 25855 9686 25875
rect 9708 25855 9710 25875
rect 9756 25855 9758 25875
rect 9780 25855 9782 25875
rect 9804 25855 9806 25875
rect 9852 25855 9854 25875
rect 9876 25855 9878 25875
rect 9900 25855 9902 25875
rect 9948 25855 9950 25875
rect 9972 25855 9974 25875
rect 9996 25855 9998 25875
rect 10068 25855 10070 25875
rect 10092 25855 10094 25875
rect 10116 25855 10118 25875
rect 10164 25855 10166 25875
rect 10188 25855 10190 25875
rect 10212 25855 10214 25875
rect 10284 25855 10286 25875
rect 10308 25855 10310 25875
rect 10332 25855 10334 25875
rect 10380 25855 10382 25875
rect 10404 25855 10406 25875
rect 10428 25855 10430 25875
rect 10476 25855 10478 25875
rect 10500 25855 10502 25875
rect 10524 25855 10526 25875
rect 10572 25855 10574 25875
rect 10596 25855 10598 25875
rect 10620 25855 10622 25875
rect 10668 25855 10670 25875
rect 10692 25855 10694 25875
rect 10716 25855 10718 25875
rect 10788 25855 10790 25875
rect 10836 25855 10838 25875
rect 10956 25855 10958 25875
rect 11004 25855 11006 25875
rect 11052 25855 11054 25875
rect 11076 25855 11078 25875
rect 11100 25855 11102 25875
rect 11172 25855 11174 25875
rect 11220 25855 11222 25875
rect 11340 25855 11342 25875
rect 11436 25855 11438 25875
rect 11532 25855 11534 25875
rect 11580 25855 11582 25875
rect 11628 25855 11630 25875
rect 11676 25855 11678 25875
rect 11724 25855 11726 25875
rect 11772 25855 11774 25875
rect 11796 25855 11798 25875
rect 11892 25855 11894 25875
rect 11988 25855 11990 25875
rect 12060 25855 12062 25875
rect 12132 25855 12134 25875
rect 12228 25855 12230 25875
rect 12276 25855 12278 25875
rect 12324 25855 12326 25875
rect 12420 25855 12422 25875
rect 12444 25855 12446 25875
rect 12492 25855 12494 25875
rect 12516 25855 12518 25875
rect 12540 25855 12542 25875
rect 12588 25855 12590 25875
rect 12636 25855 12638 25875
rect 12732 25855 12734 25875
rect 12756 25855 12758 25875
rect 12804 25855 12806 25875
rect 12828 25855 12830 25875
rect 12852 25855 12854 25875
rect 12900 25855 12902 25875
rect 12948 25855 12950 25875
rect 13044 25855 13046 25875
rect 13068 25855 13070 25875
rect 13116 25855 13118 25875
rect 13284 25855 13286 25875
rect 13332 25855 13334 25875
rect 13572 25855 13574 25875
rect 13644 25855 13646 25875
rect 13668 25855 13670 25875
rect 13764 25855 13766 25875
rect 13812 25855 13814 25875
rect 13860 25855 13862 25875
rect 13908 25855 13910 25875
rect 13956 25855 13958 25875
rect 14004 25855 14006 25875
rect 14100 25855 14102 25875
rect 14196 25855 14198 25875
rect 14292 25855 14294 25875
rect 15132 25855 15134 25875
rect 15180 25855 15182 25875
rect 15228 25855 15230 25875
rect 15252 25855 15254 25875
rect 15324 25855 15326 25875
rect 15396 25855 15398 25875
rect 15420 25855 15422 25875
rect 15492 25855 15494 25875
rect 15540 25855 15542 25875
rect 15636 25855 15638 25875
rect 15660 25855 15662 25875
rect 15708 25855 15710 25875
rect 15732 25855 15734 25875
rect 15756 25855 15758 25875
rect 15804 25855 15806 25875
rect 15828 25855 15830 25875
rect 15852 25855 15854 25875
rect 15900 25855 15902 25875
rect 15948 25855 15950 25875
rect 15996 25855 15998 25875
rect 16044 25855 16046 25875
rect 16164 25855 16166 25875
rect 16260 25855 16262 25875
rect 16308 25855 16310 25875
rect 16332 25855 16334 25875
rect 16356 25855 16358 25875
rect 16404 25855 16406 25875
rect 16452 25855 16454 25875
rect 16548 25855 16550 25875
rect 16572 25855 16574 25875
rect 16620 25855 16622 25875
rect 16668 25855 16670 25875
rect 16716 25855 16718 25875
rect 16764 25855 16766 25875
rect 16812 25855 16814 25875
rect 16884 25855 16886 25875
rect 16908 25855 16910 25875
rect 16980 25855 16982 25875
rect 17052 25855 17054 25875
rect 17196 25855 17198 25875
rect 17220 25855 17222 25875
rect 17292 25855 17294 25875
rect 17316 25855 17318 25875
rect 18084 25855 18086 25875
rect 18132 25855 18134 25875
rect 18217 25870 18220 25875
rect 18227 25856 18230 25870
rect 18228 25855 18230 25856
rect 18396 25855 18398 25875
rect 18492 25855 18494 25875
rect 18516 25855 18518 25875
rect 18564 25855 18566 25875
rect 18612 25855 18614 25875
rect 18660 25855 18662 25875
rect 18708 25855 18710 25875
rect 18756 25855 18758 25875
rect 18804 25855 18806 25875
rect 18852 25855 18854 25875
rect 18900 25855 18902 25875
rect 18996 25855 18998 25875
rect 19020 25855 19022 25875
rect 19092 25855 19094 25875
rect 19116 25855 19118 25875
rect 19140 25855 19142 25875
rect 19188 25855 19190 25875
rect 19236 25855 19238 25875
rect 19332 25855 19334 25875
rect 19476 25855 19478 25875
rect 19788 25855 19790 25875
rect 19836 25855 19838 25875
rect 19860 25855 19862 25875
rect 19884 25855 19886 25875
rect 19932 25855 19934 25875
rect 19956 25855 19958 25875
rect 19980 25855 19982 25875
rect 20028 25855 20030 25875
rect 20052 25855 20054 25875
rect 20076 25855 20078 25875
rect 20148 25855 20150 25875
rect 20172 25855 20174 25875
rect 20196 25855 20198 25875
rect 20268 25855 20270 25875
rect 20292 25855 20294 25875
rect 20388 25855 20390 25875
rect 20412 25855 20414 25875
rect 20508 25855 20510 25875
rect 20556 25855 20558 25875
rect 20604 25855 20606 25875
rect 20916 25855 20918 25875
rect 20929 25855 20963 25856
rect 20964 25855 20966 25875
rect 21012 25855 21014 25875
rect 21060 25855 21062 25875
rect 21084 25855 21086 25875
rect 21108 25855 21110 25875
rect 21204 25855 21206 25875
rect 21300 25855 21302 25875
rect 21324 25855 21326 25875
rect 21444 25855 21446 25875
rect 21468 25855 21470 25875
rect 21564 25855 21566 25875
rect 21612 25855 21614 25875
rect 21684 25855 21686 25875
rect 21708 25855 21710 25875
rect 21828 25855 21830 25875
rect 21924 25855 21926 25875
rect 22068 25855 22070 25875
rect 22188 25855 22190 25875
rect 22212 25855 22214 25875
rect 22884 25855 22886 25875
rect 22980 25855 22982 25875
rect 23076 25855 23078 25875
rect 23100 25855 23102 25875
rect 23124 25855 23126 25875
rect 23244 25855 23246 25875
rect 23340 25855 23342 25875
rect 23412 25855 23414 25875
rect 23508 25855 23510 25875
rect 23556 25855 23558 25875
rect 23652 25855 23654 25875
rect 23676 25855 23678 25875
rect 23724 25855 23726 25875
rect 23772 25855 23774 25875
rect 23820 25855 23822 25875
rect 23916 25855 23918 25875
rect 24012 25855 24014 25875
rect 24084 25855 24086 25875
rect 24396 25855 24398 25875
rect 24492 25855 24494 25875
rect 24516 25855 24518 25875
rect 24588 25855 24590 25875
rect 24612 25855 24614 25875
rect 24684 25855 24686 25875
rect 24732 25855 24734 25875
rect 24756 25855 24758 25875
rect 24780 25855 24782 25875
rect 24852 25855 24854 25875
rect 24876 25855 24878 25875
rect 24972 25855 24974 25875
rect 24996 25855 24998 25875
rect 25068 25855 25070 25875
rect 25164 25855 25166 25875
rect 25260 25855 25262 25875
rect 25308 25872 25310 25875
rect 25284 25855 25287 25872
rect 25308 25855 25311 25872
rect 25356 25855 25358 25875
rect 25380 25855 25382 25875
rect 25404 25855 25406 25875
rect 25500 25855 25502 25875
rect 25596 25855 25598 25875
rect 27036 25855 27038 25875
rect 27108 25855 27110 25875
rect 27324 25855 27326 25875
rect 27396 25855 27398 25875
rect 27420 25855 27422 25875
rect 27540 25856 27542 25875
rect 27553 25870 27556 25875
rect 27564 25870 27566 25875
rect 27563 25856 27566 25870
rect 27529 25855 27563 25856
rect -16761 25851 -12763 25855
rect -16761 25848 -16747 25851
rect -16740 25848 -16737 25851
rect -16692 25848 -16690 25851
rect -16692 25831 -16689 25848
rect -16524 25831 -16522 25851
rect -16404 25831 -16402 25851
rect -16356 25831 -16354 25851
rect -16319 25831 -16285 25832
rect -16713 25827 -16285 25831
rect -16713 25824 -16699 25827
rect -16692 25824 -16689 25827
rect -16524 25807 -16522 25827
rect -16404 25807 -16402 25827
rect -16356 25807 -16354 25827
rect -16319 25822 -16316 25827
rect -16309 25808 -16306 25822
rect -16308 25807 -16306 25808
rect -16284 25807 -16282 25851
rect -16260 25807 -16258 25851
rect -16247 25831 -16213 25832
rect -15324 25831 -15322 25851
rect -15215 25831 -15157 25832
rect -14772 25831 -14770 25851
rect -14508 25848 -14506 25851
rect -14508 25831 -14505 25848
rect -14436 25831 -14434 25851
rect -14340 25831 -14338 25851
rect -13980 25831 -13978 25851
rect -13932 25831 -13930 25851
rect -13884 25831 -13882 25851
rect -13788 25831 -13786 25851
rect -13572 25831 -13570 25851
rect -13356 25831 -13354 25851
rect -13284 25832 -13282 25851
rect -13319 25831 -13261 25832
rect -13068 25831 -13066 25851
rect -12780 25831 -12778 25851
rect -12777 25848 -12763 25851
rect -12756 25851 -9019 25855
rect -12756 25848 -12739 25851
rect -12756 25831 -12754 25848
rect -12660 25831 -12658 25851
rect -12564 25831 -12562 25851
rect -12492 25831 -12490 25851
rect -12396 25831 -12394 25851
rect -12348 25831 -12346 25851
rect -12252 25831 -12250 25851
rect -12156 25831 -12154 25851
rect -12060 25831 -12058 25851
rect -11844 25831 -11842 25851
rect -11796 25831 -11794 25851
rect -11676 25831 -11674 25851
rect -11591 25846 -11588 25851
rect -11580 25846 -11578 25851
rect -11581 25832 -11578 25846
rect -11556 25831 -11554 25851
rect -11508 25831 -11506 25851
rect -11471 25846 -11468 25851
rect -11460 25846 -11458 25851
rect -11461 25832 -11458 25846
rect -11436 25831 -11434 25851
rect -11412 25831 -11410 25851
rect -11364 25848 -11362 25851
rect -11364 25831 -11361 25848
rect -11340 25831 -11338 25851
rect -11196 25831 -11194 25851
rect -11124 25831 -11122 25851
rect -11100 25831 -11098 25851
rect -11028 25831 -11026 25851
rect -10740 25831 -10738 25851
rect -10668 25831 -10666 25851
rect -10644 25831 -10642 25851
rect -9996 25831 -9994 25851
rect -9828 25831 -9826 25851
rect -9732 25831 -9730 25851
rect -9612 25831 -9610 25851
rect -9516 25831 -9514 25851
rect -9468 25831 -9466 25851
rect -9420 25831 -9418 25851
rect -9407 25846 -9404 25851
rect -9396 25846 -9394 25851
rect -9397 25832 -9394 25846
rect -9300 25848 -9298 25851
rect -9300 25831 -9297 25848
rect -9252 25831 -9250 25851
rect -9033 25848 -9019 25851
rect -9009 25851 18317 25855
rect -9009 25848 -8995 25851
rect -8988 25848 -8985 25851
rect -8903 25846 -8900 25851
rect -8892 25846 -8890 25851
rect -8893 25832 -8890 25846
rect -8772 25832 -8770 25851
rect -8783 25831 -8749 25832
rect -8604 25831 -8602 25851
rect -8484 25831 -8482 25851
rect -8436 25831 -8434 25851
rect -8388 25831 -8386 25851
rect -8364 25831 -8362 25851
rect -8340 25831 -8338 25851
rect -8268 25831 -8266 25851
rect -8100 25831 -8098 25851
rect -8052 25831 -8050 25851
rect -7932 25831 -7930 25851
rect -7919 25831 -7885 25832
rect -7692 25831 -7690 25851
rect -7620 25831 -7618 25851
rect -7524 25831 -7522 25851
rect -7356 25831 -7354 25851
rect -7308 25831 -7306 25851
rect -7212 25831 -7210 25851
rect -7116 25831 -7114 25851
rect -7068 25831 -7066 25851
rect -6972 25831 -6970 25851
rect -6948 25831 -6946 25851
rect -6876 25831 -6874 25851
rect -6852 25831 -6850 25851
rect -6780 25831 -6778 25851
rect -6756 25831 -6754 25851
rect -6660 25831 -6658 25851
rect -6612 25831 -6610 25851
rect -6516 25831 -6514 25851
rect -6492 25832 -6490 25851
rect -6503 25831 -6469 25832
rect -6420 25831 -6418 25851
rect -6396 25831 -6394 25851
rect -6372 25831 -6370 25851
rect -6324 25831 -6322 25851
rect -6156 25831 -6154 25851
rect -6060 25831 -6058 25851
rect -6036 25831 -6034 25851
rect -5892 25831 -5890 25851
rect -5652 25831 -5650 25851
rect -5268 25831 -5266 25851
rect -5196 25831 -5194 25851
rect -5172 25831 -5170 25851
rect -5100 25831 -5098 25851
rect -5076 25831 -5074 25851
rect -4980 25831 -4978 25851
rect -4956 25831 -4954 25851
rect -4884 25832 -4882 25851
rect -4895 25831 -4861 25832
rect -4860 25831 -4858 25851
rect -4788 25831 -4786 25851
rect -4644 25831 -4642 25851
rect -4548 25831 -4546 25851
rect -4500 25831 -4498 25851
rect -4404 25831 -4402 25851
rect -4308 25831 -4306 25851
rect -4260 25831 -4258 25851
rect -4164 25831 -4162 25851
rect -4020 25831 -4018 25851
rect -3876 25831 -3874 25851
rect -3732 25831 -3730 25851
rect -3588 25831 -3586 25851
rect -3564 25831 -3562 25851
rect -3516 25831 -3514 25851
rect -3492 25831 -3490 25851
rect -3468 25831 -3466 25851
rect -3420 25831 -3418 25851
rect -3324 25831 -3322 25851
rect -3273 25848 -3259 25851
rect -3252 25848 -3249 25851
rect -3228 25831 -3226 25851
rect -3156 25831 -3154 25851
rect -3132 25831 -3130 25851
rect -3060 25831 -3058 25851
rect -3012 25831 -3010 25851
rect -2964 25831 -2962 25851
rect -2916 25831 -2914 25851
rect -2892 25831 -2890 25851
rect -2868 25831 -2866 25851
rect -2820 25831 -2818 25851
rect -2796 25831 -2794 25851
rect -2772 25831 -2770 25851
rect -2711 25846 -2708 25851
rect -2700 25846 -2698 25851
rect -2701 25832 -2698 25846
rect -2676 25831 -2674 25851
rect -2604 25848 -2602 25851
rect -2604 25831 -2601 25848
rect -2580 25831 -2578 25851
rect -2364 25831 -2362 25851
rect -2268 25831 -2266 25851
rect -2244 25831 -2242 25851
rect -2172 25831 -2170 25851
rect -2148 25831 -2146 25851
rect -2076 25831 -2074 25851
rect -2052 25831 -2050 25851
rect -1980 25831 -1978 25851
rect -1884 25831 -1882 25851
rect -1836 25831 -1834 25851
rect -1607 25846 -1604 25851
rect -1596 25846 -1594 25851
rect -1597 25832 -1594 25846
rect -1572 25831 -1570 25851
rect -1476 25831 -1474 25851
rect -1380 25831 -1378 25851
rect -1356 25831 -1354 25851
rect -1308 25831 -1306 25851
rect -1260 25831 -1258 25851
rect -1140 25831 -1138 25851
rect -852 25831 -850 25851
rect -756 25831 -754 25851
rect -708 25831 -706 25851
rect -612 25831 -610 25851
rect -588 25831 -586 25851
rect -540 25831 -538 25851
rect -492 25831 -490 25851
rect -444 25831 -442 25851
rect -396 25831 -394 25851
rect -300 25831 -298 25851
rect -276 25831 -274 25851
rect -228 25831 -226 25851
rect -12 25831 -10 25851
rect 156 25831 158 25851
rect 204 25831 206 25851
rect 217 25846 220 25851
rect 228 25846 230 25851
rect 227 25832 230 25846
rect 252 25831 254 25851
rect 348 25831 350 25851
rect 468 25831 470 25851
rect 492 25831 494 25851
rect 564 25831 566 25851
rect 588 25831 590 25851
rect 636 25831 638 25851
rect 660 25831 662 25851
rect 732 25831 734 25851
rect 745 25846 748 25851
rect 756 25846 758 25851
rect 755 25832 758 25846
rect 852 25848 854 25851
rect 852 25831 855 25848
rect 1020 25831 1022 25851
rect 1092 25831 1094 25851
rect 1116 25831 1118 25851
rect 1212 25831 1214 25851
rect 1308 25831 1310 25851
rect 1332 25831 1334 25851
rect 1380 25831 1382 25851
rect 1428 25831 1430 25851
rect 1476 25831 1478 25851
rect 1513 25846 1516 25851
rect 1524 25846 1526 25851
rect 1523 25832 1526 25846
rect 1548 25831 1550 25851
rect 1609 25846 1612 25851
rect 1620 25848 1622 25851
rect 1620 25846 1623 25848
rect 1619 25832 1623 25846
rect 1644 25831 1646 25851
rect 1692 25831 1694 25851
rect 1716 25848 1718 25851
rect 1716 25831 1719 25848
rect 1740 25831 1742 25851
rect 1788 25831 1790 25851
rect 2028 25831 2030 25851
rect 2076 25831 2078 25851
rect 2100 25831 2102 25851
rect 2124 25831 2126 25851
rect 2172 25831 2174 25851
rect 2196 25831 2198 25851
rect 2220 25831 2222 25851
rect 2268 25831 2270 25851
rect 2281 25846 2284 25851
rect 2292 25846 2294 25851
rect 2291 25832 2294 25846
rect 2316 25831 2318 25851
rect 2364 25831 2366 25851
rect 2412 25831 2414 25851
rect 2460 25831 2462 25851
rect 2508 25831 2510 25851
rect 2580 25831 2582 25851
rect 2604 25831 2606 25851
rect 2676 25831 2678 25851
rect 2700 25831 2702 25851
rect 2748 25831 2750 25851
rect 2772 25831 2774 25851
rect 2796 25831 2798 25851
rect 2844 25831 2846 25851
rect 2868 25831 2870 25851
rect 2892 25831 2894 25851
rect 2940 25831 2942 25851
rect 3012 25831 3014 25851
rect 3108 25831 3110 25851
rect 3156 25831 3158 25851
rect 3252 25831 3254 25851
rect 3348 25831 3350 25851
rect 3396 25831 3398 25851
rect 3468 25848 3470 25851
rect 3468 25831 3471 25848
rect 3481 25846 3484 25851
rect 3492 25846 3494 25851
rect 3491 25832 3494 25846
rect 3564 25831 3566 25851
rect 3612 25831 3614 25851
rect 3636 25831 3638 25851
rect 3660 25831 3662 25851
rect 3708 25831 3710 25851
rect 3732 25831 3734 25851
rect 3804 25831 3806 25851
rect 3828 25831 3830 25851
rect 3924 25831 3926 25851
rect 4020 25831 4022 25851
rect 4044 25831 4046 25851
rect 4092 25831 4094 25851
rect 4116 25831 4118 25851
rect 4140 25831 4142 25851
rect 4188 25831 4190 25851
rect 4212 25831 4214 25851
rect 4236 25831 4238 25851
rect 4308 25831 4310 25851
rect 4332 25831 4334 25851
rect 4404 25831 4406 25851
rect 4500 25831 4502 25851
rect 4596 25831 4598 25851
rect 4681 25846 4684 25851
rect 4691 25832 4694 25846
rect 4692 25831 4694 25832
rect 4860 25831 4862 25851
rect 4956 25831 4958 25851
rect 4980 25831 4982 25851
rect 5004 25831 5006 25851
rect 5076 25831 5078 25851
rect 5100 25831 5102 25851
rect 5124 25831 5126 25851
rect 5172 25831 5174 25851
rect 5220 25831 5222 25851
rect 5268 25831 5270 25851
rect 5388 25831 5390 25851
rect 5484 25831 5486 25851
rect 5508 25831 5510 25851
rect 5532 25831 5534 25851
rect 5628 25831 5630 25851
rect 5652 25831 5654 25851
rect 5748 25831 5750 25851
rect 5796 25831 5798 25851
rect 5844 25831 5846 25851
rect 5892 25831 5894 25851
rect 6132 25831 6134 25851
rect 6180 25831 6182 25851
rect 6228 25831 6230 25851
rect 6252 25831 6254 25851
rect 6276 25831 6278 25851
rect 6324 25831 6326 25851
rect 6372 25831 6374 25851
rect 6492 25831 6494 25851
rect 6588 25831 6590 25851
rect 6612 25831 6614 25851
rect 6660 25831 6662 25851
rect 6684 25831 6686 25851
rect 6708 25831 6710 25851
rect 6780 25831 6782 25851
rect 6804 25831 6806 25851
rect 6828 25831 6830 25851
rect 6900 25831 6902 25851
rect 6924 25831 6926 25851
rect 7020 25831 7022 25851
rect 7140 25831 7142 25851
rect 7236 25831 7238 25851
rect 7332 25831 7334 25851
rect 7380 25831 7382 25851
rect 7428 25831 7430 25851
rect 7452 25831 7454 25851
rect 7476 25831 7478 25851
rect 7524 25831 7526 25851
rect 7548 25831 7550 25851
rect 7572 25831 7574 25851
rect 7620 25831 7622 25851
rect 7644 25831 7646 25851
rect 7668 25831 7670 25851
rect 7740 25831 7742 25851
rect 7788 25831 7790 25851
rect 7884 25831 7886 25851
rect 7956 25831 7958 25851
rect 7980 25831 7982 25851
rect 8028 25831 8030 25851
rect 8196 25831 8198 25851
rect 8244 25831 8246 25851
rect 8268 25831 8270 25851
rect 8292 25831 8294 25851
rect 8340 25831 8342 25851
rect 8364 25831 8366 25851
rect 8388 25831 8390 25851
rect 8436 25831 8438 25851
rect 8460 25831 8462 25851
rect 8556 25831 8558 25851
rect 8604 25831 8606 25851
rect 8652 25831 8654 25851
rect 8700 25831 8702 25851
rect 8724 25831 8726 25851
rect 8748 25831 8750 25851
rect 8820 25831 8822 25851
rect 8844 25831 8846 25851
rect 8868 25831 8870 25851
rect 9516 25831 9518 25851
rect 9612 25831 9614 25851
rect 9660 25831 9662 25851
rect 9684 25831 9686 25851
rect 9708 25831 9710 25851
rect 9756 25831 9758 25851
rect 9780 25831 9782 25851
rect 9804 25831 9806 25851
rect 9852 25831 9854 25851
rect 9876 25831 9878 25851
rect 9900 25831 9902 25851
rect 9948 25831 9950 25851
rect 9972 25831 9974 25851
rect 9996 25831 9998 25851
rect 10068 25831 10070 25851
rect 10092 25831 10094 25851
rect 10116 25831 10118 25851
rect 10164 25831 10166 25851
rect 10188 25831 10190 25851
rect 10212 25831 10214 25851
rect 10284 25831 10286 25851
rect 10308 25831 10310 25851
rect 10332 25831 10334 25851
rect 10380 25831 10382 25851
rect 10404 25831 10406 25851
rect 10428 25831 10430 25851
rect 10476 25831 10478 25851
rect 10500 25831 10502 25851
rect 10524 25831 10526 25851
rect 10572 25831 10574 25851
rect 10596 25831 10598 25851
rect 10620 25831 10622 25851
rect 10668 25831 10670 25851
rect 10692 25831 10694 25851
rect 10716 25831 10718 25851
rect 10788 25831 10790 25851
rect 10836 25831 10838 25851
rect 10956 25831 10958 25851
rect 11004 25831 11006 25851
rect 11052 25831 11054 25851
rect 11076 25831 11078 25851
rect 11100 25831 11102 25851
rect 11172 25831 11174 25851
rect 11220 25831 11222 25851
rect 11340 25831 11342 25851
rect 11436 25831 11438 25851
rect 11532 25831 11534 25851
rect 11580 25831 11582 25851
rect 11628 25831 11630 25851
rect 11676 25831 11678 25851
rect 11724 25831 11726 25851
rect 11772 25831 11774 25851
rect 11796 25831 11798 25851
rect 11892 25831 11894 25851
rect 11988 25831 11990 25851
rect 12060 25831 12062 25851
rect 12132 25831 12134 25851
rect 12228 25831 12230 25851
rect 12276 25831 12278 25851
rect 12324 25831 12326 25851
rect 12420 25831 12422 25851
rect 12444 25831 12446 25851
rect 12492 25831 12494 25851
rect 12516 25831 12518 25851
rect 12540 25831 12542 25851
rect 12588 25831 12590 25851
rect 12636 25831 12638 25851
rect 12732 25831 12734 25851
rect 12756 25831 12758 25851
rect 12804 25831 12806 25851
rect 12828 25831 12830 25851
rect 12852 25831 12854 25851
rect 12900 25832 12902 25851
rect 12865 25831 12923 25832
rect 12948 25831 12950 25851
rect 13044 25831 13046 25851
rect 13068 25831 13070 25851
rect 13116 25831 13118 25851
rect 13284 25831 13286 25851
rect 13332 25831 13334 25851
rect 13572 25831 13574 25851
rect 13644 25831 13646 25851
rect 13668 25831 13670 25851
rect 13764 25831 13766 25851
rect 13812 25831 13814 25851
rect 13860 25831 13862 25851
rect 13908 25831 13910 25851
rect 13956 25831 13958 25851
rect 14004 25831 14006 25851
rect 14100 25831 14102 25851
rect 14196 25831 14198 25851
rect 14292 25831 14294 25851
rect 15132 25831 15134 25851
rect 15180 25831 15182 25851
rect 15228 25831 15230 25851
rect 15252 25831 15254 25851
rect 15324 25831 15326 25851
rect 15396 25831 15398 25851
rect 15420 25831 15422 25851
rect 15492 25831 15494 25851
rect 15540 25831 15542 25851
rect 15636 25831 15638 25851
rect 15660 25831 15662 25851
rect 15708 25831 15710 25851
rect 15732 25831 15734 25851
rect 15756 25831 15758 25851
rect 15804 25831 15806 25851
rect 15828 25831 15830 25851
rect 15852 25831 15854 25851
rect 15900 25831 15902 25851
rect 15948 25831 15950 25851
rect 15996 25831 15998 25851
rect 16044 25831 16046 25851
rect 16164 25831 16166 25851
rect 16260 25831 16262 25851
rect 16308 25831 16310 25851
rect 16332 25831 16334 25851
rect 16356 25831 16358 25851
rect 16404 25831 16406 25851
rect 16452 25831 16454 25851
rect 16548 25831 16550 25851
rect 16572 25831 16574 25851
rect 16620 25831 16622 25851
rect 16668 25831 16670 25851
rect 16716 25831 16718 25851
rect 16764 25831 16766 25851
rect 16812 25831 16814 25851
rect 16884 25831 16886 25851
rect 16908 25831 16910 25851
rect 16980 25831 16982 25851
rect 17052 25831 17054 25851
rect 17196 25831 17198 25851
rect 17220 25831 17222 25851
rect 17292 25831 17294 25851
rect 17316 25831 17318 25851
rect 18084 25831 18086 25851
rect 18132 25831 18134 25851
rect 18228 25831 18230 25851
rect 18303 25848 18317 25851
rect 18327 25851 25277 25855
rect 18327 25848 18341 25851
rect 18396 25831 18398 25851
rect 18492 25831 18494 25851
rect 18516 25831 18518 25851
rect 18564 25831 18566 25851
rect 18612 25831 18614 25851
rect 18660 25831 18662 25851
rect 18708 25831 18710 25851
rect 18756 25831 18758 25851
rect 18804 25831 18806 25851
rect 18852 25831 18854 25851
rect 18900 25831 18902 25851
rect 18996 25831 18998 25851
rect 19020 25831 19022 25851
rect 19092 25831 19094 25851
rect 19116 25831 19118 25851
rect 19140 25831 19142 25851
rect 19188 25831 19190 25851
rect 19236 25831 19238 25851
rect 19332 25831 19334 25851
rect 19476 25831 19478 25851
rect 19788 25831 19790 25851
rect 19836 25831 19838 25851
rect 19860 25831 19862 25851
rect 19884 25831 19886 25851
rect 19932 25831 19934 25851
rect 19956 25831 19958 25851
rect 19980 25831 19982 25851
rect 20028 25831 20030 25851
rect 20052 25831 20054 25851
rect 20076 25831 20078 25851
rect 20148 25831 20150 25851
rect 20172 25831 20174 25851
rect 20196 25831 20198 25851
rect 20268 25831 20270 25851
rect 20292 25831 20294 25851
rect 20388 25831 20390 25851
rect 20412 25831 20414 25851
rect 20508 25831 20510 25851
rect 20556 25831 20558 25851
rect 20604 25831 20606 25851
rect 20916 25831 20918 25851
rect 20964 25831 20966 25851
rect 21012 25831 21014 25851
rect 21060 25831 21062 25851
rect 21084 25831 21086 25851
rect 21108 25831 21110 25851
rect 21204 25831 21206 25851
rect 21300 25831 21302 25851
rect 21324 25831 21326 25851
rect 21444 25831 21446 25851
rect 21468 25831 21470 25851
rect 21564 25831 21566 25851
rect 21612 25831 21614 25851
rect 21684 25831 21686 25851
rect 21708 25831 21710 25851
rect 21828 25831 21830 25851
rect 21924 25831 21926 25851
rect 22068 25831 22070 25851
rect 22188 25831 22190 25851
rect 22212 25831 22214 25851
rect 22884 25831 22886 25851
rect 22980 25831 22982 25851
rect 23076 25831 23078 25851
rect 23100 25831 23102 25851
rect 23124 25831 23126 25851
rect 23244 25831 23246 25851
rect 23340 25831 23342 25851
rect 23412 25831 23414 25851
rect 23508 25831 23510 25851
rect 23556 25831 23558 25851
rect 23652 25831 23654 25851
rect 23676 25831 23678 25851
rect 23724 25831 23726 25851
rect 23772 25831 23774 25851
rect 23820 25831 23822 25851
rect 23916 25831 23918 25851
rect 24012 25831 24014 25851
rect 24084 25831 24086 25851
rect 24396 25831 24398 25851
rect 24492 25831 24494 25851
rect 24516 25831 24518 25851
rect 24588 25831 24590 25851
rect 24612 25831 24614 25851
rect 24684 25831 24686 25851
rect 24732 25831 24734 25851
rect 24756 25831 24758 25851
rect 24780 25831 24782 25851
rect 24852 25831 24854 25851
rect 24876 25831 24878 25851
rect 24972 25831 24974 25851
rect 24996 25831 24998 25851
rect 25068 25831 25070 25851
rect 25164 25831 25166 25851
rect 25260 25831 25262 25851
rect 25263 25848 25277 25851
rect 25284 25851 27563 25855
rect 25284 25848 25301 25851
rect 25308 25848 25311 25851
rect 25284 25831 25286 25848
rect 25356 25831 25358 25851
rect 25380 25831 25382 25851
rect 25404 25831 25406 25851
rect 25500 25831 25502 25851
rect 25596 25831 25598 25851
rect 27036 25831 27038 25851
rect 27108 25831 27110 25851
rect 27324 25831 27326 25851
rect 27396 25831 27398 25851
rect 27420 25831 27422 25851
rect 27529 25846 27532 25851
rect 27540 25846 27542 25851
rect 27539 25832 27542 25846
rect 27457 25831 27491 25832
rect -16247 25827 4781 25831
rect -16223 25814 -16219 25822
rect -16233 25808 -16223 25814
rect -15324 25807 -15322 25827
rect -15108 25807 -15105 25824
rect -14772 25807 -14770 25827
rect -14529 25824 -14515 25827
rect -14508 25824 -14505 25827
rect -14436 25807 -14434 25827
rect -14340 25807 -14338 25827
rect -13980 25807 -13978 25827
rect -13932 25807 -13930 25827
rect -13884 25807 -13882 25827
rect -13788 25807 -13786 25827
rect -13572 25807 -13570 25827
rect -13356 25807 -13354 25827
rect -13295 25822 -13292 25827
rect -13284 25822 -13282 25827
rect -13285 25808 -13282 25822
rect -13068 25807 -13066 25827
rect -12780 25807 -12778 25827
rect -12756 25807 -12754 25827
rect -12660 25807 -12658 25827
rect -12564 25807 -12562 25827
rect -12492 25807 -12490 25827
rect -12396 25807 -12394 25827
rect -12348 25807 -12346 25827
rect -12252 25807 -12250 25827
rect -12156 25807 -12154 25827
rect -12060 25807 -12058 25827
rect -11844 25807 -11842 25827
rect -11796 25808 -11794 25827
rect -11807 25807 -11773 25808
rect -11676 25807 -11674 25827
rect -11556 25807 -11554 25827
rect -11508 25807 -11506 25827
rect -11505 25824 -11491 25827
rect -11436 25807 -11434 25827
rect -11412 25807 -11410 25827
rect -11385 25824 -11371 25827
rect -11364 25824 -11361 25827
rect -11340 25807 -11338 25827
rect -11196 25807 -11194 25827
rect -11124 25807 -11122 25827
rect -11100 25807 -11098 25827
rect -11028 25807 -11026 25827
rect -10740 25807 -10738 25827
rect -10668 25807 -10666 25827
rect -10644 25807 -10642 25827
rect -9996 25807 -9994 25827
rect -9828 25807 -9826 25827
rect -9732 25807 -9730 25827
rect -9612 25807 -9610 25827
rect -9516 25807 -9514 25827
rect -9468 25807 -9466 25827
rect -9420 25807 -9418 25827
rect -9321 25824 -9307 25827
rect -9300 25824 -9297 25827
rect -9252 25807 -9250 25827
rect -8817 25824 -8803 25827
rect -8783 25822 -8780 25827
rect -8772 25822 -8770 25827
rect -8773 25808 -8770 25822
rect -8604 25807 -8602 25827
rect -8484 25807 -8482 25827
rect -8436 25807 -8434 25827
rect -8388 25807 -8386 25827
rect -8364 25807 -8362 25827
rect -8340 25807 -8338 25827
rect -8268 25807 -8266 25827
rect -8100 25807 -8098 25827
rect -8052 25807 -8050 25827
rect -7932 25807 -7930 25827
rect -7692 25807 -7690 25827
rect -7620 25807 -7618 25827
rect -7524 25807 -7522 25827
rect -7356 25807 -7354 25827
rect -7308 25807 -7306 25827
rect -7212 25807 -7210 25827
rect -7116 25807 -7114 25827
rect -7068 25807 -7066 25827
rect -6972 25807 -6970 25827
rect -6948 25807 -6946 25827
rect -6876 25807 -6874 25827
rect -6852 25807 -6850 25827
rect -6780 25807 -6778 25827
rect -6756 25807 -6754 25827
rect -6660 25807 -6658 25827
rect -6612 25807 -6610 25827
rect -6516 25807 -6514 25827
rect -6503 25822 -6500 25827
rect -6492 25822 -6490 25827
rect -6493 25808 -6490 25822
rect -6420 25807 -6418 25827
rect -6396 25824 -6394 25827
rect -6396 25807 -6393 25824
rect -6372 25807 -6370 25827
rect -6324 25807 -6322 25827
rect -6156 25807 -6154 25827
rect -6060 25807 -6058 25827
rect -6036 25807 -6034 25827
rect -5892 25807 -5890 25827
rect -5652 25807 -5650 25827
rect -5268 25807 -5266 25827
rect -5196 25807 -5194 25827
rect -5172 25807 -5170 25827
rect -5100 25807 -5098 25827
rect -5076 25807 -5074 25827
rect -4980 25807 -4978 25827
rect -4956 25807 -4954 25827
rect -4895 25822 -4892 25827
rect -4884 25822 -4882 25827
rect -4885 25808 -4882 25822
rect -4860 25807 -4858 25827
rect -4788 25824 -4786 25827
rect -4788 25807 -4785 25824
rect -4644 25807 -4642 25827
rect -4548 25807 -4546 25827
rect -4500 25807 -4498 25827
rect -4404 25807 -4402 25827
rect -4308 25807 -4306 25827
rect -4260 25807 -4258 25827
rect -4164 25807 -4162 25827
rect -4020 25807 -4018 25827
rect -3876 25807 -3874 25827
rect -3732 25807 -3730 25827
rect -3588 25807 -3586 25827
rect -3564 25807 -3562 25827
rect -3516 25807 -3514 25827
rect -3492 25807 -3490 25827
rect -3468 25807 -3466 25827
rect -3420 25807 -3418 25827
rect -3324 25807 -3322 25827
rect -3228 25807 -3226 25827
rect -3156 25807 -3154 25827
rect -3132 25807 -3130 25827
rect -3060 25807 -3058 25827
rect -3012 25807 -3010 25827
rect -2964 25807 -2962 25827
rect -2916 25807 -2914 25827
rect -2892 25807 -2890 25827
rect -2868 25807 -2866 25827
rect -2820 25807 -2818 25827
rect -2796 25807 -2794 25827
rect -2772 25807 -2770 25827
rect -2676 25807 -2674 25827
rect -2625 25824 -2611 25827
rect -2604 25824 -2601 25827
rect -2580 25807 -2578 25827
rect -2364 25807 -2362 25827
rect -2268 25807 -2266 25827
rect -2244 25807 -2242 25827
rect -2172 25807 -2170 25827
rect -2148 25807 -2146 25827
rect -2076 25807 -2074 25827
rect -2052 25807 -2050 25827
rect -1980 25807 -1978 25827
rect -1884 25807 -1882 25827
rect -1836 25807 -1834 25827
rect -1572 25807 -1570 25827
rect -1521 25824 -1507 25827
rect -1476 25807 -1474 25827
rect -1380 25807 -1378 25827
rect -1356 25807 -1354 25827
rect -1308 25807 -1306 25827
rect -1260 25807 -1258 25827
rect -1140 25807 -1138 25827
rect -852 25807 -850 25827
rect -756 25807 -754 25827
rect -708 25807 -706 25827
rect -612 25807 -610 25827
rect -588 25807 -586 25827
rect -540 25807 -538 25827
rect -492 25807 -490 25827
rect -444 25807 -442 25827
rect -396 25807 -394 25827
rect -300 25807 -298 25827
rect -276 25807 -274 25827
rect -228 25807 -226 25827
rect -12 25807 -10 25827
rect 156 25807 158 25827
rect 204 25807 206 25827
rect 252 25807 254 25827
rect 303 25824 317 25827
rect 348 25807 350 25827
rect 468 25807 470 25827
rect 492 25807 494 25827
rect 564 25807 566 25827
rect 588 25807 590 25827
rect 636 25807 638 25827
rect 660 25807 662 25827
rect 732 25807 734 25827
rect 831 25824 845 25827
rect 852 25824 855 25827
rect 1020 25807 1022 25827
rect 1092 25807 1094 25827
rect 1116 25807 1118 25827
rect 1212 25807 1214 25827
rect 1308 25807 1310 25827
rect 1332 25807 1334 25827
rect 1380 25807 1382 25827
rect 1428 25807 1430 25827
rect 1476 25807 1478 25827
rect 1548 25807 1550 25827
rect 1599 25824 1613 25827
rect 1644 25807 1646 25827
rect 1692 25807 1694 25827
rect 1695 25824 1709 25827
rect 1716 25824 1719 25827
rect 1740 25807 1742 25827
rect 1788 25807 1790 25827
rect 2028 25807 2030 25827
rect 2076 25807 2078 25827
rect 2100 25807 2102 25827
rect 2124 25807 2126 25827
rect 2172 25807 2174 25827
rect 2196 25808 2198 25827
rect 2185 25807 2219 25808
rect 2220 25807 2222 25827
rect 2268 25807 2270 25827
rect 2316 25807 2318 25827
rect 2364 25807 2366 25827
rect 2367 25824 2381 25827
rect 2412 25807 2414 25827
rect 2460 25807 2462 25827
rect 2508 25807 2510 25827
rect 2580 25807 2582 25827
rect 2604 25807 2606 25827
rect 2676 25807 2678 25827
rect 2700 25807 2702 25827
rect 2748 25807 2750 25827
rect 2772 25807 2774 25827
rect 2796 25807 2798 25827
rect 2844 25807 2846 25827
rect 2868 25807 2870 25827
rect 2892 25807 2894 25827
rect 2940 25807 2942 25827
rect 3012 25807 3014 25827
rect 3108 25807 3110 25827
rect 3156 25807 3158 25827
rect 3207 25824 3221 25827
rect 3252 25807 3254 25827
rect 3348 25807 3350 25827
rect 3396 25807 3398 25827
rect 3447 25824 3461 25827
rect 3468 25824 3471 25827
rect 3564 25807 3566 25827
rect 3567 25824 3581 25827
rect 3612 25807 3614 25827
rect 3636 25807 3638 25827
rect 3660 25807 3662 25827
rect 3708 25807 3710 25827
rect 3732 25807 3734 25827
rect 3804 25807 3806 25827
rect 3828 25807 3830 25827
rect 3924 25807 3926 25827
rect 4020 25807 4022 25827
rect 4044 25807 4046 25827
rect 4092 25807 4094 25827
rect 4116 25807 4118 25827
rect 4140 25807 4142 25827
rect 4188 25807 4190 25827
rect 4212 25807 4214 25827
rect 4236 25807 4238 25827
rect 4308 25807 4310 25827
rect 4332 25807 4334 25827
rect 4404 25807 4406 25827
rect 4500 25807 4502 25827
rect 4596 25807 4598 25827
rect 4692 25807 4694 25827
rect 4767 25824 4781 25827
rect 4791 25827 27491 25831
rect 4791 25824 4805 25827
rect 4860 25807 4862 25827
rect 4956 25807 4958 25827
rect 4980 25807 4982 25827
rect 5004 25807 5006 25827
rect 5076 25807 5078 25827
rect 5100 25807 5102 25827
rect 5124 25807 5126 25827
rect 5172 25807 5174 25827
rect 5220 25807 5222 25827
rect 5268 25807 5270 25827
rect 5388 25807 5390 25827
rect 5484 25807 5486 25827
rect 5508 25807 5510 25827
rect 5532 25807 5534 25827
rect 5628 25807 5630 25827
rect 5652 25807 5654 25827
rect 5748 25807 5750 25827
rect 5796 25807 5798 25827
rect 5844 25807 5846 25827
rect 5892 25807 5894 25827
rect 6132 25807 6134 25827
rect 6180 25807 6182 25827
rect 6228 25807 6230 25827
rect 6252 25807 6254 25827
rect 6276 25807 6278 25827
rect 6324 25807 6326 25827
rect 6372 25807 6374 25827
rect 6492 25807 6494 25827
rect 6588 25807 6590 25827
rect 6612 25807 6614 25827
rect 6660 25807 6662 25827
rect 6684 25807 6686 25827
rect 6708 25807 6710 25827
rect 6721 25807 6755 25808
rect 6780 25807 6782 25827
rect 6804 25807 6806 25827
rect 6828 25807 6830 25827
rect 6900 25807 6902 25827
rect 6924 25807 6926 25827
rect 7020 25807 7022 25827
rect 7140 25807 7142 25827
rect 7236 25807 7238 25827
rect 7332 25807 7334 25827
rect 7380 25807 7382 25827
rect 7428 25807 7430 25827
rect 7452 25807 7454 25827
rect 7476 25807 7478 25827
rect 7524 25807 7526 25827
rect 7548 25807 7550 25827
rect 7572 25807 7574 25827
rect 7620 25807 7622 25827
rect 7644 25807 7646 25827
rect 7668 25807 7670 25827
rect 7740 25807 7742 25827
rect 7788 25807 7790 25827
rect 7884 25807 7886 25827
rect 7956 25807 7958 25827
rect 7980 25807 7982 25827
rect 8028 25807 8030 25827
rect 8196 25807 8198 25827
rect 8244 25807 8246 25827
rect 8268 25807 8270 25827
rect 8292 25807 8294 25827
rect 8340 25807 8342 25827
rect 8364 25807 8366 25827
rect 8388 25807 8390 25827
rect 8436 25807 8438 25827
rect 8460 25807 8462 25827
rect 8556 25807 8558 25827
rect 8604 25807 8606 25827
rect 8652 25807 8654 25827
rect 8700 25807 8702 25827
rect 8724 25807 8726 25827
rect 8748 25807 8750 25827
rect 8820 25807 8822 25827
rect 8844 25807 8846 25827
rect 8868 25807 8870 25827
rect 9516 25807 9518 25827
rect 9612 25807 9614 25827
rect 9660 25807 9662 25827
rect 9684 25807 9686 25827
rect 9708 25807 9710 25827
rect 9756 25807 9758 25827
rect 9780 25807 9782 25827
rect 9804 25807 9806 25827
rect 9852 25807 9854 25827
rect 9876 25808 9878 25827
rect 9865 25807 9899 25808
rect 9900 25807 9902 25827
rect 9948 25807 9950 25827
rect 9972 25807 9974 25827
rect 9996 25807 9998 25827
rect 10068 25807 10070 25827
rect 10092 25807 10094 25827
rect 10116 25807 10118 25827
rect 10164 25807 10166 25827
rect 10188 25807 10190 25827
rect 10212 25807 10214 25827
rect 10284 25807 10286 25827
rect 10308 25807 10310 25827
rect 10332 25807 10334 25827
rect 10380 25807 10382 25827
rect 10404 25807 10406 25827
rect 10428 25807 10430 25827
rect 10476 25807 10478 25827
rect 10500 25807 10502 25827
rect 10524 25807 10526 25827
rect 10572 25807 10574 25827
rect 10596 25807 10598 25827
rect 10620 25807 10622 25827
rect 10668 25807 10670 25827
rect 10692 25807 10694 25827
rect 10716 25807 10718 25827
rect 10788 25807 10790 25827
rect 10836 25807 10838 25827
rect 10956 25807 10958 25827
rect 11004 25807 11006 25827
rect 11052 25807 11054 25827
rect 11076 25807 11078 25827
rect 11100 25807 11102 25827
rect 11172 25807 11174 25827
rect 11220 25807 11222 25827
rect 11340 25807 11342 25827
rect 11436 25807 11438 25827
rect 11532 25807 11534 25827
rect 11580 25807 11582 25827
rect 11628 25807 11630 25827
rect 11676 25807 11678 25827
rect 11724 25807 11726 25827
rect 11772 25807 11774 25827
rect 11796 25807 11798 25827
rect 11892 25807 11894 25827
rect 11988 25807 11990 25827
rect 12060 25807 12062 25827
rect 12132 25807 12134 25827
rect 12228 25807 12230 25827
rect 12276 25807 12278 25827
rect 12324 25807 12326 25827
rect 12420 25807 12422 25827
rect 12444 25807 12446 25827
rect 12492 25807 12494 25827
rect 12516 25807 12518 25827
rect 12540 25807 12542 25827
rect 12588 25807 12590 25827
rect 12636 25807 12638 25827
rect 12732 25807 12734 25827
rect 12756 25807 12758 25827
rect 12804 25807 12806 25827
rect 12828 25807 12830 25827
rect 12852 25807 12854 25827
rect 12889 25822 12892 25827
rect 12900 25822 12902 25827
rect 12899 25808 12902 25822
rect 12948 25807 12950 25827
rect 12972 25807 12975 25824
rect 13044 25807 13046 25827
rect 13068 25807 13070 25827
rect 13116 25807 13118 25827
rect 13284 25807 13286 25827
rect 13332 25807 13334 25827
rect 13572 25807 13574 25827
rect 13644 25807 13646 25827
rect 13668 25807 13670 25827
rect 13764 25807 13766 25827
rect 13812 25807 13814 25827
rect 13860 25807 13862 25827
rect 13908 25807 13910 25827
rect 13956 25807 13958 25827
rect 14004 25807 14006 25827
rect 14100 25807 14102 25827
rect 14196 25807 14198 25827
rect 14292 25807 14294 25827
rect 15132 25808 15134 25827
rect 15121 25807 15155 25808
rect 15180 25807 15182 25827
rect 15228 25808 15230 25827
rect 15217 25807 15251 25808
rect 15252 25807 15254 25827
rect 15265 25807 15323 25808
rect 15324 25807 15326 25827
rect 15396 25807 15398 25827
rect 15420 25807 15422 25827
rect 15492 25807 15494 25827
rect 15540 25807 15542 25827
rect 15636 25807 15638 25827
rect 15660 25807 15662 25827
rect 15708 25807 15710 25827
rect 15732 25807 15734 25827
rect 15756 25807 15758 25827
rect 15804 25807 15806 25827
rect 15828 25807 15830 25827
rect 15852 25807 15854 25827
rect 15900 25807 15902 25827
rect 15948 25807 15950 25827
rect 15996 25807 15998 25827
rect 16044 25807 16046 25827
rect 16164 25807 16166 25827
rect 16260 25807 16262 25827
rect 16308 25807 16310 25827
rect 16332 25807 16334 25827
rect 16356 25807 16358 25827
rect 16404 25807 16406 25827
rect 16452 25807 16454 25827
rect 16548 25807 16550 25827
rect 16572 25807 16574 25827
rect 16620 25807 16622 25827
rect 16668 25807 16670 25827
rect 16716 25807 16718 25827
rect 16764 25807 16766 25827
rect 16812 25807 16814 25827
rect 16884 25807 16886 25827
rect 16908 25807 16910 25827
rect 16980 25807 16982 25827
rect 17052 25807 17054 25827
rect 17196 25807 17198 25827
rect 17220 25807 17222 25827
rect 17292 25807 17294 25827
rect 17316 25807 17318 25827
rect 18084 25807 18086 25827
rect 18132 25807 18134 25827
rect 18228 25807 18230 25827
rect 18396 25807 18398 25827
rect 18492 25807 18494 25827
rect 18516 25807 18518 25827
rect 18564 25807 18566 25827
rect 18612 25807 18614 25827
rect 18660 25807 18662 25827
rect 18708 25807 18710 25827
rect 18756 25807 18758 25827
rect 18804 25807 18806 25827
rect 18852 25807 18854 25827
rect 18900 25807 18902 25827
rect 18996 25807 18998 25827
rect 19020 25807 19022 25827
rect 19092 25807 19094 25827
rect 19116 25807 19118 25827
rect 19140 25807 19142 25827
rect 19188 25807 19190 25827
rect 19236 25807 19238 25827
rect 19332 25807 19334 25827
rect 19476 25807 19478 25827
rect 19788 25807 19790 25827
rect 19836 25807 19838 25827
rect 19860 25807 19862 25827
rect 19884 25807 19886 25827
rect 19932 25807 19934 25827
rect 19956 25807 19958 25827
rect 19980 25807 19982 25827
rect 20028 25807 20030 25827
rect 20052 25807 20054 25827
rect 20076 25807 20078 25827
rect 20148 25807 20150 25827
rect 20172 25807 20174 25827
rect 20196 25807 20198 25827
rect 20268 25807 20270 25827
rect 20292 25807 20294 25827
rect 20388 25807 20390 25827
rect 20412 25807 20414 25827
rect 20508 25807 20510 25827
rect 20556 25807 20558 25827
rect 20604 25807 20606 25827
rect 20916 25807 20918 25827
rect 20964 25807 20966 25827
rect 21012 25807 21014 25827
rect 21015 25824 21029 25827
rect 21060 25807 21062 25827
rect 21084 25807 21086 25827
rect 21108 25807 21110 25827
rect 21204 25807 21206 25827
rect 21300 25807 21302 25827
rect 21324 25807 21326 25827
rect 21444 25807 21446 25827
rect 21468 25807 21470 25827
rect 21564 25807 21566 25827
rect 21612 25807 21614 25827
rect 21684 25807 21686 25827
rect 21708 25807 21710 25827
rect 21828 25807 21830 25827
rect 21924 25807 21926 25827
rect 22068 25807 22070 25827
rect 22188 25807 22190 25827
rect 22212 25807 22214 25827
rect 22884 25807 22886 25827
rect 22980 25807 22982 25827
rect 23076 25807 23078 25827
rect 23100 25807 23102 25827
rect 23124 25807 23126 25827
rect 23244 25807 23246 25827
rect 23340 25807 23342 25827
rect 23412 25807 23414 25827
rect 23508 25807 23510 25827
rect 23556 25807 23558 25827
rect 23652 25807 23654 25827
rect 23676 25807 23678 25827
rect 23724 25807 23726 25827
rect 23772 25807 23774 25827
rect 23820 25807 23822 25827
rect 23916 25807 23918 25827
rect 24012 25807 24014 25827
rect 24084 25807 24086 25827
rect 24396 25807 24398 25827
rect 24492 25807 24494 25827
rect 24516 25807 24518 25827
rect 24588 25807 24590 25827
rect 24612 25807 24614 25827
rect 24684 25807 24686 25827
rect 24732 25807 24734 25827
rect 24756 25807 24758 25827
rect 24780 25807 24782 25827
rect 24852 25807 24854 25827
rect 24876 25807 24878 25827
rect 24972 25807 24974 25827
rect 24996 25807 24998 25827
rect 25068 25807 25070 25827
rect 25164 25807 25166 25827
rect 25260 25807 25262 25827
rect 25284 25807 25286 25827
rect 25356 25807 25358 25827
rect 25380 25807 25382 25827
rect 25404 25807 25406 25827
rect 25500 25807 25502 25827
rect 25596 25807 25598 25827
rect 27036 25807 27038 25827
rect 27108 25807 27110 25827
rect 27324 25807 27326 25827
rect 27396 25807 27398 25827
rect 27420 25807 27422 25827
rect 27433 25807 27467 25808
rect -16665 25803 -16219 25807
rect -16665 25800 -16651 25803
rect -16617 25783 -16597 25784
rect -16524 25783 -16522 25803
rect -16404 25783 -16402 25803
rect -16356 25783 -16354 25803
rect -16308 25783 -16306 25803
rect -16284 25783 -16282 25803
rect -16260 25783 -16258 25803
rect -16233 25800 -16219 25803
rect -16161 25803 -15115 25807
rect -16161 25800 -16147 25803
rect -15324 25783 -15322 25803
rect -15129 25800 -15115 25803
rect -15108 25803 -13219 25807
rect -15108 25800 -15091 25803
rect -15108 25783 -15106 25800
rect -14772 25783 -14770 25803
rect -14436 25783 -14434 25803
rect -14340 25783 -14338 25803
rect -14279 25783 -14245 25784
rect -13980 25783 -13978 25803
rect -13932 25783 -13930 25803
rect -13884 25783 -13882 25803
rect -13788 25783 -13786 25803
rect -13572 25783 -13570 25803
rect -13356 25783 -13354 25803
rect -13233 25800 -13219 25803
rect -13209 25803 12965 25807
rect -13209 25800 -13195 25803
rect -13068 25783 -13066 25803
rect -12780 25783 -12778 25803
rect -12756 25783 -12754 25803
rect -12660 25783 -12658 25803
rect -12564 25783 -12562 25803
rect -12492 25783 -12490 25803
rect -12396 25783 -12394 25803
rect -12348 25783 -12346 25803
rect -12252 25783 -12250 25803
rect -12156 25783 -12154 25803
rect -12060 25783 -12058 25803
rect -11844 25783 -11842 25803
rect -11807 25798 -11804 25803
rect -11796 25798 -11794 25803
rect -11797 25784 -11794 25798
rect -11676 25783 -11674 25803
rect -11556 25783 -11554 25803
rect -11508 25783 -11506 25803
rect -11436 25783 -11434 25803
rect -11412 25783 -11410 25803
rect -11340 25783 -11338 25803
rect -11196 25783 -11194 25803
rect -11124 25783 -11122 25803
rect -11100 25783 -11098 25803
rect -11028 25783 -11026 25803
rect -10740 25783 -10738 25803
rect -10668 25783 -10666 25803
rect -10644 25783 -10642 25803
rect -9996 25783 -9994 25803
rect -9828 25783 -9826 25803
rect -9732 25783 -9730 25803
rect -9719 25783 -9685 25784
rect -9612 25783 -9610 25803
rect -9516 25783 -9514 25803
rect -9468 25783 -9466 25803
rect -9420 25783 -9418 25803
rect -9252 25783 -9250 25803
rect -8697 25800 -8683 25803
rect -8604 25783 -8602 25803
rect -8484 25783 -8482 25803
rect -8436 25783 -8434 25803
rect -8388 25783 -8386 25803
rect -8364 25783 -8362 25803
rect -8340 25783 -8338 25803
rect -8268 25783 -8266 25803
rect -8100 25783 -8098 25803
rect -8052 25783 -8050 25803
rect -7932 25783 -7930 25803
rect -7833 25800 -7819 25803
rect -7692 25783 -7690 25803
rect -7620 25783 -7618 25803
rect -7524 25783 -7522 25803
rect -7356 25783 -7354 25803
rect -7308 25783 -7306 25803
rect -7212 25783 -7210 25803
rect -7116 25783 -7114 25803
rect -7068 25783 -7066 25803
rect -6972 25783 -6970 25803
rect -6948 25783 -6946 25803
rect -6876 25783 -6874 25803
rect -6852 25783 -6850 25803
rect -6780 25783 -6778 25803
rect -6756 25783 -6754 25803
rect -6660 25783 -6658 25803
rect -6612 25783 -6610 25803
rect -6516 25783 -6514 25803
rect -6420 25783 -6418 25803
rect -6417 25800 -6403 25803
rect -6396 25800 -6393 25803
rect -6372 25783 -6370 25803
rect -6324 25783 -6322 25803
rect -6156 25783 -6154 25803
rect -6060 25783 -6058 25803
rect -6036 25783 -6034 25803
rect -5892 25783 -5890 25803
rect -5652 25783 -5650 25803
rect -5268 25783 -5266 25803
rect -5196 25783 -5194 25803
rect -5172 25783 -5170 25803
rect -5100 25783 -5098 25803
rect -5076 25783 -5074 25803
rect -4980 25783 -4978 25803
rect -4956 25783 -4954 25803
rect -4860 25783 -4858 25803
rect -4809 25800 -4795 25803
rect -4788 25800 -4785 25803
rect -4644 25783 -4642 25803
rect -4548 25783 -4546 25803
rect -4500 25783 -4498 25803
rect -4404 25783 -4402 25803
rect -4308 25783 -4306 25803
rect -4260 25783 -4258 25803
rect -4164 25783 -4162 25803
rect -4020 25783 -4018 25803
rect -3876 25783 -3874 25803
rect -3732 25783 -3730 25803
rect -3588 25783 -3586 25803
rect -3564 25783 -3562 25803
rect -3516 25783 -3514 25803
rect -3492 25783 -3490 25803
rect -3468 25783 -3466 25803
rect -3420 25783 -3418 25803
rect -3324 25783 -3322 25803
rect -3228 25783 -3226 25803
rect -3156 25783 -3154 25803
rect -3132 25783 -3130 25803
rect -3060 25783 -3058 25803
rect -3012 25783 -3010 25803
rect -2964 25783 -2962 25803
rect -2916 25783 -2914 25803
rect -2892 25783 -2890 25803
rect -2868 25783 -2866 25803
rect -2820 25783 -2818 25803
rect -2796 25783 -2794 25803
rect -2772 25783 -2770 25803
rect -2676 25783 -2674 25803
rect -2580 25783 -2578 25803
rect -2364 25783 -2362 25803
rect -2268 25783 -2266 25803
rect -2244 25783 -2242 25803
rect -2172 25783 -2170 25803
rect -2148 25783 -2146 25803
rect -2076 25783 -2074 25803
rect -2052 25783 -2050 25803
rect -1980 25783 -1978 25803
rect -1884 25783 -1882 25803
rect -1836 25783 -1834 25803
rect -1572 25783 -1570 25803
rect -1476 25783 -1474 25803
rect -1380 25783 -1378 25803
rect -1356 25783 -1354 25803
rect -1308 25783 -1306 25803
rect -1260 25783 -1258 25803
rect -1140 25783 -1138 25803
rect -852 25783 -850 25803
rect -756 25783 -754 25803
rect -708 25783 -706 25803
rect -612 25783 -610 25803
rect -588 25783 -586 25803
rect -540 25783 -538 25803
rect -492 25783 -490 25803
rect -444 25783 -442 25803
rect -396 25783 -394 25803
rect -300 25783 -298 25803
rect -276 25783 -274 25803
rect -228 25783 -226 25803
rect -12 25783 -10 25803
rect 156 25783 158 25803
rect 204 25783 206 25803
rect 252 25783 254 25803
rect 348 25783 350 25803
rect 468 25783 470 25803
rect 492 25783 494 25803
rect 564 25783 566 25803
rect 588 25783 590 25803
rect 636 25783 638 25803
rect 660 25783 662 25803
rect 732 25783 734 25803
rect 1020 25783 1022 25803
rect 1092 25783 1094 25803
rect 1116 25783 1118 25803
rect 1212 25783 1214 25803
rect 1308 25783 1310 25803
rect 1332 25783 1334 25803
rect 1380 25783 1382 25803
rect 1428 25783 1430 25803
rect 1476 25783 1478 25803
rect 1548 25783 1550 25803
rect 1644 25783 1646 25803
rect 1692 25783 1694 25803
rect 1740 25783 1742 25803
rect 1788 25783 1790 25803
rect 2028 25783 2030 25803
rect 2076 25783 2078 25803
rect 2100 25783 2102 25803
rect 2124 25783 2126 25803
rect 2172 25783 2174 25803
rect 2185 25798 2188 25803
rect 2196 25798 2198 25803
rect 2195 25784 2198 25798
rect 2220 25783 2222 25803
rect 2268 25783 2270 25803
rect 2316 25783 2318 25803
rect 2364 25783 2366 25803
rect 2412 25783 2414 25803
rect 2460 25783 2462 25803
rect 2508 25783 2510 25803
rect 2580 25783 2582 25803
rect 2604 25783 2606 25803
rect 2676 25783 2678 25803
rect 2700 25783 2702 25803
rect 2748 25783 2750 25803
rect 2772 25783 2774 25803
rect 2796 25783 2798 25803
rect 2844 25783 2846 25803
rect 2868 25783 2870 25803
rect 2892 25783 2894 25803
rect 2940 25783 2942 25803
rect 3012 25783 3014 25803
rect 3108 25783 3110 25803
rect 3156 25783 3158 25803
rect 3252 25783 3254 25803
rect 3348 25783 3350 25803
rect 3396 25783 3398 25803
rect 3564 25783 3566 25803
rect 3612 25784 3614 25803
rect 3601 25783 3635 25784
rect 3636 25783 3638 25803
rect 3660 25783 3662 25803
rect 3708 25783 3710 25803
rect 3732 25783 3734 25803
rect 3804 25783 3806 25803
rect 3828 25783 3830 25803
rect 3924 25783 3926 25803
rect 4020 25783 4022 25803
rect 4044 25783 4046 25803
rect 4092 25783 4094 25803
rect 4116 25783 4118 25803
rect 4140 25783 4142 25803
rect 4188 25783 4190 25803
rect 4212 25783 4214 25803
rect 4236 25783 4238 25803
rect 4308 25783 4310 25803
rect 4332 25783 4334 25803
rect 4404 25783 4406 25803
rect 4500 25783 4502 25803
rect 4596 25783 4598 25803
rect 4692 25783 4694 25803
rect 4860 25783 4862 25803
rect 4956 25783 4958 25803
rect 4980 25783 4982 25803
rect 5004 25783 5006 25803
rect 5076 25783 5078 25803
rect 5100 25783 5102 25803
rect 5124 25783 5126 25803
rect 5172 25783 5174 25803
rect 5220 25783 5222 25803
rect 5268 25783 5270 25803
rect 5388 25783 5390 25803
rect 5484 25783 5486 25803
rect 5508 25783 5510 25803
rect 5532 25783 5534 25803
rect 5628 25783 5630 25803
rect 5652 25783 5654 25803
rect 5748 25783 5750 25803
rect 5796 25783 5798 25803
rect 5844 25783 5846 25803
rect 5892 25783 5894 25803
rect 6132 25783 6134 25803
rect 6180 25783 6182 25803
rect 6228 25783 6230 25803
rect 6252 25783 6254 25803
rect 6276 25783 6278 25803
rect 6324 25783 6326 25803
rect 6372 25783 6374 25803
rect 6492 25783 6494 25803
rect 6588 25783 6590 25803
rect 6612 25783 6614 25803
rect 6660 25783 6662 25803
rect 6684 25783 6686 25803
rect 6708 25783 6710 25803
rect 6780 25783 6782 25803
rect 6804 25783 6806 25803
rect 6828 25800 6830 25803
rect 6828 25783 6831 25800
rect 6900 25783 6902 25803
rect 6924 25783 6926 25803
rect 7020 25783 7022 25803
rect 7140 25783 7142 25803
rect 7236 25783 7238 25803
rect 7332 25783 7334 25803
rect 7380 25783 7382 25803
rect 7428 25783 7430 25803
rect 7452 25783 7454 25803
rect 7476 25783 7478 25803
rect 7524 25783 7526 25803
rect 7548 25783 7550 25803
rect 7572 25783 7574 25803
rect 7620 25783 7622 25803
rect 7644 25783 7646 25803
rect 7668 25783 7670 25803
rect 7740 25784 7742 25803
rect 7729 25783 7763 25784
rect 7788 25783 7790 25803
rect 7884 25783 7886 25803
rect 7956 25783 7958 25803
rect 7980 25783 7982 25803
rect 8028 25783 8030 25803
rect 8196 25783 8198 25803
rect 8244 25783 8246 25803
rect 8268 25783 8270 25803
rect 8292 25783 8294 25803
rect 8340 25783 8342 25803
rect 8364 25783 8366 25803
rect 8388 25783 8390 25803
rect 8436 25783 8438 25803
rect 8460 25784 8462 25803
rect 8449 25783 8483 25784
rect 8556 25783 8558 25803
rect 8604 25783 8606 25803
rect 8652 25783 8654 25803
rect 8700 25783 8702 25803
rect 8724 25783 8726 25803
rect 8748 25783 8750 25803
rect 8820 25783 8822 25803
rect 8844 25783 8846 25803
rect 8868 25783 8870 25803
rect 9516 25783 9518 25803
rect 9612 25783 9614 25803
rect 9660 25783 9662 25803
rect 9684 25783 9686 25803
rect 9708 25783 9710 25803
rect 9756 25783 9758 25803
rect 9780 25783 9782 25803
rect 9804 25783 9806 25803
rect 9852 25783 9854 25803
rect 9865 25798 9868 25803
rect 9876 25798 9878 25803
rect 9875 25784 9878 25798
rect 9900 25783 9902 25803
rect 9948 25783 9950 25803
rect 9972 25800 9974 25803
rect 9972 25783 9975 25800
rect 9996 25783 9998 25803
rect 10068 25783 10070 25803
rect 10092 25783 10094 25803
rect 10116 25783 10118 25803
rect 10164 25783 10166 25803
rect 10188 25783 10190 25803
rect 10212 25783 10214 25803
rect 10284 25783 10286 25803
rect 10308 25783 10310 25803
rect 10332 25783 10334 25803
rect 10380 25783 10382 25803
rect 10404 25783 10406 25803
rect 10428 25783 10430 25803
rect 10476 25783 10478 25803
rect 10500 25783 10502 25803
rect 10524 25783 10526 25803
rect 10572 25783 10574 25803
rect 10596 25783 10598 25803
rect 10620 25783 10622 25803
rect 10668 25783 10670 25803
rect 10692 25783 10694 25803
rect 10716 25783 10718 25803
rect 10788 25783 10790 25803
rect 10836 25783 10838 25803
rect 10956 25783 10958 25803
rect 11004 25783 11006 25803
rect 11052 25783 11054 25803
rect 11076 25783 11078 25803
rect 11100 25783 11102 25803
rect 11172 25783 11174 25803
rect 11220 25783 11222 25803
rect 11340 25783 11342 25803
rect 11436 25783 11438 25803
rect 11532 25783 11534 25803
rect 11580 25783 11582 25803
rect 11628 25783 11630 25803
rect 11676 25783 11678 25803
rect 11724 25783 11726 25803
rect 11772 25783 11774 25803
rect 11796 25783 11798 25803
rect 11892 25783 11894 25803
rect 11988 25783 11990 25803
rect 12060 25783 12062 25803
rect 12132 25783 12134 25803
rect 12228 25783 12230 25803
rect 12276 25783 12278 25803
rect 12324 25783 12326 25803
rect 12420 25783 12422 25803
rect 12444 25783 12446 25803
rect 12492 25783 12494 25803
rect 12516 25783 12518 25803
rect 12540 25783 12542 25803
rect 12588 25783 12590 25803
rect 12636 25783 12638 25803
rect 12732 25783 12734 25803
rect 12756 25783 12758 25803
rect 12804 25783 12806 25803
rect 12828 25783 12830 25803
rect 12852 25783 12854 25803
rect 12948 25783 12950 25803
rect 12951 25800 12965 25803
rect 12972 25803 27467 25807
rect 12972 25800 12989 25803
rect 12972 25783 12974 25800
rect 13044 25783 13046 25803
rect 13068 25783 13070 25803
rect 13116 25783 13118 25803
rect 13284 25783 13286 25803
rect 13332 25783 13334 25803
rect 13572 25783 13574 25803
rect 13644 25783 13646 25803
rect 13668 25783 13670 25803
rect 13764 25783 13766 25803
rect 13812 25783 13814 25803
rect 13860 25783 13862 25803
rect 13908 25783 13910 25803
rect 13956 25783 13958 25803
rect 14004 25783 14006 25803
rect 14100 25783 14102 25803
rect 14196 25783 14198 25803
rect 14292 25783 14294 25803
rect 15121 25798 15124 25803
rect 15132 25798 15134 25803
rect 15131 25784 15134 25798
rect 15180 25783 15182 25803
rect 15217 25798 15220 25803
rect 15228 25800 15230 25803
rect 15228 25798 15231 25800
rect 15227 25784 15231 25798
rect 15252 25783 15254 25803
rect 15265 25798 15268 25803
rect 15324 25800 15326 25803
rect 15396 25800 15398 25803
rect 15275 25784 15278 25798
rect 15313 25790 15317 25798
rect 15303 25784 15313 25790
rect 15276 25783 15278 25784
rect 15324 25783 15327 25800
rect 15396 25783 15399 25800
rect 15420 25783 15422 25803
rect 15492 25783 15494 25803
rect 15540 25783 15542 25803
rect 15636 25783 15638 25803
rect 15660 25783 15662 25803
rect 15708 25783 15710 25803
rect 15732 25783 15734 25803
rect 15756 25783 15758 25803
rect 15804 25783 15806 25803
rect 15828 25783 15830 25803
rect 15852 25783 15854 25803
rect 15900 25783 15902 25803
rect 15948 25783 15950 25803
rect 15996 25783 15998 25803
rect 16044 25783 16046 25803
rect 16164 25783 16166 25803
rect 16260 25783 16262 25803
rect 16308 25783 16310 25803
rect 16332 25783 16334 25803
rect 16356 25783 16358 25803
rect 16404 25783 16406 25803
rect 16452 25783 16454 25803
rect 16548 25783 16550 25803
rect 16572 25783 16574 25803
rect 16620 25783 16622 25803
rect 16668 25783 16670 25803
rect 16716 25783 16718 25803
rect 16764 25783 16766 25803
rect 16812 25783 16814 25803
rect 16884 25783 16886 25803
rect 16908 25783 16910 25803
rect 16980 25783 16982 25803
rect 17052 25783 17054 25803
rect 17196 25783 17198 25803
rect 17220 25783 17222 25803
rect 17292 25783 17294 25803
rect 17316 25783 17318 25803
rect 18084 25783 18086 25803
rect 18132 25783 18134 25803
rect 18228 25783 18230 25803
rect 18396 25783 18398 25803
rect 18492 25783 18494 25803
rect 18516 25783 18518 25803
rect 18564 25783 18566 25803
rect 18612 25783 18614 25803
rect 18660 25783 18662 25803
rect 18708 25783 18710 25803
rect 18756 25783 18758 25803
rect 18804 25783 18806 25803
rect 18852 25783 18854 25803
rect 18900 25783 18902 25803
rect 18996 25783 18998 25803
rect 19020 25783 19022 25803
rect 19092 25783 19094 25803
rect 19116 25783 19118 25803
rect 19140 25783 19142 25803
rect 19188 25783 19190 25803
rect 19236 25783 19238 25803
rect 19332 25783 19334 25803
rect 19476 25783 19478 25803
rect 19788 25783 19790 25803
rect 19836 25783 19838 25803
rect 19860 25783 19862 25803
rect 19884 25783 19886 25803
rect 19932 25783 19934 25803
rect 19956 25783 19958 25803
rect 19980 25783 19982 25803
rect 20028 25783 20030 25803
rect 20052 25783 20054 25803
rect 20076 25783 20078 25803
rect 20148 25783 20150 25803
rect 20172 25783 20174 25803
rect 20196 25783 20198 25803
rect 20268 25783 20270 25803
rect 20292 25783 20294 25803
rect 20388 25783 20390 25803
rect 20412 25783 20414 25803
rect 20508 25783 20510 25803
rect 20556 25783 20558 25803
rect 20604 25783 20606 25803
rect 20916 25783 20918 25803
rect 20964 25783 20966 25803
rect 21012 25783 21014 25803
rect 21060 25783 21062 25803
rect 21084 25784 21086 25803
rect 21073 25783 21107 25784
rect 21108 25783 21110 25803
rect 21204 25783 21206 25803
rect 21300 25783 21302 25803
rect 21324 25783 21326 25803
rect 21444 25783 21446 25803
rect 21468 25783 21470 25803
rect 21564 25783 21566 25803
rect 21612 25783 21614 25803
rect 21684 25783 21686 25803
rect 21708 25783 21710 25803
rect 21828 25783 21830 25803
rect 21924 25783 21926 25803
rect 22068 25783 22070 25803
rect 22188 25783 22190 25803
rect 22212 25783 22214 25803
rect 22884 25783 22886 25803
rect 22980 25783 22982 25803
rect 23076 25783 23078 25803
rect 23100 25783 23102 25803
rect 23124 25783 23126 25803
rect 23244 25783 23246 25803
rect 23340 25783 23342 25803
rect 23412 25783 23414 25803
rect 23508 25783 23510 25803
rect 23556 25783 23558 25803
rect 23652 25783 23654 25803
rect 23676 25783 23678 25803
rect 23724 25783 23726 25803
rect 23772 25783 23774 25803
rect 23820 25783 23822 25803
rect 23916 25783 23918 25803
rect 23953 25783 24011 25784
rect 24012 25783 24014 25803
rect 24084 25783 24086 25803
rect 24396 25783 24398 25803
rect 24492 25783 24494 25803
rect 24516 25783 24518 25803
rect 24588 25783 24590 25803
rect 24612 25783 24614 25803
rect 24684 25783 24686 25803
rect 24732 25783 24734 25803
rect 24756 25783 24758 25803
rect 24780 25783 24782 25803
rect 24852 25783 24854 25803
rect 24876 25783 24878 25803
rect 24972 25783 24974 25803
rect 24996 25783 24998 25803
rect 25068 25783 25070 25803
rect 25164 25783 25166 25803
rect 25260 25783 25262 25803
rect 25284 25783 25286 25803
rect 25356 25783 25358 25803
rect 25380 25783 25382 25803
rect 25404 25783 25406 25803
rect 25500 25783 25502 25803
rect 25596 25783 25598 25803
rect 27036 25783 27038 25803
rect 27108 25783 27110 25803
rect 27324 25783 27326 25803
rect 27396 25783 27398 25803
rect 27420 25784 27422 25803
rect 27409 25783 27443 25784
rect -16617 25779 15365 25783
rect -16617 25776 -16603 25779
rect -16524 25776 -16522 25779
rect -16524 25760 -16521 25776
rect -16535 25759 -16501 25760
rect -16404 25759 -16402 25779
rect -16356 25759 -16354 25779
rect -16308 25759 -16306 25779
rect -16284 25759 -16282 25779
rect -16260 25759 -16258 25779
rect -15324 25759 -15322 25779
rect -15108 25759 -15106 25779
rect -14772 25759 -14770 25779
rect -14519 25759 -14485 25760
rect -14436 25759 -14434 25779
rect -14340 25759 -14338 25779
rect -13980 25759 -13978 25779
rect -13932 25759 -13930 25779
rect -13884 25759 -13882 25779
rect -13788 25759 -13786 25779
rect -13572 25759 -13570 25779
rect -13356 25759 -13354 25779
rect -13068 25759 -13066 25779
rect -12780 25759 -12778 25779
rect -12756 25759 -12754 25779
rect -12660 25759 -12658 25779
rect -12564 25759 -12562 25779
rect -12492 25759 -12490 25779
rect -12396 25759 -12394 25779
rect -12348 25759 -12346 25779
rect -12252 25759 -12250 25779
rect -12156 25759 -12154 25779
rect -12060 25759 -12058 25779
rect -11844 25759 -11842 25779
rect -11721 25776 -11707 25779
rect -11676 25759 -11674 25779
rect -11556 25759 -11554 25779
rect -11508 25759 -11506 25779
rect -11436 25759 -11434 25779
rect -11412 25759 -11410 25779
rect -11340 25759 -11338 25779
rect -11196 25759 -11194 25779
rect -11124 25759 -11122 25779
rect -11100 25759 -11098 25779
rect -11028 25759 -11026 25779
rect -10740 25759 -10738 25779
rect -10668 25759 -10666 25779
rect -10644 25759 -10642 25779
rect -9996 25759 -9994 25779
rect -9828 25759 -9826 25779
rect -9732 25759 -9730 25779
rect -9612 25776 -9610 25779
rect -9612 25759 -9609 25776
rect -9516 25759 -9514 25779
rect -9468 25759 -9466 25779
rect -9420 25759 -9418 25779
rect -9252 25759 -9250 25779
rect -8604 25759 -8602 25779
rect -8484 25759 -8482 25779
rect -8436 25759 -8434 25779
rect -8388 25759 -8386 25779
rect -8364 25759 -8362 25779
rect -8340 25759 -8338 25779
rect -8268 25759 -8266 25779
rect -8100 25759 -8098 25779
rect -8052 25759 -8050 25779
rect -7932 25759 -7930 25779
rect -7692 25759 -7690 25779
rect -7620 25759 -7618 25779
rect -7524 25759 -7522 25779
rect -7356 25759 -7354 25779
rect -7308 25759 -7306 25779
rect -7212 25759 -7210 25779
rect -7116 25759 -7114 25779
rect -7068 25759 -7066 25779
rect -6972 25759 -6970 25779
rect -6948 25759 -6946 25779
rect -6876 25759 -6874 25779
rect -6852 25759 -6850 25779
rect -6780 25759 -6778 25779
rect -6756 25759 -6754 25779
rect -6660 25759 -6658 25779
rect -6612 25759 -6610 25779
rect -6516 25759 -6514 25779
rect -6420 25759 -6418 25779
rect -6372 25759 -6370 25779
rect -6324 25759 -6322 25779
rect -6156 25759 -6154 25779
rect -6060 25759 -6058 25779
rect -6036 25759 -6034 25779
rect -5892 25759 -5890 25779
rect -5652 25759 -5650 25779
rect -5268 25759 -5266 25779
rect -5196 25759 -5194 25779
rect -5172 25759 -5170 25779
rect -5100 25759 -5098 25779
rect -5076 25759 -5074 25779
rect -4980 25759 -4978 25779
rect -4956 25759 -4954 25779
rect -4860 25759 -4858 25779
rect -4644 25759 -4642 25779
rect -4548 25759 -4546 25779
rect -4500 25759 -4498 25779
rect -4404 25759 -4402 25779
rect -4308 25759 -4306 25779
rect -4260 25759 -4258 25779
rect -4164 25759 -4162 25779
rect -4020 25759 -4018 25779
rect -3876 25759 -3874 25779
rect -3732 25759 -3730 25779
rect -3588 25759 -3586 25779
rect -3564 25759 -3562 25779
rect -3516 25759 -3514 25779
rect -3492 25759 -3490 25779
rect -3468 25759 -3466 25779
rect -3420 25759 -3418 25779
rect -3324 25759 -3322 25779
rect -3228 25759 -3226 25779
rect -3156 25760 -3154 25779
rect -3167 25759 -3133 25760
rect -3132 25759 -3130 25779
rect -3060 25759 -3058 25779
rect -3012 25759 -3010 25779
rect -2964 25759 -2962 25779
rect -2916 25759 -2914 25779
rect -2892 25759 -2890 25779
rect -2868 25759 -2866 25779
rect -2820 25759 -2818 25779
rect -2796 25759 -2794 25779
rect -2772 25759 -2770 25779
rect -2676 25759 -2674 25779
rect -2580 25759 -2578 25779
rect -2364 25759 -2362 25779
rect -2268 25759 -2266 25779
rect -2244 25759 -2242 25779
rect -2172 25759 -2170 25779
rect -2148 25759 -2146 25779
rect -2076 25759 -2074 25779
rect -2052 25759 -2050 25779
rect -1980 25759 -1978 25779
rect -1884 25759 -1882 25779
rect -1836 25760 -1834 25779
rect -1847 25759 -1813 25760
rect -1572 25759 -1570 25779
rect -1476 25759 -1474 25779
rect -1380 25759 -1378 25779
rect -1356 25759 -1354 25779
rect -1308 25759 -1306 25779
rect -1260 25759 -1258 25779
rect -1140 25759 -1138 25779
rect -852 25759 -850 25779
rect -756 25759 -754 25779
rect -708 25759 -706 25779
rect -612 25759 -610 25779
rect -588 25759 -586 25779
rect -540 25759 -538 25779
rect -492 25759 -490 25779
rect -444 25759 -442 25779
rect -396 25759 -394 25779
rect -300 25759 -298 25779
rect -276 25759 -274 25779
rect -228 25759 -226 25779
rect -12 25759 -10 25779
rect 156 25759 158 25779
rect 204 25759 206 25779
rect 252 25759 254 25779
rect 348 25759 350 25779
rect 468 25759 470 25779
rect 492 25759 494 25779
rect 564 25759 566 25779
rect 588 25759 590 25779
rect 636 25759 638 25779
rect 660 25759 662 25779
rect 732 25759 734 25779
rect 1020 25759 1022 25779
rect 1092 25759 1094 25779
rect 1116 25759 1118 25779
rect 1212 25759 1214 25779
rect 1308 25759 1310 25779
rect 1332 25759 1334 25779
rect 1380 25759 1382 25779
rect 1428 25759 1430 25779
rect 1476 25759 1478 25779
rect 1548 25759 1550 25779
rect 1644 25759 1646 25779
rect 1692 25759 1694 25779
rect 1740 25759 1742 25779
rect 1788 25759 1790 25779
rect 2028 25759 2030 25779
rect 2076 25759 2078 25779
rect 2100 25759 2102 25779
rect 2124 25759 2126 25779
rect 2172 25759 2174 25779
rect 2220 25759 2222 25779
rect 2268 25759 2270 25779
rect 2271 25776 2285 25779
rect 2316 25759 2318 25779
rect 2364 25759 2366 25779
rect 2412 25759 2414 25779
rect 2460 25759 2462 25779
rect 2508 25759 2510 25779
rect 2580 25759 2582 25779
rect 2604 25759 2606 25779
rect 2676 25759 2678 25779
rect 2700 25759 2702 25779
rect 2748 25759 2750 25779
rect 2772 25759 2774 25779
rect 2796 25759 2798 25779
rect 2844 25759 2846 25779
rect 2868 25759 2870 25779
rect 2892 25759 2894 25779
rect 2940 25759 2942 25779
rect 3012 25759 3014 25779
rect 3108 25759 3110 25779
rect 3156 25759 3158 25779
rect 3252 25759 3254 25779
rect 3348 25759 3350 25779
rect 3396 25759 3398 25779
rect 3564 25759 3566 25779
rect 3601 25774 3604 25779
rect 3612 25774 3614 25779
rect 3611 25760 3614 25774
rect 3636 25759 3638 25779
rect 3660 25759 3662 25779
rect 3708 25776 3710 25779
rect 3708 25759 3711 25776
rect 3732 25759 3734 25779
rect 3804 25760 3806 25779
rect 3769 25759 3827 25760
rect 3828 25759 3830 25779
rect 3924 25759 3926 25779
rect 4020 25759 4022 25779
rect 4044 25759 4046 25779
rect 4092 25759 4094 25779
rect 4116 25759 4118 25779
rect 4140 25759 4142 25779
rect 4188 25759 4190 25779
rect 4212 25759 4214 25779
rect 4236 25759 4238 25779
rect 4308 25759 4310 25779
rect 4332 25759 4334 25779
rect 4404 25759 4406 25779
rect 4500 25759 4502 25779
rect 4596 25759 4598 25779
rect 4692 25759 4694 25779
rect 4860 25759 4862 25779
rect 4956 25759 4958 25779
rect 4980 25759 4982 25779
rect 5004 25759 5006 25779
rect 5076 25759 5078 25779
rect 5100 25759 5102 25779
rect 5124 25759 5126 25779
rect 5172 25759 5174 25779
rect 5220 25759 5222 25779
rect 5268 25759 5270 25779
rect 5388 25759 5390 25779
rect 5484 25759 5486 25779
rect 5508 25759 5510 25779
rect 5532 25759 5534 25779
rect 5628 25759 5630 25779
rect 5652 25759 5654 25779
rect 5748 25759 5750 25779
rect 5796 25759 5798 25779
rect 5844 25759 5846 25779
rect 5892 25759 5894 25779
rect 6132 25759 6134 25779
rect 6180 25759 6182 25779
rect 6228 25759 6230 25779
rect 6252 25759 6254 25779
rect 6276 25759 6278 25779
rect 6324 25759 6326 25779
rect 6372 25759 6374 25779
rect 6492 25759 6494 25779
rect 6588 25759 6590 25779
rect 6612 25759 6614 25779
rect 6660 25759 6662 25779
rect 6684 25759 6686 25779
rect 6708 25759 6710 25779
rect 6780 25759 6782 25779
rect 6804 25759 6806 25779
rect 6807 25776 6821 25779
rect 6828 25776 6831 25779
rect 6900 25759 6902 25779
rect 6924 25759 6926 25779
rect 7020 25759 7022 25779
rect 7140 25759 7142 25779
rect 7236 25759 7238 25779
rect 7332 25759 7334 25779
rect 7380 25759 7382 25779
rect 7428 25759 7430 25779
rect 7452 25759 7454 25779
rect 7476 25759 7478 25779
rect 7524 25759 7526 25779
rect 7548 25759 7550 25779
rect 7572 25759 7574 25779
rect 7620 25759 7622 25779
rect 7644 25759 7646 25779
rect 7668 25759 7670 25779
rect 7729 25774 7732 25779
rect 7740 25774 7742 25779
rect 7739 25760 7742 25774
rect 7788 25759 7790 25779
rect 7884 25759 7886 25779
rect 7956 25759 7958 25779
rect 7980 25759 7982 25779
rect 8028 25759 8030 25779
rect 8196 25759 8198 25779
rect 8244 25759 8246 25779
rect 8268 25759 8270 25779
rect 8292 25759 8294 25779
rect 8340 25759 8342 25779
rect 8364 25759 8366 25779
rect 8388 25759 8390 25779
rect 8436 25759 8438 25779
rect 8449 25774 8452 25779
rect 8460 25774 8462 25779
rect 8459 25760 8462 25774
rect 8556 25776 8558 25779
rect 8556 25759 8559 25776
rect 8604 25759 8606 25779
rect 8652 25759 8654 25779
rect 8700 25759 8702 25779
rect 8724 25759 8726 25779
rect 8748 25759 8750 25779
rect 8820 25759 8822 25779
rect 8844 25759 8846 25779
rect 8868 25759 8870 25779
rect 9516 25759 9518 25779
rect 9612 25759 9614 25779
rect 9660 25759 9662 25779
rect 9684 25759 9686 25779
rect 9708 25759 9710 25779
rect 9756 25759 9758 25779
rect 9780 25759 9782 25779
rect 9804 25759 9806 25779
rect 9852 25759 9854 25779
rect 9900 25759 9902 25779
rect 9948 25759 9950 25779
rect 9951 25776 9965 25779
rect 9972 25776 9975 25779
rect 9996 25759 9998 25779
rect 10068 25759 10070 25779
rect 10092 25759 10094 25779
rect 10116 25759 10118 25779
rect 10164 25759 10166 25779
rect 10188 25759 10190 25779
rect 10212 25759 10214 25779
rect 10284 25759 10286 25779
rect 10308 25759 10310 25779
rect 10332 25759 10334 25779
rect 10380 25759 10382 25779
rect 10404 25759 10406 25779
rect 10428 25759 10430 25779
rect 10476 25759 10478 25779
rect 10500 25759 10502 25779
rect 10524 25759 10526 25779
rect 10572 25759 10574 25779
rect 10596 25759 10598 25779
rect 10620 25759 10622 25779
rect 10668 25759 10670 25779
rect 10692 25759 10694 25779
rect 10716 25759 10718 25779
rect 10788 25759 10790 25779
rect 10836 25759 10838 25779
rect 10956 25759 10958 25779
rect 11004 25759 11006 25779
rect 11052 25759 11054 25779
rect 11076 25759 11078 25779
rect 11100 25759 11102 25779
rect 11172 25759 11174 25779
rect 11220 25759 11222 25779
rect 11340 25759 11342 25779
rect 11436 25759 11438 25779
rect 11532 25759 11534 25779
rect 11580 25759 11582 25779
rect 11628 25759 11630 25779
rect 11676 25759 11678 25779
rect 11724 25759 11726 25779
rect 11772 25759 11774 25779
rect 11796 25759 11798 25779
rect 11892 25759 11894 25779
rect 11988 25759 11990 25779
rect 12060 25759 12062 25779
rect 12132 25759 12134 25779
rect 12228 25759 12230 25779
rect 12276 25759 12278 25779
rect 12324 25759 12326 25779
rect 12420 25759 12422 25779
rect 12444 25759 12446 25779
rect 12492 25759 12494 25779
rect 12516 25759 12518 25779
rect 12540 25759 12542 25779
rect 12588 25759 12590 25779
rect 12636 25759 12638 25779
rect 12732 25759 12734 25779
rect 12756 25759 12758 25779
rect 12804 25759 12806 25779
rect 12828 25759 12830 25779
rect 12852 25759 12854 25779
rect 12948 25759 12950 25779
rect 12972 25759 12974 25779
rect 13044 25759 13046 25779
rect 13068 25759 13070 25779
rect 13116 25759 13118 25779
rect 13284 25759 13286 25779
rect 13332 25759 13334 25779
rect 13572 25759 13574 25779
rect 13644 25759 13646 25779
rect 13668 25759 13670 25779
rect 13764 25759 13766 25779
rect 13812 25759 13814 25779
rect 13860 25759 13862 25779
rect 13908 25759 13910 25779
rect 13956 25759 13958 25779
rect 14004 25759 14006 25779
rect 14100 25759 14102 25779
rect 14196 25759 14198 25779
rect 14292 25759 14294 25779
rect 15180 25759 15182 25779
rect 15207 25776 15221 25779
rect 15252 25759 15254 25779
rect 15276 25759 15278 25779
rect 15303 25776 15317 25779
rect 15324 25776 15327 25779
rect 15351 25776 15365 25779
rect 15375 25779 27443 25783
rect 15375 25776 15389 25779
rect 15396 25776 15399 25779
rect 15420 25759 15422 25779
rect 15492 25759 15494 25779
rect 15540 25759 15542 25779
rect 15636 25759 15638 25779
rect 15660 25759 15662 25779
rect 15708 25759 15710 25779
rect 15732 25759 15734 25779
rect 15756 25759 15758 25779
rect 15804 25759 15806 25779
rect 15828 25759 15830 25779
rect 15852 25759 15854 25779
rect 15900 25759 15902 25779
rect 15948 25759 15950 25779
rect 15996 25759 15998 25779
rect 16044 25759 16046 25779
rect 16164 25759 16166 25779
rect 16260 25759 16262 25779
rect 16308 25759 16310 25779
rect 16332 25759 16334 25779
rect 16356 25759 16358 25779
rect 16404 25759 16406 25779
rect 16452 25759 16454 25779
rect 16548 25759 16550 25779
rect 16572 25759 16574 25779
rect 16620 25759 16622 25779
rect 16668 25759 16670 25779
rect 16716 25759 16718 25779
rect 16764 25759 16766 25779
rect 16812 25759 16814 25779
rect 16884 25759 16886 25779
rect 16908 25759 16910 25779
rect 16980 25759 16982 25779
rect 17052 25759 17054 25779
rect 17196 25759 17198 25779
rect 17220 25759 17222 25779
rect 17292 25759 17294 25779
rect 17316 25759 17318 25779
rect 18084 25759 18086 25779
rect 18132 25759 18134 25779
rect 18228 25759 18230 25779
rect 18396 25759 18398 25779
rect 18492 25759 18494 25779
rect 18516 25759 18518 25779
rect 18564 25759 18566 25779
rect 18612 25759 18614 25779
rect 18660 25759 18662 25779
rect 18708 25759 18710 25779
rect 18756 25759 18758 25779
rect 18804 25759 18806 25779
rect 18852 25759 18854 25779
rect 18900 25759 18902 25779
rect 18996 25759 18998 25779
rect 19020 25759 19022 25779
rect 19092 25759 19094 25779
rect 19116 25759 19118 25779
rect 19140 25759 19142 25779
rect 19188 25759 19190 25779
rect 19236 25759 19238 25779
rect 19332 25759 19334 25779
rect 19476 25759 19478 25779
rect 19788 25759 19790 25779
rect 19836 25759 19838 25779
rect 19860 25759 19862 25779
rect 19884 25759 19886 25779
rect 19932 25759 19934 25779
rect 19956 25759 19958 25779
rect 19980 25759 19982 25779
rect 20028 25759 20030 25779
rect 20052 25759 20054 25779
rect 20076 25759 20078 25779
rect 20148 25759 20150 25779
rect 20172 25759 20174 25779
rect 20196 25759 20198 25779
rect 20268 25759 20270 25779
rect 20292 25759 20294 25779
rect 20388 25759 20390 25779
rect 20412 25759 20414 25779
rect 20508 25759 20510 25779
rect 20556 25759 20558 25779
rect 20604 25759 20606 25779
rect 20916 25759 20918 25779
rect 20964 25759 20966 25779
rect 21012 25759 21014 25779
rect 21060 25759 21062 25779
rect 21073 25774 21076 25779
rect 21084 25774 21086 25779
rect 21083 25760 21086 25774
rect 21108 25759 21110 25779
rect 21204 25759 21206 25779
rect 21300 25759 21302 25779
rect 21324 25759 21326 25779
rect 21444 25759 21446 25779
rect 21468 25759 21470 25779
rect 21564 25759 21566 25779
rect 21612 25759 21614 25779
rect 21684 25759 21686 25779
rect 21708 25759 21710 25779
rect 21828 25759 21830 25779
rect 21924 25759 21926 25779
rect 22068 25759 22070 25779
rect 22188 25759 22190 25779
rect 22212 25759 22214 25779
rect 22884 25759 22886 25779
rect 22980 25759 22982 25779
rect 23076 25759 23078 25779
rect 23100 25759 23102 25779
rect 23124 25759 23126 25779
rect 23244 25759 23246 25779
rect 23340 25759 23342 25779
rect 23412 25759 23414 25779
rect 23508 25759 23510 25779
rect 23556 25759 23558 25779
rect 23652 25759 23654 25779
rect 23676 25759 23678 25779
rect 23724 25759 23726 25779
rect 23772 25759 23774 25779
rect 23820 25759 23822 25779
rect 23916 25759 23918 25779
rect 24012 25759 24014 25779
rect 24084 25776 24086 25779
rect 24084 25759 24087 25776
rect 24396 25759 24398 25779
rect 24492 25759 24494 25779
rect 24516 25759 24518 25779
rect 24588 25759 24590 25779
rect 24612 25759 24614 25779
rect 24684 25759 24686 25779
rect 24732 25759 24734 25779
rect 24756 25759 24758 25779
rect 24780 25759 24782 25779
rect 24852 25759 24854 25779
rect 24876 25759 24878 25779
rect 24972 25759 24974 25779
rect 24996 25759 24998 25779
rect 25068 25759 25070 25779
rect 25164 25759 25166 25779
rect 25260 25759 25262 25779
rect 25284 25759 25286 25779
rect 25356 25759 25358 25779
rect 25380 25759 25382 25779
rect 25404 25759 25406 25779
rect 25500 25759 25502 25779
rect 25596 25759 25598 25779
rect 27036 25759 27038 25779
rect 27108 25759 27110 25779
rect 27324 25759 27326 25779
rect 27396 25760 27398 25779
rect 27409 25774 27412 25779
rect 27420 25774 27422 25779
rect 27419 25760 27422 25774
rect 27385 25759 27419 25760
rect -16535 25755 24053 25759
rect -16535 25752 -16531 25755
rect -16524 25752 -16521 25755
rect -16404 25735 -16402 25755
rect -16356 25735 -16354 25755
rect -16308 25735 -16306 25755
rect -16284 25735 -16282 25755
rect -16260 25735 -16258 25755
rect -16079 25735 -16021 25736
rect -15324 25735 -15322 25755
rect -15108 25735 -15106 25755
rect -14772 25735 -14770 25755
rect -14436 25735 -14434 25755
rect -14340 25735 -14338 25755
rect -14193 25752 -14179 25755
rect -13980 25736 -13978 25755
rect -14015 25735 -13957 25736
rect -13932 25735 -13930 25755
rect -13884 25735 -13882 25755
rect -13788 25735 -13786 25755
rect -13572 25735 -13570 25755
rect -13356 25735 -13354 25755
rect -13068 25735 -13066 25755
rect -12780 25735 -12778 25755
rect -12756 25735 -12754 25755
rect -12660 25735 -12658 25755
rect -12564 25735 -12562 25755
rect -12492 25735 -12490 25755
rect -12396 25735 -12394 25755
rect -12348 25735 -12346 25755
rect -12252 25735 -12250 25755
rect -12156 25735 -12154 25755
rect -12119 25735 -12085 25736
rect -12060 25735 -12058 25755
rect -11844 25735 -11842 25755
rect -11676 25735 -11674 25755
rect -11556 25735 -11554 25755
rect -11508 25735 -11506 25755
rect -11436 25735 -11434 25755
rect -11412 25735 -11410 25755
rect -11340 25735 -11338 25755
rect -11196 25735 -11194 25755
rect -11124 25735 -11122 25755
rect -11100 25735 -11098 25755
rect -11028 25735 -11026 25755
rect -10740 25735 -10738 25755
rect -10668 25735 -10666 25755
rect -10644 25735 -10642 25755
rect -9996 25735 -9994 25755
rect -9828 25735 -9826 25755
rect -9732 25735 -9730 25755
rect -9633 25752 -9619 25755
rect -9612 25752 -9609 25755
rect -9516 25735 -9514 25755
rect -9468 25735 -9466 25755
rect -9420 25735 -9418 25755
rect -9252 25736 -9250 25755
rect -9287 25735 -9229 25736
rect -8604 25735 -8602 25755
rect -8484 25735 -8482 25755
rect -8436 25735 -8434 25755
rect -8388 25735 -8386 25755
rect -8364 25735 -8362 25755
rect -8340 25735 -8338 25755
rect -8268 25735 -8266 25755
rect -8100 25735 -8098 25755
rect -8052 25735 -8050 25755
rect -7932 25735 -7930 25755
rect -7692 25735 -7690 25755
rect -7620 25735 -7618 25755
rect -7524 25735 -7522 25755
rect -7356 25735 -7354 25755
rect -7308 25735 -7306 25755
rect -7212 25735 -7210 25755
rect -7116 25735 -7114 25755
rect -7068 25735 -7066 25755
rect -6972 25735 -6970 25755
rect -6948 25735 -6946 25755
rect -6876 25735 -6874 25755
rect -6852 25735 -6850 25755
rect -6780 25735 -6778 25755
rect -6756 25735 -6754 25755
rect -6660 25735 -6658 25755
rect -6612 25735 -6610 25755
rect -6516 25735 -6514 25755
rect -6420 25736 -6418 25755
rect -6455 25735 -6397 25736
rect -6372 25735 -6370 25755
rect -6324 25735 -6322 25755
rect -6156 25735 -6154 25755
rect -6060 25735 -6058 25755
rect -6036 25735 -6034 25755
rect -5892 25735 -5890 25755
rect -5652 25735 -5650 25755
rect -5268 25735 -5266 25755
rect -5196 25735 -5194 25755
rect -5172 25735 -5170 25755
rect -5100 25735 -5098 25755
rect -5076 25735 -5074 25755
rect -4980 25735 -4978 25755
rect -4956 25735 -4954 25755
rect -4860 25735 -4858 25755
rect -4644 25735 -4642 25755
rect -4548 25735 -4546 25755
rect -4500 25735 -4498 25755
rect -4404 25735 -4402 25755
rect -4308 25735 -4306 25755
rect -4260 25735 -4258 25755
rect -4164 25735 -4162 25755
rect -4020 25735 -4018 25755
rect -3876 25735 -3874 25755
rect -3732 25735 -3730 25755
rect -3588 25735 -3586 25755
rect -3564 25735 -3562 25755
rect -3516 25735 -3514 25755
rect -3492 25735 -3490 25755
rect -3468 25735 -3466 25755
rect -3420 25735 -3418 25755
rect -3324 25735 -3322 25755
rect -3228 25735 -3226 25755
rect -3167 25750 -3164 25755
rect -3156 25750 -3154 25755
rect -3157 25736 -3154 25750
rect -3132 25735 -3130 25755
rect -3060 25752 -3058 25755
rect -3060 25735 -3057 25752
rect -3012 25735 -3010 25755
rect -2964 25735 -2962 25755
rect -2916 25735 -2914 25755
rect -2892 25735 -2890 25755
rect -2868 25735 -2866 25755
rect -2820 25735 -2818 25755
rect -2796 25735 -2794 25755
rect -2772 25735 -2770 25755
rect -2676 25735 -2674 25755
rect -2580 25735 -2578 25755
rect -2364 25735 -2362 25755
rect -2327 25735 -2269 25736
rect -2268 25735 -2266 25755
rect -2244 25735 -2242 25755
rect -2172 25735 -2170 25755
rect -2148 25735 -2146 25755
rect -2076 25735 -2074 25755
rect -2052 25735 -2050 25755
rect -1980 25735 -1978 25755
rect -1884 25735 -1882 25755
rect -1847 25750 -1844 25755
rect -1836 25750 -1834 25755
rect -1837 25736 -1834 25750
rect -1572 25735 -1570 25755
rect -1476 25735 -1474 25755
rect -1380 25735 -1378 25755
rect -1356 25735 -1354 25755
rect -1308 25735 -1306 25755
rect -1260 25735 -1258 25755
rect -1140 25735 -1138 25755
rect -1031 25735 -997 25736
rect -852 25735 -850 25755
rect -756 25735 -754 25755
rect -708 25735 -706 25755
rect -612 25735 -610 25755
rect -588 25735 -586 25755
rect -540 25735 -538 25755
rect -492 25735 -490 25755
rect -444 25735 -442 25755
rect -396 25735 -394 25755
rect -300 25735 -298 25755
rect -276 25735 -274 25755
rect -228 25735 -226 25755
rect -12 25735 -10 25755
rect 156 25735 158 25755
rect 204 25735 206 25755
rect 252 25735 254 25755
rect 348 25735 350 25755
rect 468 25735 470 25755
rect 492 25735 494 25755
rect 564 25735 566 25755
rect 588 25735 590 25755
rect 636 25735 638 25755
rect 660 25735 662 25755
rect 732 25735 734 25755
rect 1020 25736 1022 25755
rect 1009 25735 1043 25736
rect 1092 25735 1094 25755
rect 1116 25736 1118 25755
rect 1105 25735 1139 25736
rect 1212 25735 1214 25755
rect 1308 25735 1310 25755
rect 1332 25735 1334 25755
rect 1380 25735 1382 25755
rect 1428 25735 1430 25755
rect 1441 25735 1475 25736
rect 1476 25735 1478 25755
rect 1548 25735 1550 25755
rect 1644 25735 1646 25755
rect 1692 25735 1694 25755
rect 1740 25735 1742 25755
rect 1788 25735 1790 25755
rect 2028 25735 2030 25755
rect 2076 25735 2078 25755
rect 2100 25735 2102 25755
rect 2124 25735 2126 25755
rect 2172 25735 2174 25755
rect 2220 25735 2222 25755
rect 2268 25735 2270 25755
rect 2316 25735 2318 25755
rect 2364 25735 2366 25755
rect 2412 25735 2414 25755
rect 2460 25735 2462 25755
rect 2508 25735 2510 25755
rect 2580 25735 2582 25755
rect 2604 25735 2606 25755
rect 2676 25735 2678 25755
rect 2700 25735 2702 25755
rect 2748 25735 2750 25755
rect 2772 25735 2774 25755
rect 2796 25735 2798 25755
rect 2844 25735 2846 25755
rect 2868 25735 2870 25755
rect 2892 25735 2894 25755
rect 2940 25735 2942 25755
rect 3012 25735 3014 25755
rect 3108 25735 3110 25755
rect 3156 25735 3158 25755
rect 3252 25735 3254 25755
rect 3348 25735 3350 25755
rect 3396 25735 3398 25755
rect 3564 25735 3566 25755
rect 3636 25735 3638 25755
rect 3660 25735 3662 25755
rect 3687 25752 3701 25755
rect 3708 25752 3711 25755
rect 3732 25735 3734 25755
rect 3793 25750 3796 25755
rect 3804 25750 3806 25755
rect 3803 25736 3806 25750
rect 3828 25735 3830 25755
rect 3924 25735 3926 25755
rect 4020 25735 4022 25755
rect 4044 25735 4046 25755
rect 4092 25735 4094 25755
rect 4116 25735 4118 25755
rect 4140 25735 4142 25755
rect 4188 25735 4190 25755
rect 4212 25735 4214 25755
rect 4236 25735 4238 25755
rect 4308 25735 4310 25755
rect 4332 25735 4334 25755
rect 4404 25735 4406 25755
rect 4500 25735 4502 25755
rect 4596 25735 4598 25755
rect 4692 25735 4694 25755
rect 4860 25735 4862 25755
rect 4956 25735 4958 25755
rect 4980 25735 4982 25755
rect 5004 25735 5006 25755
rect 5076 25736 5078 25755
rect 5041 25735 5099 25736
rect 5100 25735 5102 25755
rect 5124 25735 5126 25755
rect 5172 25735 5174 25755
rect 5220 25735 5222 25755
rect 5268 25735 5270 25755
rect 5388 25735 5390 25755
rect 5484 25735 5486 25755
rect 5508 25735 5510 25755
rect 5532 25735 5534 25755
rect 5628 25735 5630 25755
rect 5652 25735 5654 25755
rect 5748 25735 5750 25755
rect 5796 25735 5798 25755
rect 5844 25735 5846 25755
rect 5892 25735 5894 25755
rect 6132 25735 6134 25755
rect 6180 25735 6182 25755
rect 6228 25735 6230 25755
rect 6252 25735 6254 25755
rect 6276 25735 6278 25755
rect 6324 25735 6326 25755
rect 6372 25735 6374 25755
rect 6492 25735 6494 25755
rect 6588 25735 6590 25755
rect 6612 25735 6614 25755
rect 6660 25735 6662 25755
rect 6684 25735 6686 25755
rect 6708 25735 6710 25755
rect 6780 25735 6782 25755
rect 6804 25735 6806 25755
rect 6900 25735 6902 25755
rect 6924 25735 6926 25755
rect 7020 25735 7022 25755
rect 7140 25735 7142 25755
rect 7236 25735 7238 25755
rect 7332 25735 7334 25755
rect 7380 25735 7382 25755
rect 7428 25735 7430 25755
rect 7452 25735 7454 25755
rect 7476 25735 7478 25755
rect 7524 25735 7526 25755
rect 7548 25735 7550 25755
rect 7572 25735 7574 25755
rect 7620 25735 7622 25755
rect 7644 25735 7646 25755
rect 7668 25735 7670 25755
rect 7788 25735 7790 25755
rect 7815 25752 7829 25755
rect 7884 25735 7886 25755
rect 7956 25735 7958 25755
rect 7980 25735 7982 25755
rect 8028 25735 8030 25755
rect 8196 25735 8198 25755
rect 8244 25735 8246 25755
rect 8268 25735 8270 25755
rect 8292 25735 8294 25755
rect 8340 25735 8342 25755
rect 8364 25735 8366 25755
rect 8388 25735 8390 25755
rect 8436 25735 8438 25755
rect 8535 25752 8549 25755
rect 8556 25752 8559 25755
rect 8604 25735 8606 25755
rect 8652 25735 8654 25755
rect 8700 25735 8702 25755
rect 8724 25735 8726 25755
rect 8748 25735 8750 25755
rect 8820 25735 8822 25755
rect 8844 25735 8846 25755
rect 8868 25735 8870 25755
rect 9516 25735 9518 25755
rect 9612 25735 9614 25755
rect 9660 25735 9662 25755
rect 9684 25735 9686 25755
rect 9708 25735 9710 25755
rect 9756 25735 9758 25755
rect 9780 25735 9782 25755
rect 9804 25735 9806 25755
rect 9852 25735 9854 25755
rect 9900 25735 9902 25755
rect 9948 25735 9950 25755
rect 9996 25735 9998 25755
rect 10068 25735 10070 25755
rect 10092 25735 10094 25755
rect 10116 25735 10118 25755
rect 10164 25735 10166 25755
rect 10188 25735 10190 25755
rect 10212 25735 10214 25755
rect 10284 25735 10286 25755
rect 10308 25735 10310 25755
rect 10332 25735 10334 25755
rect 10380 25735 10382 25755
rect 10404 25735 10406 25755
rect 10428 25735 10430 25755
rect 10476 25735 10478 25755
rect 10500 25735 10502 25755
rect 10524 25735 10526 25755
rect 10572 25735 10574 25755
rect 10596 25735 10598 25755
rect 10620 25735 10622 25755
rect 10668 25735 10670 25755
rect 10692 25735 10694 25755
rect 10716 25735 10718 25755
rect 10788 25735 10790 25755
rect 10836 25735 10838 25755
rect 10956 25735 10958 25755
rect 11004 25735 11006 25755
rect 11052 25735 11054 25755
rect 11076 25735 11078 25755
rect 11100 25735 11102 25755
rect 11172 25735 11174 25755
rect 11220 25735 11222 25755
rect 11340 25735 11342 25755
rect 11436 25735 11438 25755
rect 11532 25735 11534 25755
rect 11580 25735 11582 25755
rect 11628 25735 11630 25755
rect 11676 25735 11678 25755
rect 11724 25735 11726 25755
rect 11772 25735 11774 25755
rect 11796 25735 11798 25755
rect 11892 25735 11894 25755
rect 11988 25735 11990 25755
rect 12060 25735 12062 25755
rect 12132 25735 12134 25755
rect 12228 25735 12230 25755
rect 12276 25735 12278 25755
rect 12324 25735 12326 25755
rect 12420 25735 12422 25755
rect 12444 25735 12446 25755
rect 12492 25735 12494 25755
rect 12516 25735 12518 25755
rect 12540 25735 12542 25755
rect 12588 25735 12590 25755
rect 12636 25735 12638 25755
rect 12732 25735 12734 25755
rect 12756 25735 12758 25755
rect 12804 25735 12806 25755
rect 12828 25735 12830 25755
rect 12852 25735 12854 25755
rect 12948 25735 12950 25755
rect 12972 25735 12974 25755
rect 13044 25735 13046 25755
rect 13068 25735 13070 25755
rect 13116 25735 13118 25755
rect 13284 25735 13286 25755
rect 13332 25735 13334 25755
rect 13572 25735 13574 25755
rect 13644 25736 13646 25755
rect 13609 25735 13667 25736
rect 13668 25735 13670 25755
rect 13764 25735 13766 25755
rect 13812 25735 13814 25755
rect 13860 25735 13862 25755
rect 13908 25735 13910 25755
rect 13956 25735 13958 25755
rect 14004 25735 14006 25755
rect 14100 25735 14102 25755
rect 14196 25735 14198 25755
rect 14292 25735 14294 25755
rect 15180 25735 15182 25755
rect 15252 25735 15254 25755
rect 15276 25735 15278 25755
rect 15420 25735 15422 25755
rect 15492 25735 15494 25755
rect 15540 25735 15542 25755
rect 15636 25735 15638 25755
rect 15660 25735 15662 25755
rect 15708 25735 15710 25755
rect 15732 25735 15734 25755
rect 15756 25735 15758 25755
rect 15804 25735 15806 25755
rect 15828 25735 15830 25755
rect 15852 25735 15854 25755
rect 15900 25735 15902 25755
rect 15948 25735 15950 25755
rect 15996 25735 15998 25755
rect 16044 25735 16046 25755
rect 16164 25735 16166 25755
rect 16260 25735 16262 25755
rect 16308 25735 16310 25755
rect 16332 25735 16334 25755
rect 16356 25735 16358 25755
rect 16404 25735 16406 25755
rect 16452 25735 16454 25755
rect 16548 25735 16550 25755
rect 16572 25735 16574 25755
rect 16620 25735 16622 25755
rect 16668 25735 16670 25755
rect 16716 25735 16718 25755
rect 16764 25735 16766 25755
rect 16812 25735 16814 25755
rect 16884 25735 16886 25755
rect 16908 25735 16910 25755
rect 16980 25735 16982 25755
rect 17052 25735 17054 25755
rect 17196 25735 17198 25755
rect 17220 25735 17222 25755
rect 17292 25735 17294 25755
rect 17316 25735 17318 25755
rect 18084 25735 18086 25755
rect 18132 25735 18134 25755
rect 18228 25735 18230 25755
rect 18396 25735 18398 25755
rect 18492 25735 18494 25755
rect 18516 25735 18518 25755
rect 18564 25735 18566 25755
rect 18612 25735 18614 25755
rect 18660 25735 18662 25755
rect 18708 25735 18710 25755
rect 18756 25735 18758 25755
rect 18804 25735 18806 25755
rect 18852 25735 18854 25755
rect 18900 25735 18902 25755
rect 18996 25735 18998 25755
rect 19020 25735 19022 25755
rect 19092 25735 19094 25755
rect 19116 25735 19118 25755
rect 19140 25735 19142 25755
rect 19188 25735 19190 25755
rect 19236 25735 19238 25755
rect 19332 25735 19334 25755
rect 19476 25735 19478 25755
rect 19788 25735 19790 25755
rect 19836 25735 19838 25755
rect 19860 25735 19862 25755
rect 19884 25735 19886 25755
rect 19932 25735 19934 25755
rect 19956 25735 19958 25755
rect 19980 25735 19982 25755
rect 20028 25735 20030 25755
rect 20052 25735 20054 25755
rect 20076 25735 20078 25755
rect 20148 25735 20150 25755
rect 20172 25735 20174 25755
rect 20196 25735 20198 25755
rect 20268 25735 20270 25755
rect 20292 25735 20294 25755
rect 20388 25735 20390 25755
rect 20412 25735 20414 25755
rect 20508 25735 20510 25755
rect 20556 25735 20558 25755
rect 20604 25735 20606 25755
rect 20916 25735 20918 25755
rect 20964 25735 20966 25755
rect 21012 25735 21014 25755
rect 21060 25735 21062 25755
rect 21108 25735 21110 25755
rect 21159 25752 21173 25755
rect 21204 25735 21206 25755
rect 21300 25735 21302 25755
rect 21324 25735 21326 25755
rect 21444 25735 21446 25755
rect 21468 25735 21470 25755
rect 21481 25735 21539 25736
rect 21564 25735 21566 25755
rect 21612 25735 21614 25755
rect 21684 25735 21686 25755
rect 21708 25735 21710 25755
rect 21828 25735 21830 25755
rect 21924 25735 21926 25755
rect 22068 25735 22070 25755
rect 22188 25735 22190 25755
rect 22212 25735 22214 25755
rect 22884 25735 22886 25755
rect 22980 25735 22982 25755
rect 23076 25735 23078 25755
rect 23100 25735 23102 25755
rect 23124 25735 23126 25755
rect 23244 25735 23246 25755
rect 23340 25735 23342 25755
rect 23412 25735 23414 25755
rect 23508 25735 23510 25755
rect 23556 25735 23558 25755
rect 23652 25735 23654 25755
rect 23676 25735 23678 25755
rect 23724 25735 23726 25755
rect 23772 25735 23774 25755
rect 23820 25735 23822 25755
rect 23916 25735 23918 25755
rect 24012 25735 24014 25755
rect 24039 25752 24053 25755
rect 24063 25755 27419 25759
rect 24063 25752 24077 25755
rect 24084 25752 24087 25755
rect 24049 25735 24107 25736
rect 24396 25735 24398 25755
rect 24492 25735 24494 25755
rect 24516 25735 24518 25755
rect 24588 25735 24590 25755
rect 24612 25735 24614 25755
rect 24684 25735 24686 25755
rect 24732 25735 24734 25755
rect 24756 25735 24758 25755
rect 24780 25735 24782 25755
rect 24852 25735 24854 25755
rect 24876 25735 24878 25755
rect 24972 25735 24974 25755
rect 24996 25735 24998 25755
rect 25068 25735 25070 25755
rect 25164 25735 25166 25755
rect 25260 25735 25262 25755
rect 25284 25735 25286 25755
rect 25356 25735 25358 25755
rect 25380 25735 25382 25755
rect 25404 25735 25406 25755
rect 25500 25735 25502 25755
rect 25596 25735 25598 25755
rect 27036 25735 27038 25755
rect 27108 25735 27110 25755
rect 27324 25736 27326 25755
rect 27385 25750 27388 25755
rect 27396 25750 27398 25755
rect 27395 25736 27398 25750
rect 27313 25735 27347 25736
rect -16449 25731 3869 25735
rect -16449 25728 -16435 25731
rect -16404 25728 -16402 25731
rect -16404 25711 -16401 25728
rect -16356 25711 -16354 25731
rect -16308 25711 -16306 25731
rect -16284 25711 -16282 25731
rect -16260 25711 -16258 25731
rect -15324 25711 -15322 25731
rect -15108 25711 -15106 25731
rect -14772 25711 -14770 25731
rect -14436 25711 -14434 25731
rect -14433 25728 -14419 25731
rect -14340 25711 -14338 25731
rect -13991 25726 -13988 25731
rect -13980 25726 -13978 25731
rect -13981 25712 -13978 25726
rect -13932 25711 -13930 25731
rect -13884 25728 -13882 25731
rect -13884 25711 -13881 25728
rect -13788 25711 -13786 25731
rect -13572 25711 -13570 25731
rect -13356 25711 -13354 25731
rect -13199 25711 -13141 25712
rect -13068 25711 -13066 25731
rect -12780 25711 -12778 25731
rect -12756 25711 -12754 25731
rect -12660 25711 -12658 25731
rect -12564 25711 -12562 25731
rect -12492 25711 -12490 25731
rect -12396 25711 -12394 25731
rect -12348 25711 -12346 25731
rect -12252 25711 -12250 25731
rect -12156 25711 -12154 25731
rect -12060 25711 -12058 25731
rect -11844 25711 -11842 25731
rect -11676 25711 -11674 25731
rect -11556 25711 -11554 25731
rect -11508 25711 -11506 25731
rect -11436 25711 -11434 25731
rect -11412 25711 -11410 25731
rect -11340 25711 -11338 25731
rect -11196 25711 -11194 25731
rect -11124 25711 -11122 25731
rect -11100 25711 -11098 25731
rect -11028 25711 -11026 25731
rect -10740 25711 -10738 25731
rect -10668 25711 -10666 25731
rect -10644 25711 -10642 25731
rect -9996 25711 -9994 25731
rect -9828 25711 -9826 25731
rect -9732 25711 -9730 25731
rect -9516 25711 -9514 25731
rect -9468 25711 -9466 25731
rect -9420 25712 -9418 25731
rect -9263 25726 -9260 25731
rect -9252 25726 -9250 25731
rect -9253 25712 -9250 25726
rect -9455 25711 -9397 25712
rect -9180 25711 -9177 25728
rect -8604 25711 -8602 25731
rect -8484 25711 -8482 25731
rect -8436 25711 -8434 25731
rect -8388 25711 -8386 25731
rect -8364 25711 -8362 25731
rect -8340 25711 -8338 25731
rect -8268 25711 -8266 25731
rect -8100 25711 -8098 25731
rect -8052 25711 -8050 25731
rect -7932 25711 -7930 25731
rect -7692 25711 -7690 25731
rect -7620 25711 -7618 25731
rect -7524 25711 -7522 25731
rect -7356 25711 -7354 25731
rect -7308 25711 -7306 25731
rect -7212 25711 -7210 25731
rect -7116 25711 -7114 25731
rect -7068 25711 -7066 25731
rect -6972 25711 -6970 25731
rect -6948 25711 -6946 25731
rect -6876 25711 -6874 25731
rect -6852 25711 -6850 25731
rect -6780 25711 -6778 25731
rect -6756 25711 -6754 25731
rect -6660 25711 -6658 25731
rect -6612 25711 -6610 25731
rect -6516 25711 -6514 25731
rect -6431 25726 -6428 25731
rect -6420 25726 -6418 25731
rect -6421 25712 -6418 25726
rect -6372 25711 -6370 25731
rect -6324 25728 -6322 25731
rect -6324 25711 -6321 25728
rect -6156 25711 -6154 25731
rect -6060 25711 -6058 25731
rect -6036 25711 -6034 25731
rect -5892 25711 -5890 25731
rect -5652 25711 -5650 25731
rect -5268 25711 -5266 25731
rect -5196 25711 -5194 25731
rect -5172 25711 -5170 25731
rect -5100 25711 -5098 25731
rect -5076 25711 -5074 25731
rect -4980 25711 -4978 25731
rect -4956 25711 -4954 25731
rect -4860 25711 -4858 25731
rect -4644 25711 -4642 25731
rect -4548 25711 -4546 25731
rect -4500 25711 -4498 25731
rect -4404 25711 -4402 25731
rect -4308 25711 -4306 25731
rect -4260 25711 -4258 25731
rect -4164 25711 -4162 25731
rect -4020 25711 -4018 25731
rect -3876 25711 -3874 25731
rect -3732 25711 -3730 25731
rect -3588 25711 -3586 25731
rect -3564 25711 -3562 25731
rect -3516 25711 -3514 25731
rect -3492 25711 -3490 25731
rect -3468 25711 -3466 25731
rect -3420 25711 -3418 25731
rect -3324 25711 -3322 25731
rect -3228 25711 -3226 25731
rect -3132 25711 -3130 25731
rect -3081 25728 -3067 25731
rect -3060 25728 -3057 25731
rect -3012 25711 -3010 25731
rect -2964 25711 -2962 25731
rect -2916 25711 -2914 25731
rect -2892 25711 -2890 25731
rect -2868 25711 -2866 25731
rect -2820 25711 -2818 25731
rect -2796 25711 -2794 25731
rect -2772 25711 -2770 25731
rect -2676 25711 -2674 25731
rect -2580 25711 -2578 25731
rect -2364 25711 -2362 25731
rect -2327 25726 -2324 25731
rect -2317 25712 -2314 25726
rect -2316 25711 -2314 25712
rect -2268 25711 -2266 25731
rect -2244 25711 -2242 25731
rect -2172 25711 -2170 25731
rect -2148 25711 -2146 25731
rect -2076 25711 -2074 25731
rect -2052 25711 -2050 25731
rect -1980 25711 -1978 25731
rect -1884 25711 -1882 25731
rect -1761 25728 -1747 25731
rect -1572 25711 -1570 25731
rect -1476 25711 -1474 25731
rect -1380 25711 -1378 25731
rect -1356 25711 -1354 25731
rect -1308 25711 -1306 25731
rect -1260 25711 -1258 25731
rect -1140 25711 -1138 25731
rect -852 25712 -850 25731
rect -887 25711 -829 25712
rect -756 25711 -754 25731
rect -708 25711 -706 25731
rect -612 25711 -610 25731
rect -588 25711 -586 25731
rect -540 25711 -538 25731
rect -492 25711 -490 25731
rect -444 25711 -442 25731
rect -396 25711 -394 25731
rect -300 25711 -298 25731
rect -276 25711 -274 25731
rect -228 25711 -226 25731
rect -12 25711 -10 25731
rect 156 25711 158 25731
rect 204 25711 206 25731
rect 252 25711 254 25731
rect 348 25711 350 25731
rect 468 25711 470 25731
rect 492 25711 494 25731
rect 564 25711 566 25731
rect 588 25711 590 25731
rect 636 25711 638 25731
rect 660 25711 662 25731
rect 732 25711 734 25731
rect 1009 25726 1012 25731
rect 1020 25726 1022 25731
rect 1019 25712 1022 25726
rect 1092 25711 1094 25731
rect 1105 25726 1108 25731
rect 1116 25728 1118 25731
rect 1212 25728 1214 25731
rect 1116 25726 1119 25728
rect 1115 25712 1119 25726
rect 1212 25711 1215 25728
rect 1308 25711 1310 25731
rect 1332 25711 1334 25731
rect 1380 25711 1382 25731
rect 1428 25711 1430 25731
rect 1476 25711 1478 25731
rect 1548 25728 1550 25731
rect 1548 25711 1551 25728
rect 1644 25711 1646 25731
rect 1692 25711 1694 25731
rect 1740 25711 1742 25731
rect 1788 25711 1790 25731
rect 2028 25711 2030 25731
rect 2076 25711 2078 25731
rect 2100 25711 2102 25731
rect 2124 25711 2126 25731
rect 2172 25711 2174 25731
rect 2220 25711 2222 25731
rect 2268 25712 2270 25731
rect 2233 25711 2291 25712
rect 2316 25711 2318 25731
rect 2364 25711 2366 25731
rect 2412 25711 2414 25731
rect 2460 25711 2462 25731
rect 2508 25711 2510 25731
rect 2580 25711 2582 25731
rect 2604 25711 2606 25731
rect 2676 25711 2678 25731
rect 2700 25711 2702 25731
rect 2748 25711 2750 25731
rect 2772 25711 2774 25731
rect 2796 25711 2798 25731
rect 2844 25711 2846 25731
rect 2868 25711 2870 25731
rect 2892 25711 2894 25731
rect 2940 25711 2942 25731
rect 3012 25711 3014 25731
rect 3049 25711 3083 25712
rect 3108 25711 3110 25731
rect 3156 25711 3158 25731
rect 3252 25711 3254 25731
rect 3348 25711 3350 25731
rect 3396 25711 3398 25731
rect 3564 25711 3566 25731
rect 3636 25711 3638 25731
rect 3660 25711 3662 25731
rect 3732 25711 3734 25731
rect 3828 25711 3830 25731
rect 3855 25728 3869 25731
rect 3879 25731 27347 25735
rect 3879 25728 3893 25731
rect 3924 25711 3926 25731
rect 4020 25711 4022 25731
rect 4044 25711 4046 25731
rect 4092 25711 4094 25731
rect 4116 25711 4118 25731
rect 4140 25711 4142 25731
rect 4188 25711 4190 25731
rect 4212 25711 4214 25731
rect 4236 25711 4238 25731
rect 4308 25711 4310 25731
rect 4332 25711 4334 25731
rect 4404 25711 4406 25731
rect 4500 25711 4502 25731
rect 4596 25711 4598 25731
rect 4692 25711 4694 25731
rect 4860 25711 4862 25731
rect 4956 25711 4958 25731
rect 4980 25711 4982 25731
rect 5004 25711 5006 25731
rect 5041 25726 5044 25731
rect 5065 25726 5068 25731
rect 5076 25726 5078 25731
rect 5051 25712 5054 25726
rect 5075 25712 5078 25726
rect 5052 25711 5054 25712
rect 5100 25711 5102 25731
rect 5124 25711 5126 25731
rect 5172 25728 5174 25731
rect 5172 25711 5175 25728
rect 5220 25711 5222 25731
rect 5268 25711 5270 25731
rect 5388 25711 5390 25731
rect 5484 25711 5486 25731
rect 5508 25711 5510 25731
rect 5532 25711 5534 25731
rect 5628 25711 5630 25731
rect 5652 25711 5654 25731
rect 5748 25711 5750 25731
rect 5796 25711 5798 25731
rect 5844 25711 5846 25731
rect 5892 25711 5894 25731
rect 6132 25711 6134 25731
rect 6180 25711 6182 25731
rect 6228 25711 6230 25731
rect 6252 25711 6254 25731
rect 6276 25711 6278 25731
rect 6324 25711 6326 25731
rect 6372 25711 6374 25731
rect 6492 25711 6494 25731
rect 6588 25711 6590 25731
rect 6612 25711 6614 25731
rect 6660 25711 6662 25731
rect 6684 25711 6686 25731
rect 6708 25711 6710 25731
rect 6780 25711 6782 25731
rect 6804 25711 6806 25731
rect 6900 25711 6902 25731
rect 6924 25711 6926 25731
rect 7020 25711 7022 25731
rect 7033 25711 7115 25712
rect 7140 25711 7142 25731
rect 7236 25711 7238 25731
rect 7332 25711 7334 25731
rect 7380 25711 7382 25731
rect 7428 25711 7430 25731
rect 7452 25711 7454 25731
rect 7476 25711 7478 25731
rect 7524 25711 7526 25731
rect 7548 25711 7550 25731
rect 7572 25711 7574 25731
rect 7620 25711 7622 25731
rect 7644 25711 7646 25731
rect 7668 25711 7670 25731
rect 7788 25711 7790 25731
rect 7884 25711 7886 25731
rect 7956 25711 7958 25731
rect 7980 25711 7982 25731
rect 8028 25711 8030 25731
rect 8196 25711 8198 25731
rect 8244 25711 8246 25731
rect 8268 25711 8270 25731
rect 8292 25711 8294 25731
rect 8340 25711 8342 25731
rect 8364 25711 8366 25731
rect 8388 25711 8390 25731
rect 8436 25711 8438 25731
rect 8604 25711 8606 25731
rect 8652 25711 8654 25731
rect 8700 25711 8702 25731
rect 8724 25711 8726 25731
rect 8748 25711 8750 25731
rect 8820 25711 8822 25731
rect 8844 25711 8846 25731
rect 8868 25711 8870 25731
rect 9516 25711 9518 25731
rect 9612 25711 9614 25731
rect 9660 25711 9662 25731
rect 9684 25711 9686 25731
rect 9708 25711 9710 25731
rect 9756 25711 9758 25731
rect 9780 25711 9782 25731
rect 9804 25711 9806 25731
rect 9852 25711 9854 25731
rect 9900 25711 9902 25731
rect 9948 25711 9950 25731
rect 9996 25711 9998 25731
rect 10068 25711 10070 25731
rect 10092 25711 10094 25731
rect 10116 25711 10118 25731
rect 10164 25711 10166 25731
rect 10188 25711 10190 25731
rect 10212 25711 10214 25731
rect 10284 25711 10286 25731
rect 10308 25711 10310 25731
rect 10332 25711 10334 25731
rect 10380 25711 10382 25731
rect 10404 25711 10406 25731
rect 10428 25711 10430 25731
rect 10476 25711 10478 25731
rect 10500 25711 10502 25731
rect 10524 25711 10526 25731
rect 10572 25711 10574 25731
rect 10596 25711 10598 25731
rect 10620 25711 10622 25731
rect 10668 25711 10670 25731
rect 10692 25711 10694 25731
rect 10716 25711 10718 25731
rect 10788 25711 10790 25731
rect 10836 25711 10838 25731
rect 10956 25711 10958 25731
rect 11004 25711 11006 25731
rect 11052 25711 11054 25731
rect 11076 25711 11078 25731
rect 11100 25711 11102 25731
rect 11172 25711 11174 25731
rect 11220 25711 11222 25731
rect 11340 25711 11342 25731
rect 11436 25711 11438 25731
rect 11532 25711 11534 25731
rect 11580 25711 11582 25731
rect 11628 25711 11630 25731
rect 11676 25711 11678 25731
rect 11724 25711 11726 25731
rect 11772 25711 11774 25731
rect 11796 25711 11798 25731
rect 11892 25711 11894 25731
rect 11988 25711 11990 25731
rect 12060 25711 12062 25731
rect 12132 25711 12134 25731
rect 12228 25711 12230 25731
rect 12276 25711 12278 25731
rect 12324 25711 12326 25731
rect 12420 25711 12422 25731
rect 12444 25711 12446 25731
rect 12492 25711 12494 25731
rect 12516 25711 12518 25731
rect 12540 25711 12542 25731
rect 12588 25711 12590 25731
rect 12636 25711 12638 25731
rect 12732 25711 12734 25731
rect 12756 25711 12758 25731
rect 12804 25711 12806 25731
rect 12828 25711 12830 25731
rect 12852 25711 12854 25731
rect 12948 25711 12950 25731
rect 12972 25711 12974 25731
rect 13044 25711 13046 25731
rect 13068 25711 13070 25731
rect 13116 25711 13118 25731
rect 13284 25711 13286 25731
rect 13332 25711 13334 25731
rect 13572 25711 13574 25731
rect 13609 25726 13612 25731
rect 13633 25726 13636 25731
rect 13644 25726 13646 25731
rect 13619 25712 13622 25726
rect 13643 25712 13646 25726
rect 13620 25711 13622 25712
rect 13668 25711 13670 25731
rect 13716 25711 13719 25728
rect 13764 25711 13766 25731
rect 13812 25712 13814 25731
rect 13801 25711 13835 25712
rect 13860 25711 13862 25731
rect 13908 25711 13910 25731
rect 13956 25711 13958 25731
rect 14004 25711 14006 25731
rect 14100 25711 14102 25731
rect 14196 25711 14198 25731
rect 14292 25711 14294 25731
rect 15180 25711 15182 25731
rect 15252 25712 15254 25731
rect 15241 25711 15275 25712
rect 15276 25711 15278 25731
rect 15420 25711 15422 25731
rect 15492 25711 15494 25731
rect 15540 25711 15542 25731
rect 15636 25711 15638 25731
rect 15660 25711 15662 25731
rect 15708 25711 15710 25731
rect 15732 25711 15734 25731
rect 15756 25711 15758 25731
rect 15804 25711 15806 25731
rect 15828 25711 15830 25731
rect 15852 25711 15854 25731
rect 15900 25711 15902 25731
rect 15948 25711 15950 25731
rect 15996 25712 15998 25731
rect 15961 25711 16019 25712
rect 16044 25711 16046 25731
rect 16164 25711 16166 25731
rect 16260 25711 16262 25731
rect 16308 25711 16310 25731
rect 16332 25711 16334 25731
rect 16356 25711 16358 25731
rect 16404 25711 16406 25731
rect 16452 25711 16454 25731
rect 16548 25711 16550 25731
rect 16572 25711 16574 25731
rect 16620 25711 16622 25731
rect 16668 25711 16670 25731
rect 16716 25711 16718 25731
rect 16764 25711 16766 25731
rect 16812 25711 16814 25731
rect 16884 25711 16886 25731
rect 16908 25711 16910 25731
rect 16980 25711 16982 25731
rect 17052 25711 17054 25731
rect 17196 25711 17198 25731
rect 17220 25711 17222 25731
rect 17292 25711 17294 25731
rect 17316 25711 17318 25731
rect 18084 25711 18086 25731
rect 18132 25711 18134 25731
rect 18228 25711 18230 25731
rect 18396 25711 18398 25731
rect 18492 25711 18494 25731
rect 18516 25711 18518 25731
rect 18564 25711 18566 25731
rect 18612 25711 18614 25731
rect 18660 25711 18662 25731
rect 18708 25711 18710 25731
rect 18756 25711 18758 25731
rect 18804 25711 18806 25731
rect 18852 25711 18854 25731
rect 18900 25711 18902 25731
rect 18996 25711 18998 25731
rect 19020 25711 19022 25731
rect 19092 25711 19094 25731
rect 19116 25711 19118 25731
rect 19140 25711 19142 25731
rect 19188 25711 19190 25731
rect 19236 25711 19238 25731
rect 19332 25711 19334 25731
rect 19476 25711 19478 25731
rect 19788 25711 19790 25731
rect 19836 25711 19838 25731
rect 19860 25711 19862 25731
rect 19884 25711 19886 25731
rect 19932 25711 19934 25731
rect 19956 25711 19958 25731
rect 19980 25711 19982 25731
rect 20028 25711 20030 25731
rect 20052 25711 20054 25731
rect 20076 25711 20078 25731
rect 20148 25711 20150 25731
rect 20172 25711 20174 25731
rect 20196 25711 20198 25731
rect 20268 25711 20270 25731
rect 20292 25711 20294 25731
rect 20388 25711 20390 25731
rect 20412 25711 20414 25731
rect 20508 25711 20510 25731
rect 20556 25711 20558 25731
rect 20604 25711 20606 25731
rect 20916 25711 20918 25731
rect 20964 25711 20966 25731
rect 21012 25711 21014 25731
rect 21060 25711 21062 25731
rect 21108 25711 21110 25731
rect 21204 25711 21206 25731
rect 21300 25711 21302 25731
rect 21324 25711 21326 25731
rect 21444 25711 21446 25731
rect 21468 25711 21470 25731
rect 21564 25711 21566 25731
rect 21612 25728 21614 25731
rect 21588 25711 21591 25728
rect 21612 25711 21615 25728
rect 21684 25711 21686 25731
rect 21708 25711 21710 25731
rect 21828 25711 21830 25731
rect 21924 25711 21926 25731
rect 22068 25711 22070 25731
rect 22188 25711 22190 25731
rect 22212 25711 22214 25731
rect 22884 25711 22886 25731
rect 22980 25711 22982 25731
rect 23076 25711 23078 25731
rect 23100 25711 23102 25731
rect 23124 25711 23126 25731
rect 23244 25711 23246 25731
rect 23340 25711 23342 25731
rect 23412 25711 23414 25731
rect 23508 25711 23510 25731
rect 23556 25711 23558 25731
rect 23652 25711 23654 25731
rect 23676 25711 23678 25731
rect 23724 25711 23726 25731
rect 23772 25711 23774 25731
rect 23820 25711 23822 25731
rect 23916 25711 23918 25731
rect 24012 25711 24014 25731
rect 24049 25726 24052 25731
rect 24059 25712 24062 25726
rect 24060 25711 24062 25712
rect 24156 25711 24159 25728
rect 24289 25711 24323 25712
rect 24396 25711 24398 25731
rect 24492 25711 24494 25731
rect 24516 25711 24518 25731
rect 24588 25711 24590 25731
rect 24612 25711 24614 25731
rect 24684 25711 24686 25731
rect 24732 25711 24734 25731
rect 24756 25711 24758 25731
rect 24780 25711 24782 25731
rect 24852 25711 24854 25731
rect 24876 25711 24878 25731
rect 24972 25711 24974 25731
rect 24996 25712 24998 25731
rect 24985 25711 25019 25712
rect 25068 25711 25070 25731
rect 25164 25711 25166 25731
rect 25260 25711 25262 25731
rect 25284 25711 25286 25731
rect 25356 25711 25358 25731
rect 25380 25711 25382 25731
rect 25404 25711 25406 25731
rect 25500 25711 25502 25731
rect 25596 25711 25598 25731
rect 27036 25711 27038 25731
rect 27108 25711 27110 25731
rect 27313 25726 27316 25731
rect 27324 25726 27326 25731
rect 27323 25712 27326 25726
rect 27289 25711 27323 25712
rect -16425 25707 -15979 25711
rect -16425 25704 -16411 25707
rect -16404 25704 -16401 25707
rect -16356 25704 -16354 25707
rect -16377 25687 -16357 25688
rect -16356 25687 -16353 25704
rect -16308 25687 -16306 25707
rect -16284 25687 -16282 25707
rect -16260 25687 -16258 25707
rect -15993 25704 -15979 25707
rect -15969 25707 -13915 25711
rect -15969 25704 -15955 25707
rect -15324 25687 -15322 25707
rect -15108 25687 -15106 25707
rect -14807 25687 -14773 25688
rect -14772 25687 -14770 25707
rect -14687 25687 -14629 25688
rect -14436 25687 -14434 25707
rect -14340 25687 -14338 25707
rect -13932 25687 -13930 25707
rect -13929 25704 -13915 25707
rect -13905 25707 -9187 25711
rect -13905 25704 -13891 25707
rect -13884 25704 -13881 25707
rect -13788 25687 -13786 25707
rect -13572 25687 -13570 25707
rect -13356 25687 -13354 25707
rect -13068 25704 -13066 25707
rect -13068 25687 -13065 25704
rect -12780 25687 -12778 25707
rect -12756 25687 -12754 25707
rect -12660 25687 -12658 25707
rect -12564 25687 -12562 25707
rect -12492 25687 -12490 25707
rect -12396 25687 -12394 25707
rect -12348 25687 -12346 25707
rect -12252 25687 -12250 25707
rect -12156 25687 -12154 25707
rect -12060 25687 -12058 25707
rect -12033 25704 -12019 25707
rect -11844 25687 -11842 25707
rect -11676 25687 -11674 25707
rect -11556 25687 -11554 25707
rect -11508 25687 -11506 25707
rect -11436 25687 -11434 25707
rect -11412 25687 -11410 25707
rect -11340 25687 -11338 25707
rect -11196 25687 -11194 25707
rect -11124 25687 -11122 25707
rect -11100 25687 -11098 25707
rect -11028 25687 -11026 25707
rect -10740 25687 -10738 25707
rect -10668 25687 -10666 25707
rect -10644 25687 -10642 25707
rect -9996 25687 -9994 25707
rect -9911 25687 -9853 25688
rect -9828 25687 -9826 25707
rect -9732 25687 -9730 25707
rect -9516 25687 -9514 25707
rect -9468 25687 -9466 25707
rect -9431 25702 -9428 25707
rect -9420 25702 -9418 25707
rect -9201 25704 -9187 25707
rect -9180 25707 -6355 25711
rect -9180 25704 -9163 25707
rect -9421 25688 -9418 25702
rect -9348 25687 -9345 25704
rect -9180 25687 -9178 25704
rect -8604 25687 -8602 25707
rect -8484 25687 -8482 25707
rect -8436 25687 -8434 25707
rect -8388 25687 -8386 25707
rect -8364 25687 -8362 25707
rect -8340 25687 -8338 25707
rect -8268 25687 -8266 25707
rect -8100 25687 -8098 25707
rect -8052 25687 -8050 25707
rect -8015 25687 -7957 25688
rect -7932 25687 -7930 25707
rect -7692 25687 -7690 25707
rect -7620 25687 -7618 25707
rect -7524 25687 -7522 25707
rect -7356 25687 -7354 25707
rect -7308 25687 -7306 25707
rect -7212 25687 -7210 25707
rect -7116 25687 -7114 25707
rect -7068 25687 -7066 25707
rect -6972 25687 -6970 25707
rect -6948 25687 -6946 25707
rect -6876 25687 -6874 25707
rect -6852 25687 -6850 25707
rect -6780 25687 -6778 25707
rect -6756 25687 -6754 25707
rect -6660 25687 -6658 25707
rect -6612 25687 -6610 25707
rect -6516 25687 -6514 25707
rect -6372 25687 -6370 25707
rect -6369 25704 -6355 25707
rect -6345 25707 -2227 25711
rect -6345 25704 -6331 25707
rect -6324 25704 -6321 25707
rect -6156 25687 -6154 25707
rect -6060 25687 -6058 25707
rect -6036 25687 -6034 25707
rect -5892 25687 -5890 25707
rect -5652 25687 -5650 25707
rect -5268 25687 -5266 25707
rect -5196 25687 -5194 25707
rect -5172 25687 -5170 25707
rect -5100 25687 -5098 25707
rect -5076 25687 -5074 25707
rect -4980 25687 -4978 25707
rect -4956 25687 -4954 25707
rect -4860 25687 -4858 25707
rect -4644 25687 -4642 25707
rect -4548 25687 -4546 25707
rect -4500 25687 -4498 25707
rect -4404 25687 -4402 25707
rect -4308 25687 -4306 25707
rect -4260 25687 -4258 25707
rect -4164 25687 -4162 25707
rect -4020 25687 -4018 25707
rect -3876 25687 -3874 25707
rect -3732 25687 -3730 25707
rect -3588 25687 -3586 25707
rect -3564 25687 -3562 25707
rect -3516 25687 -3514 25707
rect -3492 25687 -3490 25707
rect -3468 25687 -3466 25707
rect -3420 25687 -3418 25707
rect -3324 25687 -3322 25707
rect -3228 25687 -3226 25707
rect -3132 25687 -3130 25707
rect -3012 25687 -3010 25707
rect -2964 25687 -2962 25707
rect -2916 25687 -2914 25707
rect -2892 25687 -2890 25707
rect -2868 25687 -2866 25707
rect -2820 25687 -2818 25707
rect -2796 25687 -2794 25707
rect -2772 25687 -2770 25707
rect -2676 25687 -2674 25707
rect -2580 25687 -2578 25707
rect -2364 25687 -2362 25707
rect -2316 25687 -2314 25707
rect -2268 25687 -2266 25707
rect -2244 25687 -2242 25707
rect -2241 25704 -2227 25707
rect -2217 25707 5141 25711
rect -2217 25704 -2203 25707
rect -2172 25687 -2170 25707
rect -2148 25687 -2146 25707
rect -2076 25687 -2074 25707
rect -2052 25687 -2050 25707
rect -1980 25687 -1978 25707
rect -1884 25687 -1882 25707
rect -1572 25687 -1570 25707
rect -1476 25687 -1474 25707
rect -1380 25687 -1378 25707
rect -1356 25687 -1354 25707
rect -1308 25687 -1306 25707
rect -1260 25687 -1258 25707
rect -1140 25687 -1138 25707
rect -945 25704 -931 25707
rect -863 25702 -860 25707
rect -852 25702 -850 25707
rect -853 25688 -850 25702
rect -756 25704 -754 25707
rect -756 25687 -753 25704
rect -708 25687 -706 25707
rect -612 25687 -610 25707
rect -588 25687 -586 25707
rect -540 25687 -538 25707
rect -492 25687 -490 25707
rect -444 25687 -442 25707
rect -396 25687 -394 25707
rect -300 25687 -298 25707
rect -276 25687 -274 25707
rect -228 25687 -226 25707
rect -12 25687 -10 25707
rect 156 25687 158 25707
rect 204 25687 206 25707
rect 252 25687 254 25707
rect 348 25687 350 25707
rect 468 25687 470 25707
rect 492 25687 494 25707
rect 564 25687 566 25707
rect 588 25687 590 25707
rect 636 25687 638 25707
rect 660 25687 662 25707
rect 732 25687 734 25707
rect 1092 25687 1094 25707
rect 1095 25704 1109 25707
rect 1191 25704 1205 25707
rect 1212 25704 1215 25707
rect 1308 25687 1310 25707
rect 1332 25687 1334 25707
rect 1380 25687 1382 25707
rect 1428 25687 1430 25707
rect 1476 25687 1478 25707
rect 1527 25704 1541 25707
rect 1548 25704 1551 25707
rect 1644 25687 1646 25707
rect 1692 25687 1694 25707
rect 1740 25687 1742 25707
rect 1788 25687 1790 25707
rect 2028 25687 2030 25707
rect 2076 25687 2078 25707
rect 2100 25687 2102 25707
rect 2124 25687 2126 25707
rect 2172 25687 2174 25707
rect 2220 25687 2222 25707
rect 2257 25702 2260 25707
rect 2268 25702 2270 25707
rect 2267 25688 2270 25702
rect 2316 25687 2318 25707
rect 2364 25704 2366 25707
rect 2364 25687 2367 25704
rect 2412 25687 2414 25707
rect 2460 25687 2462 25707
rect 2508 25687 2510 25707
rect 2580 25687 2582 25707
rect 2604 25687 2606 25707
rect 2676 25687 2678 25707
rect 2700 25687 2702 25707
rect 2748 25687 2750 25707
rect 2772 25687 2774 25707
rect 2796 25687 2798 25707
rect 2844 25687 2846 25707
rect 2868 25687 2870 25707
rect 2892 25687 2894 25707
rect 2940 25687 2942 25707
rect 3012 25687 3014 25707
rect 3108 25687 3110 25707
rect 3156 25704 3158 25707
rect 3156 25687 3159 25704
rect 3252 25687 3254 25707
rect 3348 25687 3350 25707
rect 3396 25687 3398 25707
rect 3564 25687 3566 25707
rect 3636 25687 3638 25707
rect 3660 25687 3662 25707
rect 3732 25687 3734 25707
rect 3828 25687 3830 25707
rect 3924 25687 3926 25707
rect 4020 25687 4022 25707
rect 4044 25687 4046 25707
rect 4092 25687 4094 25707
rect 4116 25687 4118 25707
rect 4140 25687 4142 25707
rect 4188 25687 4190 25707
rect 4212 25687 4214 25707
rect 4236 25687 4238 25707
rect 4308 25687 4310 25707
rect 4332 25687 4334 25707
rect 4404 25687 4406 25707
rect 4500 25687 4502 25707
rect 4596 25687 4598 25707
rect 4692 25687 4694 25707
rect 4860 25687 4862 25707
rect 4956 25687 4958 25707
rect 4980 25687 4982 25707
rect 5004 25687 5006 25707
rect 5052 25687 5054 25707
rect 5100 25687 5102 25707
rect 5124 25687 5126 25707
rect 5127 25704 5141 25707
rect 5151 25707 13709 25711
rect 5151 25704 5165 25707
rect 5172 25704 5175 25707
rect 5220 25687 5222 25707
rect 5268 25687 5270 25707
rect 5388 25687 5390 25707
rect 5484 25687 5486 25707
rect 5508 25687 5510 25707
rect 5532 25687 5534 25707
rect 5628 25687 5630 25707
rect 5652 25687 5654 25707
rect 5748 25687 5750 25707
rect 5796 25687 5798 25707
rect 5844 25687 5846 25707
rect 5892 25687 5894 25707
rect 6132 25687 6134 25707
rect 6180 25687 6182 25707
rect 6228 25687 6230 25707
rect 6252 25687 6254 25707
rect 6276 25687 6278 25707
rect 6324 25687 6326 25707
rect 6372 25687 6374 25707
rect 6492 25687 6494 25707
rect 6588 25687 6590 25707
rect 6612 25687 6614 25707
rect 6660 25687 6662 25707
rect 6684 25687 6686 25707
rect 6708 25687 6710 25707
rect 6780 25687 6782 25707
rect 6804 25687 6806 25707
rect 6900 25687 6902 25707
rect 6924 25687 6926 25707
rect 7020 25687 7022 25707
rect 7057 25702 7060 25707
rect 7140 25704 7142 25707
rect 7067 25688 7070 25702
rect 7068 25687 7070 25688
rect 7140 25687 7143 25704
rect 7164 25687 7167 25704
rect 7236 25687 7238 25707
rect 7332 25687 7334 25707
rect 7380 25687 7382 25707
rect 7428 25687 7430 25707
rect 7452 25687 7454 25707
rect 7476 25687 7478 25707
rect 7524 25687 7526 25707
rect 7548 25687 7550 25707
rect 7572 25687 7574 25707
rect 7620 25687 7622 25707
rect 7644 25687 7646 25707
rect 7668 25687 7670 25707
rect 7788 25687 7790 25707
rect 7884 25687 7886 25707
rect 7956 25687 7958 25707
rect 7980 25687 7982 25707
rect 8028 25687 8030 25707
rect 8196 25687 8198 25707
rect 8244 25687 8246 25707
rect 8268 25687 8270 25707
rect 8292 25687 8294 25707
rect 8340 25687 8342 25707
rect 8364 25687 8366 25707
rect 8388 25687 8390 25707
rect 8436 25687 8438 25707
rect 8604 25687 8606 25707
rect 8652 25687 8654 25707
rect 8700 25687 8702 25707
rect 8724 25687 8726 25707
rect 8748 25687 8750 25707
rect 8820 25687 8822 25707
rect 8844 25687 8846 25707
rect 8868 25687 8870 25707
rect 9516 25687 9518 25707
rect 9612 25687 9614 25707
rect 9660 25687 9662 25707
rect 9684 25687 9686 25707
rect 9708 25687 9710 25707
rect 9756 25687 9758 25707
rect 9780 25687 9782 25707
rect 9804 25687 9806 25707
rect 9852 25687 9854 25707
rect 9900 25687 9902 25707
rect 9948 25687 9950 25707
rect 9996 25687 9998 25707
rect 10068 25687 10070 25707
rect 10092 25687 10094 25707
rect 10116 25687 10118 25707
rect 10164 25687 10166 25707
rect 10188 25687 10190 25707
rect 10212 25687 10214 25707
rect 10284 25687 10286 25707
rect 10308 25687 10310 25707
rect 10332 25687 10334 25707
rect 10380 25687 10382 25707
rect 10404 25687 10406 25707
rect 10428 25687 10430 25707
rect 10476 25687 10478 25707
rect 10500 25687 10502 25707
rect 10524 25687 10526 25707
rect 10572 25687 10574 25707
rect 10596 25687 10598 25707
rect 10620 25687 10622 25707
rect 10668 25687 10670 25707
rect 10692 25687 10694 25707
rect 10716 25687 10718 25707
rect 10788 25687 10790 25707
rect 10836 25687 10838 25707
rect 10956 25687 10958 25707
rect 10969 25687 11003 25688
rect 11004 25687 11006 25707
rect 11052 25687 11054 25707
rect 11076 25687 11078 25707
rect 11100 25687 11102 25707
rect 11172 25687 11174 25707
rect 11220 25687 11222 25707
rect 11340 25687 11342 25707
rect 11436 25687 11438 25707
rect 11532 25687 11534 25707
rect 11580 25687 11582 25707
rect 11628 25687 11630 25707
rect 11676 25687 11678 25707
rect 11724 25687 11726 25707
rect 11772 25687 11774 25707
rect 11796 25687 11798 25707
rect 11892 25687 11894 25707
rect 11988 25687 11990 25707
rect 12060 25687 12062 25707
rect 12132 25687 12134 25707
rect 12228 25687 12230 25707
rect 12276 25687 12278 25707
rect 12324 25687 12326 25707
rect 12420 25687 12422 25707
rect 12444 25687 12446 25707
rect 12492 25687 12494 25707
rect 12516 25687 12518 25707
rect 12540 25687 12542 25707
rect 12588 25687 12590 25707
rect 12636 25687 12638 25707
rect 12732 25687 12734 25707
rect 12756 25687 12758 25707
rect 12804 25687 12806 25707
rect 12828 25687 12830 25707
rect 12852 25687 12854 25707
rect 12948 25687 12950 25707
rect 12972 25687 12974 25707
rect 13044 25687 13046 25707
rect 13068 25687 13070 25707
rect 13116 25687 13118 25707
rect 13284 25687 13286 25707
rect 13332 25687 13334 25707
rect 13572 25687 13574 25707
rect 13620 25687 13622 25707
rect 13668 25687 13670 25707
rect 13695 25704 13709 25707
rect 13716 25707 21581 25711
rect 13716 25704 13733 25707
rect 13716 25687 13718 25704
rect 13764 25687 13766 25707
rect 13801 25702 13804 25707
rect 13812 25702 13814 25707
rect 13811 25688 13814 25702
rect 13860 25687 13862 25707
rect 13908 25704 13910 25707
rect 13908 25687 13911 25704
rect 13956 25687 13958 25707
rect 14004 25687 14006 25707
rect 14100 25687 14102 25707
rect 14196 25687 14198 25707
rect 14292 25687 14294 25707
rect 15180 25687 15182 25707
rect 15241 25702 15244 25707
rect 15252 25702 15254 25707
rect 15251 25688 15254 25702
rect 15276 25687 15278 25707
rect 15420 25687 15422 25707
rect 15492 25687 15494 25707
rect 15540 25687 15542 25707
rect 15636 25687 15638 25707
rect 15660 25687 15662 25707
rect 15708 25687 15710 25707
rect 15732 25687 15734 25707
rect 15756 25687 15758 25707
rect 15804 25687 15806 25707
rect 15828 25687 15830 25707
rect 15852 25687 15854 25707
rect 15900 25687 15902 25707
rect 15948 25687 15950 25707
rect 15985 25702 15988 25707
rect 15996 25702 15998 25707
rect 15995 25688 15998 25702
rect 16044 25687 16046 25707
rect 16068 25687 16071 25704
rect 16164 25687 16166 25707
rect 16260 25687 16262 25707
rect 16308 25687 16310 25707
rect 16332 25687 16334 25707
rect 16356 25687 16358 25707
rect 16404 25687 16406 25707
rect 16452 25687 16454 25707
rect 16548 25687 16550 25707
rect 16572 25687 16574 25707
rect 16620 25687 16622 25707
rect 16668 25687 16670 25707
rect 16716 25687 16718 25707
rect 16764 25687 16766 25707
rect 16812 25687 16814 25707
rect 16884 25687 16886 25707
rect 16908 25687 16910 25707
rect 16980 25687 16982 25707
rect 17052 25687 17054 25707
rect 17196 25687 17198 25707
rect 17220 25687 17222 25707
rect 17292 25687 17294 25707
rect 17316 25687 17318 25707
rect 18084 25687 18086 25707
rect 18132 25687 18134 25707
rect 18228 25687 18230 25707
rect 18396 25687 18398 25707
rect 18492 25687 18494 25707
rect 18516 25687 18518 25707
rect 18564 25687 18566 25707
rect 18612 25687 18614 25707
rect 18660 25687 18662 25707
rect 18708 25687 18710 25707
rect 18756 25687 18758 25707
rect 18804 25687 18806 25707
rect 18852 25687 18854 25707
rect 18900 25687 18902 25707
rect 18996 25687 18998 25707
rect 19020 25687 19022 25707
rect 19092 25687 19094 25707
rect 19116 25687 19118 25707
rect 19140 25687 19142 25707
rect 19188 25687 19190 25707
rect 19236 25687 19238 25707
rect 19332 25687 19334 25707
rect 19476 25687 19478 25707
rect 19788 25687 19790 25707
rect 19836 25687 19838 25707
rect 19860 25687 19862 25707
rect 19884 25687 19886 25707
rect 19932 25687 19934 25707
rect 19956 25687 19958 25707
rect 19980 25687 19982 25707
rect 20028 25687 20030 25707
rect 20052 25687 20054 25707
rect 20076 25687 20078 25707
rect 20148 25687 20150 25707
rect 20172 25687 20174 25707
rect 20196 25687 20198 25707
rect 20268 25687 20270 25707
rect 20292 25687 20294 25707
rect 20388 25687 20390 25707
rect 20412 25687 20414 25707
rect 20508 25687 20510 25707
rect 20556 25687 20558 25707
rect 20604 25687 20606 25707
rect 20916 25687 20918 25707
rect 20964 25687 20966 25707
rect 21012 25687 21014 25707
rect 21060 25687 21062 25707
rect 21108 25687 21110 25707
rect 21204 25687 21206 25707
rect 21300 25687 21302 25707
rect 21324 25687 21326 25707
rect 21444 25687 21446 25707
rect 21468 25687 21470 25707
rect 21564 25687 21566 25707
rect 21567 25704 21581 25707
rect 21588 25707 24149 25711
rect 21588 25704 21605 25707
rect 21612 25704 21615 25707
rect 21588 25687 21590 25704
rect 21684 25687 21686 25707
rect 21708 25687 21710 25707
rect 21828 25687 21830 25707
rect 21924 25687 21926 25707
rect 22068 25687 22070 25707
rect 22188 25687 22190 25707
rect 22212 25687 22214 25707
rect 22884 25687 22886 25707
rect 22980 25687 22982 25707
rect 23076 25687 23078 25707
rect 23100 25687 23102 25707
rect 23124 25687 23126 25707
rect 23244 25687 23246 25707
rect 23340 25687 23342 25707
rect 23412 25687 23414 25707
rect 23508 25687 23510 25707
rect 23556 25687 23558 25707
rect 23652 25687 23654 25707
rect 23676 25687 23678 25707
rect 23724 25687 23726 25707
rect 23772 25687 23774 25707
rect 23820 25687 23822 25707
rect 23916 25687 23918 25707
rect 24012 25687 24014 25707
rect 24060 25687 24062 25707
rect 24135 25704 24149 25707
rect 24156 25707 27323 25711
rect 24156 25704 24173 25707
rect 24396 25704 24398 25707
rect 24156 25687 24158 25704
rect 24396 25687 24399 25704
rect 24492 25687 24494 25707
rect 24516 25687 24518 25707
rect 24588 25687 24590 25707
rect 24612 25687 24614 25707
rect 24684 25687 24686 25707
rect 24732 25687 24734 25707
rect 24756 25687 24758 25707
rect 24780 25687 24782 25707
rect 24852 25687 24854 25707
rect 24876 25687 24878 25707
rect 24972 25687 24974 25707
rect 24985 25702 24988 25707
rect 24996 25702 24998 25707
rect 24995 25688 24998 25702
rect 25068 25687 25070 25707
rect 25164 25687 25166 25707
rect 25260 25687 25262 25707
rect 25284 25687 25286 25707
rect 25356 25687 25358 25707
rect 25380 25687 25382 25707
rect 25404 25687 25406 25707
rect 25500 25687 25502 25707
rect 25596 25687 25598 25707
rect 27036 25687 27038 25707
rect 27108 25688 27110 25707
rect 27097 25687 27131 25688
rect -16377 25683 -13099 25687
rect -16377 25680 -16363 25683
rect -16356 25680 -16353 25683
rect -16308 25680 -16306 25683
rect -16284 25680 -16282 25683
rect -16308 25663 -16305 25680
rect -16284 25663 -16281 25680
rect -16260 25663 -16258 25683
rect -15324 25663 -15322 25683
rect -15108 25663 -15106 25683
rect -14903 25663 -14845 25664
rect -14772 25663 -14770 25683
rect -14687 25678 -14684 25683
rect -14677 25664 -14674 25678
rect -14676 25663 -14674 25664
rect -14567 25663 -14509 25664
rect -14436 25663 -14434 25683
rect -14340 25663 -14338 25683
rect -13932 25663 -13930 25683
rect -13788 25663 -13786 25683
rect -13572 25663 -13570 25683
rect -13356 25663 -13354 25683
rect -13113 25680 -13099 25683
rect -13089 25683 -9355 25687
rect -13089 25680 -13075 25683
rect -13068 25680 -13065 25683
rect -12887 25663 -12853 25664
rect -12780 25663 -12778 25683
rect -12756 25663 -12754 25683
rect -12660 25663 -12658 25683
rect -12564 25663 -12562 25683
rect -12492 25663 -12490 25683
rect -12396 25663 -12394 25683
rect -12348 25663 -12346 25683
rect -12252 25663 -12250 25683
rect -12156 25663 -12154 25683
rect -12060 25663 -12058 25683
rect -11844 25663 -11842 25683
rect -11676 25663 -11674 25683
rect -11556 25663 -11554 25683
rect -11508 25663 -11506 25683
rect -11436 25663 -11434 25683
rect -11412 25663 -11410 25683
rect -11340 25663 -11338 25683
rect -11196 25663 -11194 25683
rect -11124 25664 -11122 25683
rect -11135 25663 -11101 25664
rect -11100 25663 -11098 25683
rect -11028 25664 -11026 25683
rect -11039 25663 -11005 25664
rect -10740 25663 -10738 25683
rect -10668 25663 -10666 25683
rect -10644 25663 -10642 25683
rect -9996 25663 -9994 25683
rect -9911 25678 -9908 25683
rect -9901 25664 -9898 25678
rect -9900 25663 -9898 25664
rect -9828 25663 -9826 25683
rect -9732 25663 -9730 25683
rect -9516 25663 -9514 25683
rect -9468 25663 -9466 25683
rect -9369 25680 -9355 25683
rect -9348 25683 -787 25687
rect -9348 25680 -9331 25683
rect -9348 25663 -9346 25680
rect -9180 25663 -9178 25683
rect -8604 25663 -8602 25683
rect -8484 25663 -8482 25683
rect -8436 25663 -8434 25683
rect -8388 25663 -8386 25683
rect -8364 25663 -8362 25683
rect -8340 25663 -8338 25683
rect -8268 25663 -8266 25683
rect -8100 25663 -8098 25683
rect -8052 25663 -8050 25683
rect -8015 25678 -8012 25683
rect -8005 25664 -8002 25678
rect -8004 25663 -8002 25664
rect -7932 25663 -7930 25683
rect -7692 25663 -7690 25683
rect -7620 25663 -7618 25683
rect -7524 25663 -7522 25683
rect -7356 25663 -7354 25683
rect -7308 25663 -7306 25683
rect -7212 25663 -7210 25683
rect -7116 25663 -7114 25683
rect -7068 25663 -7066 25683
rect -6972 25663 -6970 25683
rect -6948 25663 -6946 25683
rect -6876 25663 -6874 25683
rect -6852 25663 -6850 25683
rect -6780 25663 -6778 25683
rect -6756 25663 -6754 25683
rect -6660 25663 -6658 25683
rect -6612 25663 -6610 25683
rect -6516 25663 -6514 25683
rect -6372 25663 -6370 25683
rect -6156 25663 -6154 25683
rect -6060 25663 -6058 25683
rect -6036 25663 -6034 25683
rect -5892 25663 -5890 25683
rect -5652 25664 -5650 25683
rect -5687 25663 -5629 25664
rect -5268 25663 -5266 25683
rect -5196 25663 -5194 25683
rect -5172 25663 -5170 25683
rect -5100 25663 -5098 25683
rect -5076 25663 -5074 25683
rect -4980 25663 -4978 25683
rect -4956 25663 -4954 25683
rect -4943 25663 -4885 25664
rect -4860 25663 -4858 25683
rect -4644 25663 -4642 25683
rect -4548 25663 -4546 25683
rect -4500 25663 -4498 25683
rect -4404 25663 -4402 25683
rect -4308 25663 -4306 25683
rect -4260 25663 -4258 25683
rect -4164 25663 -4162 25683
rect -4020 25663 -4018 25683
rect -3876 25663 -3874 25683
rect -3732 25663 -3730 25683
rect -3588 25663 -3586 25683
rect -3564 25663 -3562 25683
rect -3516 25663 -3514 25683
rect -3492 25663 -3490 25683
rect -3468 25663 -3466 25683
rect -3420 25663 -3418 25683
rect -3324 25663 -3322 25683
rect -3228 25663 -3226 25683
rect -3132 25663 -3130 25683
rect -3012 25663 -3010 25683
rect -2964 25663 -2962 25683
rect -2916 25663 -2914 25683
rect -2892 25663 -2890 25683
rect -2868 25663 -2866 25683
rect -2820 25663 -2818 25683
rect -2796 25663 -2794 25683
rect -2772 25663 -2770 25683
rect -2676 25663 -2674 25683
rect -2580 25663 -2578 25683
rect -2364 25663 -2362 25683
rect -2316 25663 -2314 25683
rect -2268 25663 -2266 25683
rect -2244 25663 -2242 25683
rect -2172 25663 -2170 25683
rect -2148 25663 -2146 25683
rect -2076 25663 -2074 25683
rect -2052 25663 -2050 25683
rect -1980 25663 -1978 25683
rect -1884 25663 -1882 25683
rect -1572 25663 -1570 25683
rect -1476 25663 -1474 25683
rect -1380 25663 -1378 25683
rect -1356 25663 -1354 25683
rect -1308 25663 -1306 25683
rect -1260 25663 -1258 25683
rect -1140 25663 -1138 25683
rect -801 25680 -787 25683
rect -777 25683 2333 25687
rect -777 25680 -763 25683
rect -756 25680 -753 25683
rect -708 25663 -706 25683
rect -612 25663 -610 25683
rect -588 25663 -586 25683
rect -540 25663 -538 25683
rect -492 25663 -490 25683
rect -444 25663 -442 25683
rect -396 25663 -394 25683
rect -300 25663 -298 25683
rect -276 25663 -274 25683
rect -228 25663 -226 25683
rect -12 25663 -10 25683
rect 156 25663 158 25683
rect 204 25663 206 25683
rect 252 25663 254 25683
rect 348 25663 350 25683
rect 468 25663 470 25683
rect 492 25663 494 25683
rect 564 25663 566 25683
rect 588 25663 590 25683
rect 636 25663 638 25683
rect 660 25663 662 25683
rect 732 25663 734 25683
rect 1092 25663 1094 25683
rect 1308 25663 1310 25683
rect 1332 25663 1334 25683
rect 1380 25663 1382 25683
rect 1428 25663 1430 25683
rect 1476 25663 1478 25683
rect 1644 25663 1646 25683
rect 1692 25663 1694 25683
rect 1740 25663 1742 25683
rect 1788 25663 1790 25683
rect 2028 25663 2030 25683
rect 2076 25663 2078 25683
rect 2100 25663 2102 25683
rect 2124 25663 2126 25683
rect 2172 25663 2174 25683
rect 2220 25663 2222 25683
rect 2316 25663 2318 25683
rect 2319 25680 2333 25683
rect 2343 25683 7157 25687
rect 2343 25680 2357 25683
rect 2364 25680 2367 25683
rect 2412 25663 2414 25683
rect 2460 25663 2462 25683
rect 2508 25663 2510 25683
rect 2580 25663 2582 25683
rect 2604 25663 2606 25683
rect 2676 25663 2678 25683
rect 2700 25663 2702 25683
rect 2748 25663 2750 25683
rect 2772 25663 2774 25683
rect 2796 25663 2798 25683
rect 2844 25663 2846 25683
rect 2868 25663 2870 25683
rect 2892 25663 2894 25683
rect 2940 25663 2942 25683
rect 3012 25663 3014 25683
rect 3108 25663 3110 25683
rect 3135 25680 3149 25683
rect 3156 25680 3159 25683
rect 3252 25663 3254 25683
rect 3348 25663 3350 25683
rect 3396 25663 3398 25683
rect 3564 25663 3566 25683
rect 3636 25663 3638 25683
rect 3660 25663 3662 25683
rect 3732 25663 3734 25683
rect 3828 25663 3830 25683
rect 3924 25663 3926 25683
rect 4020 25663 4022 25683
rect 4044 25663 4046 25683
rect 4092 25663 4094 25683
rect 4116 25663 4118 25683
rect 4140 25663 4142 25683
rect 4188 25663 4190 25683
rect 4212 25663 4214 25683
rect 4236 25663 4238 25683
rect 4308 25663 4310 25683
rect 4332 25663 4334 25683
rect 4404 25663 4406 25683
rect 4500 25663 4502 25683
rect 4596 25663 4598 25683
rect 4692 25663 4694 25683
rect 4860 25663 4862 25683
rect 4956 25663 4958 25683
rect 4980 25663 4982 25683
rect 5004 25663 5006 25683
rect 5052 25663 5054 25683
rect 5100 25663 5102 25683
rect 5124 25663 5126 25683
rect 5220 25663 5222 25683
rect 5268 25663 5270 25683
rect 5388 25663 5390 25683
rect 5484 25663 5486 25683
rect 5508 25663 5510 25683
rect 5532 25663 5534 25683
rect 5628 25663 5630 25683
rect 5652 25663 5654 25683
rect 5748 25663 5750 25683
rect 5796 25663 5798 25683
rect 5844 25663 5846 25683
rect 5892 25663 5894 25683
rect 6132 25663 6134 25683
rect 6180 25663 6182 25683
rect 6228 25663 6230 25683
rect 6252 25663 6254 25683
rect 6276 25663 6278 25683
rect 6324 25663 6326 25683
rect 6372 25663 6374 25683
rect 6492 25663 6494 25683
rect 6588 25663 6590 25683
rect 6612 25663 6614 25683
rect 6660 25663 6662 25683
rect 6684 25663 6686 25683
rect 6708 25663 6710 25683
rect 6780 25663 6782 25683
rect 6804 25663 6806 25683
rect 6900 25663 6902 25683
rect 6924 25663 6926 25683
rect 7020 25663 7022 25683
rect 7068 25663 7070 25683
rect 7119 25680 7133 25683
rect 7140 25680 7157 25683
rect 7164 25683 16061 25687
rect 7164 25680 7181 25683
rect 7164 25663 7166 25680
rect 7236 25663 7238 25683
rect 7332 25663 7334 25683
rect 7380 25663 7382 25683
rect 7428 25663 7430 25683
rect 7452 25663 7454 25683
rect 7476 25663 7478 25683
rect 7524 25663 7526 25683
rect 7548 25663 7550 25683
rect 7572 25663 7574 25683
rect 7620 25663 7622 25683
rect 7644 25663 7646 25683
rect 7668 25663 7670 25683
rect 7788 25663 7790 25683
rect 7884 25663 7886 25683
rect 7956 25663 7958 25683
rect 7980 25663 7982 25683
rect 8028 25663 8030 25683
rect 8196 25663 8198 25683
rect 8244 25663 8246 25683
rect 8268 25663 8270 25683
rect 8292 25663 8294 25683
rect 8340 25663 8342 25683
rect 8364 25663 8366 25683
rect 8388 25663 8390 25683
rect 8436 25663 8438 25683
rect 8604 25663 8606 25683
rect 8652 25663 8654 25683
rect 8700 25663 8702 25683
rect 8724 25663 8726 25683
rect 8748 25663 8750 25683
rect 8820 25663 8822 25683
rect 8844 25663 8846 25683
rect 8868 25663 8870 25683
rect 9516 25663 9518 25683
rect 9612 25663 9614 25683
rect 9660 25663 9662 25683
rect 9684 25663 9686 25683
rect 9708 25663 9710 25683
rect 9756 25663 9758 25683
rect 9780 25663 9782 25683
rect 9804 25663 9806 25683
rect 9852 25663 9854 25683
rect 9900 25663 9902 25683
rect 9948 25663 9950 25683
rect 9996 25663 9998 25683
rect 10068 25663 10070 25683
rect 10092 25663 10094 25683
rect 10116 25663 10118 25683
rect 10164 25663 10166 25683
rect 10188 25663 10190 25683
rect 10212 25663 10214 25683
rect 10284 25663 10286 25683
rect 10308 25663 10310 25683
rect 10332 25663 10334 25683
rect 10380 25663 10382 25683
rect 10404 25663 10406 25683
rect 10428 25663 10430 25683
rect 10476 25663 10478 25683
rect 10500 25663 10502 25683
rect 10524 25663 10526 25683
rect 10572 25663 10574 25683
rect 10596 25663 10598 25683
rect 10620 25663 10622 25683
rect 10668 25663 10670 25683
rect 10692 25663 10694 25683
rect 10716 25663 10718 25683
rect 10788 25663 10790 25683
rect 10836 25663 10838 25683
rect 10956 25663 10958 25683
rect 11004 25663 11006 25683
rect 11052 25663 11054 25683
rect 11076 25680 11078 25683
rect 11076 25663 11079 25680
rect 11100 25663 11102 25683
rect 11172 25663 11174 25683
rect 11220 25663 11222 25683
rect 11340 25663 11342 25683
rect 11436 25663 11438 25683
rect 11532 25663 11534 25683
rect 11580 25663 11582 25683
rect 11628 25663 11630 25683
rect 11676 25663 11678 25683
rect 11724 25663 11726 25683
rect 11772 25663 11774 25683
rect 11796 25663 11798 25683
rect 11892 25663 11894 25683
rect 11988 25663 11990 25683
rect 12060 25663 12062 25683
rect 12132 25663 12134 25683
rect 12228 25663 12230 25683
rect 12276 25663 12278 25683
rect 12324 25663 12326 25683
rect 12420 25663 12422 25683
rect 12444 25663 12446 25683
rect 12492 25663 12494 25683
rect 12516 25663 12518 25683
rect 12540 25663 12542 25683
rect 12588 25663 12590 25683
rect 12636 25663 12638 25683
rect 12732 25663 12734 25683
rect 12756 25663 12758 25683
rect 12804 25663 12806 25683
rect 12828 25663 12830 25683
rect 12852 25663 12854 25683
rect 12948 25663 12950 25683
rect 12972 25663 12974 25683
rect 13044 25663 13046 25683
rect 13068 25663 13070 25683
rect 13116 25663 13118 25683
rect 13284 25663 13286 25683
rect 13332 25663 13334 25683
rect 13572 25663 13574 25683
rect 13620 25663 13622 25683
rect 13668 25663 13670 25683
rect 13716 25663 13718 25683
rect 13764 25663 13766 25683
rect 13860 25663 13862 25683
rect 13887 25680 13901 25683
rect 13908 25680 13911 25683
rect 13956 25663 13958 25683
rect 14004 25663 14006 25683
rect 14100 25663 14102 25683
rect 14196 25663 14198 25683
rect 14292 25663 14294 25683
rect 15180 25663 15182 25683
rect 15276 25663 15278 25683
rect 15327 25680 15341 25683
rect 15420 25663 15422 25683
rect 15492 25663 15494 25683
rect 15540 25664 15542 25683
rect 15529 25663 15563 25664
rect 15636 25663 15638 25683
rect 15660 25663 15662 25683
rect 15708 25663 15710 25683
rect 15732 25663 15734 25683
rect 15756 25663 15758 25683
rect 15804 25663 15806 25683
rect 15828 25663 15830 25683
rect 15852 25663 15854 25683
rect 15900 25663 15902 25683
rect 15948 25663 15950 25683
rect 16044 25663 16046 25683
rect 16047 25680 16061 25683
rect 16068 25683 27131 25687
rect 27145 25687 27179 25688
rect 27217 25687 27251 25688
rect 27145 25683 27251 25687
rect 16068 25680 16085 25683
rect 16068 25663 16070 25680
rect 16164 25663 16166 25683
rect 16260 25663 16262 25683
rect 16308 25663 16310 25683
rect 16332 25663 16334 25683
rect 16356 25663 16358 25683
rect 16404 25663 16406 25683
rect 16452 25663 16454 25683
rect 16548 25663 16550 25683
rect 16572 25663 16574 25683
rect 16620 25663 16622 25683
rect 16668 25663 16670 25683
rect 16716 25663 16718 25683
rect 16764 25663 16766 25683
rect 16812 25663 16814 25683
rect 16884 25663 16886 25683
rect 16908 25663 16910 25683
rect 16980 25663 16982 25683
rect 17052 25663 17054 25683
rect 17196 25663 17198 25683
rect 17220 25663 17222 25683
rect 17292 25663 17294 25683
rect 17316 25663 17318 25683
rect 18084 25663 18086 25683
rect 18132 25663 18134 25683
rect 18228 25663 18230 25683
rect 18396 25663 18398 25683
rect 18492 25663 18494 25683
rect 18516 25663 18518 25683
rect 18564 25663 18566 25683
rect 18612 25663 18614 25683
rect 18660 25663 18662 25683
rect 18708 25663 18710 25683
rect 18756 25663 18758 25683
rect 18804 25663 18806 25683
rect 18852 25663 18854 25683
rect 18900 25663 18902 25683
rect 18996 25663 18998 25683
rect 19020 25663 19022 25683
rect 19092 25663 19094 25683
rect 19116 25663 19118 25683
rect 19140 25663 19142 25683
rect 19188 25663 19190 25683
rect 19236 25663 19238 25683
rect 19332 25663 19334 25683
rect 19441 25663 19475 25664
rect 19476 25663 19478 25683
rect 19788 25663 19790 25683
rect 19836 25663 19838 25683
rect 19860 25663 19862 25683
rect 19884 25663 19886 25683
rect 19932 25663 19934 25683
rect 19956 25663 19958 25683
rect 19980 25663 19982 25683
rect 20028 25663 20030 25683
rect 20052 25663 20054 25683
rect 20076 25663 20078 25683
rect 20148 25663 20150 25683
rect 20172 25663 20174 25683
rect 20196 25663 20198 25683
rect 20268 25663 20270 25683
rect 20292 25663 20294 25683
rect 20388 25663 20390 25683
rect 20412 25663 20414 25683
rect 20508 25663 20510 25683
rect 20556 25663 20558 25683
rect 20604 25663 20606 25683
rect 20916 25663 20918 25683
rect 20964 25663 20966 25683
rect 21012 25663 21014 25683
rect 21060 25663 21062 25683
rect 21108 25663 21110 25683
rect 21204 25663 21206 25683
rect 21300 25663 21302 25683
rect 21324 25663 21326 25683
rect 21444 25663 21446 25683
rect 21468 25663 21470 25683
rect 21564 25663 21566 25683
rect 21588 25663 21590 25683
rect 21684 25663 21686 25683
rect 21708 25663 21710 25683
rect 21828 25663 21830 25683
rect 21924 25663 21926 25683
rect 22068 25663 22070 25683
rect 22188 25663 22190 25683
rect 22212 25663 22214 25683
rect 22884 25663 22886 25683
rect 22980 25663 22982 25683
rect 23076 25663 23078 25683
rect 23100 25663 23102 25683
rect 23124 25663 23126 25683
rect 23244 25663 23246 25683
rect 23340 25663 23342 25683
rect 23412 25663 23414 25683
rect 23508 25663 23510 25683
rect 23556 25663 23558 25683
rect 23593 25663 23651 25664
rect 23652 25663 23654 25683
rect 23676 25663 23678 25683
rect 23724 25663 23726 25683
rect 23772 25663 23774 25683
rect 23820 25663 23822 25683
rect 23916 25663 23918 25683
rect 24012 25663 24014 25683
rect 24060 25663 24062 25683
rect 24156 25663 24158 25683
rect 24375 25680 24389 25683
rect 24396 25680 24399 25683
rect 24492 25663 24494 25683
rect 24516 25663 24518 25683
rect 24588 25663 24590 25683
rect 24612 25663 24614 25683
rect 24684 25663 24686 25683
rect 24732 25663 24734 25683
rect 24756 25663 24758 25683
rect 24780 25663 24782 25683
rect 24852 25663 24854 25683
rect 24876 25663 24878 25683
rect 24972 25663 24974 25683
rect 25068 25663 25070 25683
rect 25071 25680 25085 25683
rect 25164 25663 25166 25683
rect 25260 25663 25262 25683
rect 25284 25663 25286 25683
rect 25356 25663 25358 25683
rect 25380 25663 25382 25683
rect 25404 25663 25406 25683
rect 25500 25663 25502 25683
rect 25596 25663 25598 25683
rect 27036 25664 27038 25683
rect 27097 25678 27100 25683
rect 27108 25678 27110 25683
rect 27107 25664 27110 25678
rect 27241 25670 27245 25678
rect 27231 25664 27241 25670
rect 26809 25663 26843 25664
rect -16329 25656 -16326 25663
rect -16316 25656 -16315 25663
rect -16308 25659 -14587 25663
rect -16308 25656 -16291 25659
rect -16284 25656 -16281 25659
rect -16260 25639 -16258 25659
rect -15324 25639 -15322 25659
rect -15108 25639 -15106 25659
rect -14903 25654 -14900 25659
rect -14772 25656 -14770 25659
rect -14721 25656 -14707 25659
rect -14893 25640 -14890 25654
rect -14892 25639 -14890 25640
rect -14772 25639 -14769 25656
rect -14676 25639 -14674 25659
rect -14601 25656 -14587 25659
rect -14577 25659 -9811 25663
rect -14577 25656 -14563 25659
rect -14436 25656 -14434 25659
rect -14436 25639 -14433 25656
rect -14340 25639 -14338 25659
rect -13932 25640 -13930 25659
rect -14039 25639 -14005 25640
rect -13943 25639 -13909 25640
rect -13788 25639 -13786 25659
rect -13572 25640 -13570 25659
rect -13356 25640 -13354 25659
rect -12780 25656 -12778 25659
rect -13583 25639 -13549 25640
rect -13367 25639 -13333 25640
rect -12780 25639 -12777 25656
rect -12756 25639 -12754 25659
rect -12660 25639 -12658 25659
rect -12564 25640 -12562 25659
rect -12575 25639 -12541 25640
rect -12492 25639 -12490 25659
rect -12396 25639 -12394 25659
rect -12348 25639 -12346 25659
rect -12252 25639 -12250 25659
rect -12156 25639 -12154 25659
rect -12060 25639 -12058 25659
rect -11844 25639 -11842 25659
rect -11676 25639 -11674 25659
rect -11556 25640 -11554 25659
rect -11567 25639 -11533 25640
rect -11508 25639 -11506 25659
rect -11436 25639 -11434 25659
rect -11412 25639 -11410 25659
rect -11375 25639 -11341 25640
rect -11340 25639 -11338 25659
rect -11196 25639 -11194 25659
rect -11135 25654 -11132 25659
rect -11124 25654 -11122 25659
rect -11125 25640 -11122 25654
rect -11100 25639 -11098 25659
rect -11039 25654 -11036 25659
rect -11028 25656 -11026 25659
rect -11028 25654 -11025 25656
rect -11029 25640 -11025 25654
rect -10740 25639 -10738 25659
rect -10668 25640 -10666 25659
rect -10679 25639 -10645 25640
rect -10644 25639 -10642 25659
rect -10535 25639 -10477 25640
rect -9996 25639 -9994 25659
rect -9900 25639 -9898 25659
rect -9828 25639 -9826 25659
rect -9825 25656 -9811 25659
rect -9801 25659 -7915 25663
rect -9801 25656 -9787 25659
rect -9732 25639 -9730 25659
rect -9516 25639 -9514 25659
rect -9468 25639 -9466 25659
rect -9348 25639 -9346 25659
rect -9180 25639 -9178 25659
rect -8604 25639 -8602 25659
rect -8484 25639 -8482 25659
rect -8436 25639 -8434 25659
rect -8388 25639 -8386 25659
rect -8364 25639 -8362 25659
rect -8340 25639 -8338 25659
rect -8268 25639 -8266 25659
rect -8100 25639 -8098 25659
rect -8052 25639 -8050 25659
rect -8004 25639 -8002 25659
rect -7932 25639 -7930 25659
rect -7929 25656 -7915 25659
rect -7905 25659 26843 25663
rect 26929 25663 26963 25664
rect 27001 25663 27059 25664
rect 27073 25663 27107 25664
rect 26929 25659 27107 25663
rect -7905 25656 -7891 25659
rect -7692 25639 -7690 25659
rect -7620 25639 -7618 25659
rect -7524 25639 -7522 25659
rect -7356 25639 -7354 25659
rect -7308 25639 -7306 25659
rect -7212 25639 -7210 25659
rect -7199 25639 -7141 25640
rect -7116 25639 -7114 25659
rect -7068 25639 -7066 25659
rect -6972 25639 -6970 25659
rect -6948 25639 -6946 25659
rect -6876 25639 -6874 25659
rect -6852 25639 -6850 25659
rect -6780 25639 -6778 25659
rect -6756 25639 -6754 25659
rect -6660 25639 -6658 25659
rect -6612 25639 -6610 25659
rect -6516 25639 -6514 25659
rect -6372 25639 -6370 25659
rect -6156 25639 -6154 25659
rect -6060 25639 -6058 25659
rect -6036 25639 -6034 25659
rect -5892 25639 -5890 25659
rect -5663 25654 -5660 25659
rect -5652 25654 -5650 25659
rect -5653 25640 -5650 25654
rect -5268 25639 -5266 25659
rect -5196 25639 -5194 25659
rect -5172 25639 -5170 25659
rect -5100 25639 -5098 25659
rect -5076 25639 -5074 25659
rect -4980 25639 -4978 25659
rect -4956 25639 -4954 25659
rect -4860 25639 -4858 25659
rect -4644 25639 -4642 25659
rect -4548 25639 -4546 25659
rect -4500 25639 -4498 25659
rect -4404 25639 -4402 25659
rect -4308 25639 -4306 25659
rect -4260 25639 -4258 25659
rect -4164 25639 -4162 25659
rect -4020 25639 -4018 25659
rect -3876 25639 -3874 25659
rect -3732 25639 -3730 25659
rect -3588 25639 -3586 25659
rect -3564 25639 -3562 25659
rect -3516 25639 -3514 25659
rect -3492 25639 -3490 25659
rect -3468 25639 -3466 25659
rect -3420 25639 -3418 25659
rect -3324 25639 -3322 25659
rect -3228 25639 -3226 25659
rect -3132 25639 -3130 25659
rect -3012 25639 -3010 25659
rect -2964 25639 -2962 25659
rect -2916 25639 -2914 25659
rect -2892 25639 -2890 25659
rect -2868 25639 -2866 25659
rect -2820 25639 -2818 25659
rect -2796 25639 -2794 25659
rect -2772 25639 -2770 25659
rect -2676 25639 -2674 25659
rect -2580 25639 -2578 25659
rect -2364 25639 -2362 25659
rect -2316 25639 -2314 25659
rect -2268 25639 -2266 25659
rect -2244 25639 -2242 25659
rect -2172 25639 -2170 25659
rect -2148 25639 -2146 25659
rect -2076 25639 -2074 25659
rect -2052 25639 -2050 25659
rect -1980 25639 -1978 25659
rect -1884 25639 -1882 25659
rect -1572 25639 -1570 25659
rect -1476 25639 -1474 25659
rect -1380 25639 -1378 25659
rect -1356 25639 -1354 25659
rect -1308 25639 -1306 25659
rect -1260 25639 -1258 25659
rect -1140 25639 -1138 25659
rect -708 25639 -706 25659
rect -612 25639 -610 25659
rect -588 25639 -586 25659
rect -540 25639 -538 25659
rect -492 25639 -490 25659
rect -444 25639 -442 25659
rect -396 25639 -394 25659
rect -300 25639 -298 25659
rect -276 25639 -274 25659
rect -228 25639 -226 25659
rect -12 25639 -10 25659
rect 156 25639 158 25659
rect 204 25639 206 25659
rect 252 25639 254 25659
rect 348 25639 350 25659
rect 468 25639 470 25659
rect 492 25639 494 25659
rect 564 25639 566 25659
rect 588 25639 590 25659
rect 636 25639 638 25659
rect 660 25639 662 25659
rect 732 25639 734 25659
rect 1092 25639 1094 25659
rect 1308 25639 1310 25659
rect 1332 25639 1334 25659
rect 1380 25639 1382 25659
rect 1428 25639 1430 25659
rect 1476 25639 1478 25659
rect 1644 25639 1646 25659
rect 1692 25639 1694 25659
rect 1740 25639 1742 25659
rect 1788 25639 1790 25659
rect 2028 25639 2030 25659
rect 2076 25639 2078 25659
rect 2100 25639 2102 25659
rect 2124 25639 2126 25659
rect 2172 25639 2174 25659
rect 2220 25639 2222 25659
rect 2316 25639 2318 25659
rect 2412 25639 2414 25659
rect 2460 25639 2462 25659
rect 2508 25639 2510 25659
rect 2580 25639 2582 25659
rect 2604 25639 2606 25659
rect 2676 25639 2678 25659
rect 2700 25639 2702 25659
rect 2748 25639 2750 25659
rect 2772 25639 2774 25659
rect 2796 25639 2798 25659
rect 2844 25639 2846 25659
rect 2868 25639 2870 25659
rect 2892 25639 2894 25659
rect 2940 25639 2942 25659
rect 3012 25639 3014 25659
rect 3108 25639 3110 25659
rect 3252 25639 3254 25659
rect 3348 25639 3350 25659
rect 3396 25639 3398 25659
rect 3564 25639 3566 25659
rect 3636 25639 3638 25659
rect 3660 25639 3662 25659
rect 3732 25639 3734 25659
rect 3828 25639 3830 25659
rect 3924 25639 3926 25659
rect 4020 25639 4022 25659
rect 4044 25639 4046 25659
rect 4092 25639 4094 25659
rect 4116 25639 4118 25659
rect 4140 25639 4142 25659
rect 4188 25639 4190 25659
rect 4212 25639 4214 25659
rect 4236 25639 4238 25659
rect 4308 25639 4310 25659
rect 4332 25639 4334 25659
rect 4404 25639 4406 25659
rect 4500 25639 4502 25659
rect 4596 25639 4598 25659
rect 4692 25639 4694 25659
rect 4860 25639 4862 25659
rect 4956 25639 4958 25659
rect 4980 25639 4982 25659
rect 5004 25639 5006 25659
rect 5052 25639 5054 25659
rect 5100 25639 5102 25659
rect 5124 25639 5126 25659
rect 5220 25639 5222 25659
rect 5268 25639 5270 25659
rect 5388 25639 5390 25659
rect 5484 25639 5486 25659
rect 5508 25639 5510 25659
rect 5532 25639 5534 25659
rect 5628 25639 5630 25659
rect 5652 25639 5654 25659
rect 5748 25639 5750 25659
rect 5796 25639 5798 25659
rect 5844 25639 5846 25659
rect 5892 25639 5894 25659
rect 6132 25639 6134 25659
rect 6180 25639 6182 25659
rect 6228 25639 6230 25659
rect 6252 25639 6254 25659
rect 6276 25639 6278 25659
rect 6324 25639 6326 25659
rect 6372 25639 6374 25659
rect 6492 25639 6494 25659
rect 6588 25639 6590 25659
rect 6612 25639 6614 25659
rect 6660 25639 6662 25659
rect 6684 25639 6686 25659
rect 6708 25639 6710 25659
rect 6780 25639 6782 25659
rect 6804 25639 6806 25659
rect 6900 25639 6902 25659
rect 6924 25639 6926 25659
rect 7020 25639 7022 25659
rect 7068 25639 7070 25659
rect 7164 25639 7166 25659
rect 7236 25639 7238 25659
rect 7332 25639 7334 25659
rect 7380 25639 7382 25659
rect 7428 25639 7430 25659
rect 7452 25639 7454 25659
rect 7476 25639 7478 25659
rect 7524 25639 7526 25659
rect 7548 25639 7550 25659
rect 7572 25639 7574 25659
rect 7620 25639 7622 25659
rect 7644 25639 7646 25659
rect 7668 25639 7670 25659
rect 7788 25639 7790 25659
rect 7884 25639 7886 25659
rect 7956 25639 7958 25659
rect 7980 25639 7982 25659
rect 8028 25639 8030 25659
rect 8196 25639 8198 25659
rect 8244 25639 8246 25659
rect 8268 25639 8270 25659
rect 8292 25639 8294 25659
rect 8340 25639 8342 25659
rect 8364 25639 8366 25659
rect 8388 25639 8390 25659
rect 8436 25639 8438 25659
rect 8604 25639 8606 25659
rect 8652 25639 8654 25659
rect 8700 25639 8702 25659
rect 8724 25639 8726 25659
rect 8748 25639 8750 25659
rect 8820 25639 8822 25659
rect 8844 25639 8846 25659
rect 8868 25639 8870 25659
rect 9516 25639 9518 25659
rect 9612 25639 9614 25659
rect 9660 25639 9662 25659
rect 9684 25639 9686 25659
rect 9708 25639 9710 25659
rect 9756 25639 9758 25659
rect 9780 25639 9782 25659
rect 9804 25639 9806 25659
rect 9852 25639 9854 25659
rect 9900 25639 9902 25659
rect 9948 25639 9950 25659
rect 9996 25639 9998 25659
rect 10068 25639 10070 25659
rect 10092 25639 10094 25659
rect 10116 25639 10118 25659
rect 10164 25639 10166 25659
rect 10188 25639 10190 25659
rect 10212 25639 10214 25659
rect 10284 25639 10286 25659
rect 10308 25639 10310 25659
rect 10332 25639 10334 25659
rect 10380 25639 10382 25659
rect 10404 25639 10406 25659
rect 10428 25639 10430 25659
rect 10476 25639 10478 25659
rect 10500 25639 10502 25659
rect 10524 25639 10526 25659
rect 10572 25639 10574 25659
rect 10596 25639 10598 25659
rect 10620 25639 10622 25659
rect 10668 25639 10670 25659
rect 10692 25639 10694 25659
rect 10716 25639 10718 25659
rect 10788 25639 10790 25659
rect 10836 25639 10838 25659
rect 10956 25639 10958 25659
rect 11004 25639 11006 25659
rect 11052 25639 11054 25659
rect 11055 25656 11069 25659
rect 11076 25656 11079 25659
rect 11100 25639 11102 25659
rect 11172 25639 11174 25659
rect 11220 25639 11222 25659
rect 11340 25639 11342 25659
rect 11436 25639 11438 25659
rect 11532 25639 11534 25659
rect 11580 25639 11582 25659
rect 11628 25639 11630 25659
rect 11676 25639 11678 25659
rect 11724 25639 11726 25659
rect 11772 25639 11774 25659
rect 11796 25639 11798 25659
rect 11892 25639 11894 25659
rect 11988 25639 11990 25659
rect 12060 25639 12062 25659
rect 12132 25639 12134 25659
rect 12228 25639 12230 25659
rect 12276 25639 12278 25659
rect 12324 25639 12326 25659
rect 12420 25639 12422 25659
rect 12444 25639 12446 25659
rect 12492 25639 12494 25659
rect 12516 25639 12518 25659
rect 12540 25639 12542 25659
rect 12588 25639 12590 25659
rect 12636 25639 12638 25659
rect 12732 25639 12734 25659
rect 12756 25639 12758 25659
rect 12804 25639 12806 25659
rect 12828 25639 12830 25659
rect 12852 25639 12854 25659
rect 12948 25639 12950 25659
rect 12972 25639 12974 25659
rect 13044 25639 13046 25659
rect 13068 25639 13070 25659
rect 13116 25639 13118 25659
rect 13284 25639 13286 25659
rect 13332 25639 13334 25659
rect 13572 25639 13574 25659
rect 13620 25639 13622 25659
rect 13668 25639 13670 25659
rect 13716 25639 13718 25659
rect 13764 25639 13766 25659
rect 13860 25639 13862 25659
rect 13956 25639 13958 25659
rect 14004 25639 14006 25659
rect 14100 25639 14102 25659
rect 14196 25639 14198 25659
rect 14292 25639 14294 25659
rect 15180 25639 15182 25659
rect 15276 25639 15278 25659
rect 15420 25639 15422 25659
rect 15492 25639 15494 25659
rect 15529 25654 15532 25659
rect 15540 25654 15542 25659
rect 15539 25640 15542 25654
rect 15636 25656 15638 25659
rect 15636 25639 15639 25656
rect 15660 25639 15662 25659
rect 15708 25639 15710 25659
rect 15732 25639 15734 25659
rect 15756 25639 15758 25659
rect 15804 25639 15806 25659
rect 15828 25639 15830 25659
rect 15852 25639 15854 25659
rect 15900 25639 15902 25659
rect 15948 25639 15950 25659
rect 16044 25639 16046 25659
rect 16068 25639 16070 25659
rect 16164 25639 16166 25659
rect 16260 25639 16262 25659
rect 16308 25639 16310 25659
rect 16332 25639 16334 25659
rect 16356 25639 16358 25659
rect 16404 25639 16406 25659
rect 16452 25639 16454 25659
rect 16548 25639 16550 25659
rect 16572 25639 16574 25659
rect 16620 25639 16622 25659
rect 16668 25639 16670 25659
rect 16716 25639 16718 25659
rect 16764 25639 16766 25659
rect 16812 25639 16814 25659
rect 16884 25639 16886 25659
rect 16908 25639 16910 25659
rect 16980 25639 16982 25659
rect 17052 25639 17054 25659
rect 17196 25639 17198 25659
rect 17220 25639 17222 25659
rect 17292 25639 17294 25659
rect 17316 25639 17318 25659
rect 18084 25639 18086 25659
rect 18132 25639 18134 25659
rect 18228 25639 18230 25659
rect 18396 25639 18398 25659
rect 18492 25639 18494 25659
rect 18516 25639 18518 25659
rect 18564 25639 18566 25659
rect 18612 25639 18614 25659
rect 18660 25639 18662 25659
rect 18708 25639 18710 25659
rect 18756 25639 18758 25659
rect 18804 25639 18806 25659
rect 18852 25639 18854 25659
rect 18900 25639 18902 25659
rect 18996 25639 18998 25659
rect 19020 25639 19022 25659
rect 19092 25639 19094 25659
rect 19116 25639 19118 25659
rect 19140 25639 19142 25659
rect 19188 25639 19190 25659
rect 19236 25639 19238 25659
rect 19332 25639 19334 25659
rect 19476 25639 19478 25659
rect 19788 25639 19790 25659
rect 19836 25639 19838 25659
rect 19860 25639 19862 25659
rect 19884 25639 19886 25659
rect 19932 25639 19934 25659
rect 19956 25639 19958 25659
rect 19980 25639 19982 25659
rect 20028 25639 20030 25659
rect 20052 25639 20054 25659
rect 20076 25639 20078 25659
rect 20148 25639 20150 25659
rect 20172 25639 20174 25659
rect 20196 25639 20198 25659
rect 20268 25639 20270 25659
rect 20292 25639 20294 25659
rect 20388 25639 20390 25659
rect 20412 25639 20414 25659
rect 20508 25639 20510 25659
rect 20556 25639 20558 25659
rect 20604 25639 20606 25659
rect 20916 25639 20918 25659
rect 20964 25639 20966 25659
rect 21012 25639 21014 25659
rect 21060 25639 21062 25659
rect 21108 25639 21110 25659
rect 21204 25639 21206 25659
rect 21300 25639 21302 25659
rect 21324 25639 21326 25659
rect 21444 25639 21446 25659
rect 21468 25639 21470 25659
rect 21564 25639 21566 25659
rect 21588 25639 21590 25659
rect 21684 25639 21686 25659
rect 21708 25639 21710 25659
rect 21828 25639 21830 25659
rect 21924 25639 21926 25659
rect 22068 25639 22070 25659
rect 22188 25639 22190 25659
rect 22212 25639 22214 25659
rect 22884 25639 22886 25659
rect 22980 25639 22982 25659
rect 23076 25639 23078 25659
rect 23100 25639 23102 25659
rect 23124 25639 23126 25659
rect 23244 25639 23246 25659
rect 23340 25639 23342 25659
rect 23412 25639 23414 25659
rect 23508 25639 23510 25659
rect 23556 25639 23558 25659
rect 23593 25654 23596 25659
rect 23603 25640 23606 25654
rect 23604 25639 23606 25640
rect 23652 25639 23654 25659
rect 23676 25639 23678 25659
rect 23724 25656 23726 25659
rect 23724 25639 23727 25656
rect 23772 25639 23774 25659
rect 23820 25639 23822 25659
rect 23916 25639 23918 25659
rect 24012 25639 24014 25659
rect 24060 25639 24062 25659
rect 24156 25639 24158 25659
rect 24492 25639 24494 25659
rect 24516 25639 24518 25659
rect 24588 25639 24590 25659
rect 24612 25639 24614 25659
rect 24684 25639 24686 25659
rect 24732 25639 24734 25659
rect 24756 25639 24758 25659
rect 24780 25639 24782 25659
rect 24852 25639 24854 25659
rect 24876 25639 24878 25659
rect 24972 25639 24974 25659
rect 25068 25639 25070 25659
rect 25164 25639 25166 25659
rect 25260 25639 25262 25659
rect 25284 25639 25286 25659
rect 25356 25639 25358 25659
rect 25380 25639 25382 25659
rect 25404 25639 25406 25659
rect 25500 25639 25502 25659
rect 25596 25639 25598 25659
rect 27025 25654 27028 25659
rect 27036 25656 27038 25659
rect 27036 25654 27039 25656
rect 27025 25646 27029 25654
rect 27015 25640 27025 25646
rect 27035 25640 27039 25654
rect 27097 25646 27101 25654
rect 27087 25640 27097 25646
rect 26449 25639 26483 25640
rect -16326 25635 -14803 25639
rect -16260 25632 -16258 25635
rect -16260 25615 -16257 25632
rect -15324 25615 -15322 25635
rect -15108 25615 -15106 25635
rect -14892 25615 -14890 25635
rect -14817 25632 -14803 25635
rect -14793 25635 -14467 25639
rect -14793 25632 -14779 25635
rect -14772 25632 -14769 25635
rect -14676 25615 -14674 25635
rect -14481 25632 -14467 25635
rect -14457 25635 -5587 25639
rect -14457 25632 -14443 25635
rect -14436 25632 -14433 25635
rect -14340 25615 -14338 25635
rect -13943 25630 -13940 25635
rect -13932 25632 -13930 25635
rect -13932 25630 -13929 25632
rect -13933 25616 -13929 25630
rect -13788 25615 -13786 25635
rect -13583 25630 -13580 25635
rect -13572 25630 -13570 25635
rect -13367 25630 -13364 25635
rect -13356 25630 -13354 25635
rect -12801 25632 -12787 25635
rect -12780 25632 -12777 25635
rect -13573 25616 -13570 25630
rect -13357 25616 -13354 25630
rect -13535 25615 -13477 25616
rect -12756 25615 -12754 25635
rect -12660 25615 -12658 25635
rect -12575 25630 -12572 25635
rect -12564 25630 -12562 25635
rect -12565 25616 -12562 25630
rect -12492 25615 -12490 25635
rect -12396 25615 -12394 25635
rect -12348 25615 -12346 25635
rect -12252 25615 -12250 25635
rect -12156 25615 -12154 25635
rect -12060 25615 -12058 25635
rect -11844 25615 -11842 25635
rect -11676 25615 -11674 25635
rect -11567 25630 -11564 25635
rect -11556 25630 -11554 25635
rect -11557 25616 -11554 25630
rect -11508 25615 -11506 25635
rect -11436 25615 -11434 25635
rect -11412 25615 -11410 25635
rect -11340 25615 -11338 25635
rect -11196 25615 -11194 25635
rect -11100 25615 -11098 25635
rect -11049 25632 -11035 25635
rect -10953 25632 -10939 25635
rect -10740 25615 -10738 25635
rect -10679 25630 -10676 25635
rect -10668 25630 -10666 25635
rect -10669 25616 -10666 25630
rect -10644 25615 -10642 25635
rect -9996 25615 -9994 25635
rect -9900 25615 -9898 25635
rect -9828 25615 -9826 25635
rect -9732 25615 -9730 25635
rect -9516 25615 -9514 25635
rect -9468 25615 -9466 25635
rect -9348 25615 -9346 25635
rect -9180 25615 -9178 25635
rect -8604 25615 -8602 25635
rect -8484 25615 -8482 25635
rect -8436 25615 -8434 25635
rect -8388 25615 -8386 25635
rect -8364 25615 -8362 25635
rect -8340 25615 -8338 25635
rect -8268 25615 -8266 25635
rect -8100 25615 -8098 25635
rect -8052 25615 -8050 25635
rect -8004 25615 -8002 25635
rect -7932 25615 -7930 25635
rect -7692 25615 -7690 25635
rect -7620 25615 -7618 25635
rect -7524 25615 -7522 25635
rect -7356 25615 -7354 25635
rect -7308 25615 -7306 25635
rect -7212 25615 -7210 25635
rect -7116 25615 -7114 25635
rect -7068 25632 -7066 25635
rect -7068 25615 -7065 25632
rect -6972 25615 -6970 25635
rect -6948 25615 -6946 25635
rect -6876 25615 -6874 25635
rect -6852 25615 -6850 25635
rect -6780 25615 -6778 25635
rect -6756 25615 -6754 25635
rect -6660 25615 -6658 25635
rect -6612 25615 -6610 25635
rect -6516 25615 -6514 25635
rect -6372 25615 -6370 25635
rect -6156 25615 -6154 25635
rect -6060 25615 -6058 25635
rect -6036 25615 -6034 25635
rect -5892 25615 -5890 25635
rect -5601 25632 -5587 25635
rect -5577 25635 -4843 25639
rect -5577 25632 -5563 25635
rect -5268 25615 -5266 25635
rect -5196 25615 -5194 25635
rect -5172 25615 -5170 25635
rect -5100 25615 -5098 25635
rect -5076 25615 -5074 25635
rect -4980 25615 -4978 25635
rect -4956 25615 -4954 25635
rect -4860 25615 -4858 25635
rect -4857 25632 -4843 25635
rect -4833 25635 23693 25639
rect -4833 25632 -4819 25635
rect -4644 25615 -4642 25635
rect -4548 25615 -4546 25635
rect -4500 25615 -4498 25635
rect -4404 25615 -4402 25635
rect -4308 25615 -4306 25635
rect -4260 25615 -4258 25635
rect -4164 25615 -4162 25635
rect -4020 25615 -4018 25635
rect -3876 25615 -3874 25635
rect -3732 25615 -3730 25635
rect -3588 25615 -3586 25635
rect -3564 25615 -3562 25635
rect -3516 25615 -3514 25635
rect -3492 25615 -3490 25635
rect -3468 25615 -3466 25635
rect -3420 25615 -3418 25635
rect -3324 25615 -3322 25635
rect -3228 25615 -3226 25635
rect -3132 25615 -3130 25635
rect -3012 25615 -3010 25635
rect -2964 25615 -2962 25635
rect -2916 25615 -2914 25635
rect -2892 25615 -2890 25635
rect -2868 25615 -2866 25635
rect -2820 25615 -2818 25635
rect -2796 25615 -2794 25635
rect -2772 25615 -2770 25635
rect -2676 25615 -2674 25635
rect -2580 25615 -2578 25635
rect -2364 25615 -2362 25635
rect -2316 25615 -2314 25635
rect -2268 25615 -2266 25635
rect -2244 25615 -2242 25635
rect -2172 25615 -2170 25635
rect -2148 25615 -2146 25635
rect -2076 25615 -2074 25635
rect -2052 25615 -2050 25635
rect -1980 25615 -1978 25635
rect -1884 25615 -1882 25635
rect -1572 25615 -1570 25635
rect -1476 25615 -1474 25635
rect -1380 25615 -1378 25635
rect -1356 25615 -1354 25635
rect -1308 25615 -1306 25635
rect -1260 25615 -1258 25635
rect -1140 25615 -1138 25635
rect -708 25615 -706 25635
rect -612 25615 -610 25635
rect -588 25615 -586 25635
rect -540 25615 -538 25635
rect -492 25615 -490 25635
rect -444 25615 -442 25635
rect -396 25615 -394 25635
rect -300 25615 -298 25635
rect -276 25615 -274 25635
rect -228 25615 -226 25635
rect -12 25615 -10 25635
rect 156 25615 158 25635
rect 204 25615 206 25635
rect 252 25615 254 25635
rect 348 25615 350 25635
rect 468 25615 470 25635
rect 492 25615 494 25635
rect 564 25615 566 25635
rect 588 25615 590 25635
rect 636 25615 638 25635
rect 660 25615 662 25635
rect 732 25615 734 25635
rect 1092 25615 1094 25635
rect 1308 25615 1310 25635
rect 1332 25615 1334 25635
rect 1380 25615 1382 25635
rect 1428 25615 1430 25635
rect 1476 25615 1478 25635
rect 1644 25615 1646 25635
rect 1692 25615 1694 25635
rect 1740 25615 1742 25635
rect 1788 25615 1790 25635
rect 2028 25615 2030 25635
rect 2076 25615 2078 25635
rect 2100 25615 2102 25635
rect 2124 25615 2126 25635
rect 2172 25615 2174 25635
rect 2220 25615 2222 25635
rect 2316 25615 2318 25635
rect 2412 25615 2414 25635
rect 2460 25615 2462 25635
rect 2508 25615 2510 25635
rect 2580 25615 2582 25635
rect 2604 25615 2606 25635
rect 2676 25615 2678 25635
rect 2700 25615 2702 25635
rect 2748 25615 2750 25635
rect 2772 25615 2774 25635
rect 2796 25615 2798 25635
rect 2844 25615 2846 25635
rect 2868 25615 2870 25635
rect 2892 25615 2894 25635
rect 2940 25615 2942 25635
rect 3012 25615 3014 25635
rect 3108 25615 3110 25635
rect 3252 25615 3254 25635
rect 3348 25615 3350 25635
rect 3396 25615 3398 25635
rect 3564 25615 3566 25635
rect 3636 25615 3638 25635
rect 3660 25615 3662 25635
rect 3732 25615 3734 25635
rect 3828 25615 3830 25635
rect 3924 25615 3926 25635
rect 4020 25615 4022 25635
rect 4044 25615 4046 25635
rect 4092 25615 4094 25635
rect 4116 25615 4118 25635
rect 4140 25615 4142 25635
rect 4188 25615 4190 25635
rect 4212 25615 4214 25635
rect 4236 25615 4238 25635
rect 4308 25615 4310 25635
rect 4332 25615 4334 25635
rect 4404 25615 4406 25635
rect 4500 25615 4502 25635
rect 4596 25615 4598 25635
rect 4692 25615 4694 25635
rect 4860 25615 4862 25635
rect 4956 25615 4958 25635
rect 4980 25615 4982 25635
rect 5004 25615 5006 25635
rect 5052 25615 5054 25635
rect 5100 25615 5102 25635
rect 5124 25615 5126 25635
rect 5220 25615 5222 25635
rect 5268 25615 5270 25635
rect 5388 25615 5390 25635
rect 5484 25615 5486 25635
rect 5508 25615 5510 25635
rect 5532 25615 5534 25635
rect 5628 25615 5630 25635
rect 5652 25615 5654 25635
rect 5748 25615 5750 25635
rect 5796 25615 5798 25635
rect 5844 25615 5846 25635
rect 5892 25615 5894 25635
rect 6132 25615 6134 25635
rect 6180 25615 6182 25635
rect 6228 25615 6230 25635
rect 6252 25615 6254 25635
rect 6276 25615 6278 25635
rect 6324 25615 6326 25635
rect 6372 25615 6374 25635
rect 6492 25615 6494 25635
rect 6588 25615 6590 25635
rect 6612 25615 6614 25635
rect 6660 25615 6662 25635
rect 6684 25615 6686 25635
rect 6708 25615 6710 25635
rect 6780 25615 6782 25635
rect 6804 25615 6806 25635
rect 6900 25615 6902 25635
rect 6924 25615 6926 25635
rect 7020 25615 7022 25635
rect 7068 25615 7070 25635
rect 7164 25615 7166 25635
rect 7236 25615 7238 25635
rect 7332 25615 7334 25635
rect 7380 25615 7382 25635
rect 7428 25615 7430 25635
rect 7452 25615 7454 25635
rect 7476 25615 7478 25635
rect 7524 25615 7526 25635
rect 7548 25615 7550 25635
rect 7572 25615 7574 25635
rect 7620 25615 7622 25635
rect 7644 25615 7646 25635
rect 7668 25615 7670 25635
rect 7788 25615 7790 25635
rect 7884 25615 7886 25635
rect 7956 25615 7958 25635
rect 7980 25615 7982 25635
rect 8028 25615 8030 25635
rect 8196 25615 8198 25635
rect 8244 25615 8246 25635
rect 8268 25615 8270 25635
rect 8292 25615 8294 25635
rect 8340 25615 8342 25635
rect 8364 25615 8366 25635
rect 8388 25615 8390 25635
rect 8436 25615 8438 25635
rect 8604 25615 8606 25635
rect 8652 25615 8654 25635
rect 8700 25615 8702 25635
rect 8724 25615 8726 25635
rect 8748 25615 8750 25635
rect 8820 25615 8822 25635
rect 8844 25615 8846 25635
rect 8868 25615 8870 25635
rect 9516 25615 9518 25635
rect 9612 25615 9614 25635
rect 9660 25615 9662 25635
rect 9684 25615 9686 25635
rect 9708 25615 9710 25635
rect 9756 25615 9758 25635
rect 9780 25615 9782 25635
rect 9804 25615 9806 25635
rect 9852 25615 9854 25635
rect 9900 25615 9902 25635
rect 9948 25615 9950 25635
rect 9996 25615 9998 25635
rect 10068 25615 10070 25635
rect 10092 25615 10094 25635
rect 10116 25615 10118 25635
rect 10164 25615 10166 25635
rect 10188 25615 10190 25635
rect 10212 25615 10214 25635
rect 10284 25615 10286 25635
rect 10308 25615 10310 25635
rect 10332 25615 10334 25635
rect 10380 25615 10382 25635
rect 10404 25615 10406 25635
rect 10428 25615 10430 25635
rect 10476 25615 10478 25635
rect 10500 25615 10502 25635
rect 10524 25615 10526 25635
rect 10572 25615 10574 25635
rect 10596 25615 10598 25635
rect 10620 25615 10622 25635
rect 10668 25615 10670 25635
rect 10692 25615 10694 25635
rect 10716 25615 10718 25635
rect 10788 25615 10790 25635
rect 10836 25615 10838 25635
rect 10956 25615 10958 25635
rect 11004 25615 11006 25635
rect 11052 25615 11054 25635
rect 11100 25615 11102 25635
rect 11172 25615 11174 25635
rect 11220 25615 11222 25635
rect 11340 25615 11342 25635
rect 11436 25615 11438 25635
rect 11532 25615 11534 25635
rect 11580 25615 11582 25635
rect 11628 25615 11630 25635
rect 11676 25615 11678 25635
rect 11724 25615 11726 25635
rect 11772 25615 11774 25635
rect 11796 25615 11798 25635
rect 11892 25615 11894 25635
rect 11988 25615 11990 25635
rect 12060 25615 12062 25635
rect 12132 25615 12134 25635
rect 12228 25615 12230 25635
rect 12276 25615 12278 25635
rect 12324 25615 12326 25635
rect 12420 25615 12422 25635
rect 12444 25615 12446 25635
rect 12492 25615 12494 25635
rect 12516 25615 12518 25635
rect 12540 25615 12542 25635
rect 12588 25615 12590 25635
rect 12636 25615 12638 25635
rect 12732 25615 12734 25635
rect 12756 25615 12758 25635
rect 12804 25615 12806 25635
rect 12828 25615 12830 25635
rect 12852 25615 12854 25635
rect 12948 25615 12950 25635
rect 12972 25615 12974 25635
rect 13044 25615 13046 25635
rect 13068 25615 13070 25635
rect 13116 25615 13118 25635
rect 13284 25615 13286 25635
rect 13332 25615 13334 25635
rect 13572 25615 13574 25635
rect 13620 25615 13622 25635
rect 13668 25615 13670 25635
rect 13716 25615 13718 25635
rect 13764 25615 13766 25635
rect 13860 25615 13862 25635
rect 13956 25615 13958 25635
rect 14004 25615 14006 25635
rect 14100 25615 14102 25635
rect 14196 25616 14198 25635
rect 14161 25615 14219 25616
rect 14292 25615 14294 25635
rect 15180 25615 15182 25635
rect 15276 25615 15278 25635
rect 15420 25615 15422 25635
rect 15492 25615 15494 25635
rect 15615 25632 15629 25635
rect 15636 25632 15639 25635
rect 15660 25615 15662 25635
rect 15708 25615 15710 25635
rect 15732 25615 15734 25635
rect 15756 25615 15758 25635
rect 15804 25615 15806 25635
rect 15828 25615 15830 25635
rect 15852 25615 15854 25635
rect 15900 25615 15902 25635
rect 15948 25615 15950 25635
rect 16044 25615 16046 25635
rect 16068 25615 16070 25635
rect 16164 25615 16166 25635
rect 16260 25615 16262 25635
rect 16308 25615 16310 25635
rect 16332 25615 16334 25635
rect 16356 25615 16358 25635
rect 16404 25615 16406 25635
rect 16452 25615 16454 25635
rect 16548 25615 16550 25635
rect 16572 25615 16574 25635
rect 16620 25615 16622 25635
rect 16668 25615 16670 25635
rect 16716 25615 16718 25635
rect 16764 25615 16766 25635
rect 16812 25615 16814 25635
rect 16884 25615 16886 25635
rect 16908 25615 16910 25635
rect 16980 25615 16982 25635
rect 17052 25615 17054 25635
rect 17196 25615 17198 25635
rect 17220 25615 17222 25635
rect 17292 25615 17294 25635
rect 17316 25615 17318 25635
rect 18084 25615 18086 25635
rect 18132 25615 18134 25635
rect 18228 25615 18230 25635
rect 18396 25615 18398 25635
rect 18492 25615 18494 25635
rect 18516 25615 18518 25635
rect 18564 25615 18566 25635
rect 18612 25615 18614 25635
rect 18660 25615 18662 25635
rect 18708 25616 18710 25635
rect 18673 25615 18731 25616
rect 18756 25615 18758 25635
rect 18804 25615 18806 25635
rect 18852 25615 18854 25635
rect 18900 25615 18902 25635
rect 18996 25615 18998 25635
rect 19020 25615 19022 25635
rect 19092 25615 19094 25635
rect 19116 25615 19118 25635
rect 19140 25615 19142 25635
rect 19188 25615 19190 25635
rect 19236 25615 19238 25635
rect 19332 25615 19334 25635
rect 19476 25615 19478 25635
rect 19527 25632 19541 25635
rect 19788 25615 19790 25635
rect 19836 25615 19838 25635
rect 19860 25615 19862 25635
rect 19884 25615 19886 25635
rect 19932 25615 19934 25635
rect 19956 25615 19958 25635
rect 19980 25615 19982 25635
rect 20028 25615 20030 25635
rect 20052 25615 20054 25635
rect 20076 25615 20078 25635
rect 20148 25615 20150 25635
rect 20172 25615 20174 25635
rect 20196 25615 20198 25635
rect 20268 25615 20270 25635
rect 20292 25615 20294 25635
rect 20388 25615 20390 25635
rect 20412 25615 20414 25635
rect 20508 25615 20510 25635
rect 20556 25615 20558 25635
rect 20604 25615 20606 25635
rect 20916 25615 20918 25635
rect 20964 25615 20966 25635
rect 21012 25615 21014 25635
rect 21060 25615 21062 25635
rect 21108 25615 21110 25635
rect 21204 25615 21206 25635
rect 21300 25615 21302 25635
rect 21324 25615 21326 25635
rect 21444 25615 21446 25635
rect 21468 25615 21470 25635
rect 21564 25615 21566 25635
rect 21588 25615 21590 25635
rect 21684 25615 21686 25635
rect 21708 25615 21710 25635
rect 21828 25615 21830 25635
rect 21924 25615 21926 25635
rect 22068 25615 22070 25635
rect 22188 25615 22190 25635
rect 22212 25615 22214 25635
rect 22884 25615 22886 25635
rect 22980 25615 22982 25635
rect 23076 25615 23078 25635
rect 23100 25615 23102 25635
rect 23124 25615 23126 25635
rect 23244 25615 23246 25635
rect 23340 25615 23342 25635
rect 23412 25615 23414 25635
rect 23508 25615 23510 25635
rect 23556 25615 23558 25635
rect 23604 25615 23606 25635
rect 23652 25615 23654 25635
rect 23676 25615 23678 25635
rect 23679 25632 23693 25635
rect 23703 25635 26483 25639
rect 23703 25632 23717 25635
rect 23724 25632 23727 25635
rect 23772 25615 23774 25635
rect 23820 25615 23822 25635
rect 23916 25615 23918 25635
rect 24012 25615 24014 25635
rect 24060 25615 24062 25635
rect 24156 25615 24158 25635
rect 24492 25615 24494 25635
rect 24516 25615 24518 25635
rect 24588 25615 24590 25635
rect 24612 25615 24614 25635
rect 24684 25615 24686 25635
rect 24732 25615 24734 25635
rect 24756 25615 24758 25635
rect 24780 25615 24782 25635
rect 24852 25615 24854 25635
rect 24876 25615 24878 25635
rect 24972 25615 24974 25635
rect 25068 25615 25070 25635
rect 25164 25615 25166 25635
rect 25260 25615 25262 25635
rect 25284 25615 25286 25635
rect 25356 25615 25358 25635
rect 25380 25615 25382 25635
rect 25404 25615 25406 25635
rect 25500 25615 25502 25635
rect 25596 25615 25598 25635
rect 26401 25615 26435 25616
rect -16281 25611 -10435 25615
rect -16281 25608 -16267 25611
rect -16260 25608 -16257 25611
rect -15455 25591 -15397 25592
rect -15324 25591 -15322 25611
rect -15108 25591 -15106 25611
rect -14892 25591 -14890 25611
rect -14676 25591 -14674 25611
rect -14340 25591 -14338 25611
rect -13953 25608 -13939 25611
rect -13857 25608 -13843 25611
rect -13788 25591 -13786 25611
rect -13497 25608 -13483 25611
rect -13281 25608 -13267 25611
rect -13428 25591 -13425 25608
rect -13007 25591 -12973 25592
rect -12756 25591 -12754 25611
rect -12660 25591 -12658 25611
rect -12492 25591 -12490 25611
rect -12489 25608 -12475 25611
rect -12396 25591 -12394 25611
rect -12348 25591 -12346 25611
rect -12252 25591 -12250 25611
rect -12156 25591 -12154 25611
rect -12060 25591 -12058 25611
rect -11844 25591 -11842 25611
rect -11676 25591 -11674 25611
rect -11508 25591 -11506 25611
rect -11481 25608 -11467 25611
rect -11436 25591 -11434 25611
rect -11412 25591 -11410 25611
rect -11340 25591 -11338 25611
rect -11289 25608 -11275 25611
rect -11196 25591 -11194 25611
rect -11100 25591 -11098 25611
rect -10740 25591 -10738 25611
rect -10644 25591 -10642 25611
rect -10593 25608 -10579 25611
rect -10449 25608 -10435 25611
rect -10425 25611 -7099 25615
rect -10425 25608 -10411 25611
rect -9996 25591 -9994 25611
rect -9935 25591 -9901 25592
rect -9900 25591 -9898 25611
rect -9828 25591 -9826 25611
rect -9732 25591 -9730 25611
rect -9516 25591 -9514 25611
rect -9468 25591 -9466 25611
rect -9348 25591 -9346 25611
rect -9180 25591 -9178 25611
rect -8604 25591 -8602 25611
rect -8484 25591 -8482 25611
rect -8436 25591 -8434 25611
rect -8388 25591 -8386 25611
rect -8364 25591 -8362 25611
rect -8340 25591 -8338 25611
rect -8268 25591 -8266 25611
rect -8100 25591 -8098 25611
rect -8052 25591 -8050 25611
rect -8004 25591 -8002 25611
rect -7932 25591 -7930 25611
rect -7692 25591 -7690 25611
rect -7620 25591 -7618 25611
rect -7524 25591 -7522 25611
rect -7356 25591 -7354 25611
rect -7308 25591 -7306 25611
rect -7212 25591 -7210 25611
rect -7116 25592 -7114 25611
rect -7113 25608 -7099 25611
rect -7089 25611 26435 25615
rect -7089 25608 -7075 25611
rect -7068 25608 -7065 25611
rect -7151 25591 -7093 25592
rect -6972 25591 -6970 25611
rect -6948 25591 -6946 25611
rect -6876 25591 -6874 25611
rect -6852 25591 -6850 25611
rect -6780 25591 -6778 25611
rect -6756 25591 -6754 25611
rect -6660 25591 -6658 25611
rect -6612 25591 -6610 25611
rect -6516 25591 -6514 25611
rect -6372 25591 -6370 25611
rect -6156 25591 -6154 25611
rect -6060 25591 -6058 25611
rect -6036 25591 -6034 25611
rect -5892 25591 -5890 25611
rect -5268 25591 -5266 25611
rect -5196 25591 -5194 25611
rect -5172 25591 -5170 25611
rect -5100 25591 -5098 25611
rect -5076 25591 -5074 25611
rect -4980 25591 -4978 25611
rect -4956 25591 -4954 25611
rect -4860 25591 -4858 25611
rect -4644 25591 -4642 25611
rect -4548 25591 -4546 25611
rect -4500 25591 -4498 25611
rect -4404 25591 -4402 25611
rect -4308 25591 -4306 25611
rect -4260 25591 -4258 25611
rect -4164 25591 -4162 25611
rect -4020 25591 -4018 25611
rect -3876 25591 -3874 25611
rect -3732 25591 -3730 25611
rect -3588 25591 -3586 25611
rect -3564 25591 -3562 25611
rect -3516 25591 -3514 25611
rect -3492 25591 -3490 25611
rect -3468 25591 -3466 25611
rect -3420 25591 -3418 25611
rect -3324 25591 -3322 25611
rect -3228 25591 -3226 25611
rect -3132 25591 -3130 25611
rect -3012 25591 -3010 25611
rect -2964 25591 -2962 25611
rect -2916 25591 -2914 25611
rect -2892 25591 -2890 25611
rect -2868 25591 -2866 25611
rect -2820 25591 -2818 25611
rect -2796 25591 -2794 25611
rect -2772 25591 -2770 25611
rect -2676 25591 -2674 25611
rect -2580 25591 -2578 25611
rect -2364 25591 -2362 25611
rect -2316 25591 -2314 25611
rect -2268 25591 -2266 25611
rect -2244 25591 -2242 25611
rect -2172 25591 -2170 25611
rect -2148 25591 -2146 25611
rect -2076 25591 -2074 25611
rect -2052 25591 -2050 25611
rect -1980 25591 -1978 25611
rect -1884 25591 -1882 25611
rect -1572 25591 -1570 25611
rect -1476 25591 -1474 25611
rect -1380 25591 -1378 25611
rect -1356 25591 -1354 25611
rect -1308 25591 -1306 25611
rect -1260 25591 -1258 25611
rect -1140 25591 -1138 25611
rect -708 25591 -706 25611
rect -612 25591 -610 25611
rect -588 25591 -586 25611
rect -540 25591 -538 25611
rect -492 25591 -490 25611
rect -444 25591 -442 25611
rect -396 25591 -394 25611
rect -300 25591 -298 25611
rect -276 25591 -274 25611
rect -228 25591 -226 25611
rect -12 25591 -10 25611
rect 156 25591 158 25611
rect 204 25591 206 25611
rect 252 25591 254 25611
rect 348 25591 350 25611
rect 468 25591 470 25611
rect 492 25591 494 25611
rect 564 25591 566 25611
rect 588 25591 590 25611
rect 636 25591 638 25611
rect 660 25591 662 25611
rect 732 25591 734 25611
rect 1092 25591 1094 25611
rect 1308 25591 1310 25611
rect 1332 25591 1334 25611
rect 1380 25591 1382 25611
rect 1428 25591 1430 25611
rect 1476 25591 1478 25611
rect 1644 25591 1646 25611
rect 1692 25591 1694 25611
rect 1740 25591 1742 25611
rect 1788 25591 1790 25611
rect 2028 25591 2030 25611
rect 2076 25591 2078 25611
rect 2100 25591 2102 25611
rect 2124 25591 2126 25611
rect 2172 25591 2174 25611
rect 2220 25591 2222 25611
rect 2316 25591 2318 25611
rect 2412 25591 2414 25611
rect 2460 25591 2462 25611
rect 2508 25591 2510 25611
rect 2580 25591 2582 25611
rect 2604 25591 2606 25611
rect 2676 25591 2678 25611
rect 2700 25591 2702 25611
rect 2748 25591 2750 25611
rect 2772 25591 2774 25611
rect 2796 25591 2798 25611
rect 2844 25591 2846 25611
rect 2868 25591 2870 25611
rect 2892 25591 2894 25611
rect 2940 25591 2942 25611
rect 3012 25591 3014 25611
rect 3108 25591 3110 25611
rect 3252 25591 3254 25611
rect 3348 25591 3350 25611
rect 3396 25591 3398 25611
rect 3564 25591 3566 25611
rect 3636 25591 3638 25611
rect 3660 25591 3662 25611
rect 3732 25591 3734 25611
rect 3828 25591 3830 25611
rect 3924 25591 3926 25611
rect 4020 25591 4022 25611
rect 4044 25591 4046 25611
rect 4092 25591 4094 25611
rect 4116 25591 4118 25611
rect 4140 25591 4142 25611
rect 4188 25591 4190 25611
rect 4212 25591 4214 25611
rect 4236 25591 4238 25611
rect 4308 25591 4310 25611
rect 4332 25591 4334 25611
rect 4404 25591 4406 25611
rect 4500 25591 4502 25611
rect 4596 25591 4598 25611
rect 4692 25591 4694 25611
rect 4860 25591 4862 25611
rect 4956 25591 4958 25611
rect 4980 25591 4982 25611
rect 5004 25591 5006 25611
rect 5052 25591 5054 25611
rect 5100 25591 5102 25611
rect 5124 25591 5126 25611
rect 5220 25591 5222 25611
rect 5268 25591 5270 25611
rect 5388 25591 5390 25611
rect 5484 25591 5486 25611
rect 5508 25591 5510 25611
rect 5532 25591 5534 25611
rect 5628 25591 5630 25611
rect 5652 25591 5654 25611
rect 5748 25591 5750 25611
rect 5796 25591 5798 25611
rect 5844 25591 5846 25611
rect 5892 25591 5894 25611
rect 6132 25591 6134 25611
rect 6180 25591 6182 25611
rect 6228 25591 6230 25611
rect 6252 25591 6254 25611
rect 6276 25591 6278 25611
rect 6324 25591 6326 25611
rect 6372 25591 6374 25611
rect 6492 25591 6494 25611
rect 6588 25591 6590 25611
rect 6612 25591 6614 25611
rect 6660 25591 6662 25611
rect 6684 25591 6686 25611
rect 6708 25591 6710 25611
rect 6780 25591 6782 25611
rect 6804 25591 6806 25611
rect 6900 25591 6902 25611
rect 6924 25591 6926 25611
rect 7020 25591 7022 25611
rect 7068 25591 7070 25611
rect 7164 25591 7166 25611
rect 7236 25591 7238 25611
rect 7332 25591 7334 25611
rect 7380 25591 7382 25611
rect 7428 25591 7430 25611
rect 7452 25591 7454 25611
rect 7476 25591 7478 25611
rect 7524 25591 7526 25611
rect 7548 25591 7550 25611
rect 7572 25591 7574 25611
rect 7620 25591 7622 25611
rect 7644 25591 7646 25611
rect 7668 25591 7670 25611
rect 7788 25591 7790 25611
rect 7884 25591 7886 25611
rect 7956 25591 7958 25611
rect 7980 25591 7982 25611
rect 8028 25591 8030 25611
rect 8196 25591 8198 25611
rect 8244 25591 8246 25611
rect 8268 25591 8270 25611
rect 8292 25591 8294 25611
rect 8340 25591 8342 25611
rect 8364 25591 8366 25611
rect 8388 25591 8390 25611
rect 8436 25591 8438 25611
rect 8604 25591 8606 25611
rect 8652 25591 8654 25611
rect 8700 25591 8702 25611
rect 8724 25591 8726 25611
rect 8748 25591 8750 25611
rect 8820 25591 8822 25611
rect 8844 25591 8846 25611
rect 8868 25591 8870 25611
rect 9516 25591 9518 25611
rect 9612 25591 9614 25611
rect 9660 25591 9662 25611
rect 9684 25591 9686 25611
rect 9708 25591 9710 25611
rect 9756 25591 9758 25611
rect 9780 25591 9782 25611
rect 9804 25591 9806 25611
rect 9852 25591 9854 25611
rect 9900 25591 9902 25611
rect 9948 25591 9950 25611
rect 9996 25591 9998 25611
rect 10068 25591 10070 25611
rect 10092 25591 10094 25611
rect 10116 25591 10118 25611
rect 10164 25591 10166 25611
rect 10188 25591 10190 25611
rect 10212 25591 10214 25611
rect 10284 25591 10286 25611
rect 10308 25591 10310 25611
rect 10332 25591 10334 25611
rect 10380 25591 10382 25611
rect 10404 25591 10406 25611
rect 10428 25591 10430 25611
rect 10476 25591 10478 25611
rect 10500 25591 10502 25611
rect 10524 25591 10526 25611
rect 10572 25591 10574 25611
rect 10596 25591 10598 25611
rect 10620 25591 10622 25611
rect 10668 25591 10670 25611
rect 10692 25591 10694 25611
rect 10716 25591 10718 25611
rect 10788 25591 10790 25611
rect 10836 25591 10838 25611
rect 10956 25591 10958 25611
rect 11004 25591 11006 25611
rect 11052 25591 11054 25611
rect 11100 25591 11102 25611
rect 11172 25591 11174 25611
rect 11220 25591 11222 25611
rect 11340 25591 11342 25611
rect 11436 25591 11438 25611
rect 11532 25591 11534 25611
rect 11580 25591 11582 25611
rect 11628 25591 11630 25611
rect 11676 25591 11678 25611
rect 11724 25591 11726 25611
rect 11772 25591 11774 25611
rect 11796 25591 11798 25611
rect 11892 25591 11894 25611
rect 11988 25591 11990 25611
rect 12060 25591 12062 25611
rect 12132 25591 12134 25611
rect 12228 25591 12230 25611
rect 12276 25591 12278 25611
rect 12324 25591 12326 25611
rect 12420 25591 12422 25611
rect 12444 25591 12446 25611
rect 12492 25591 12494 25611
rect 12516 25591 12518 25611
rect 12540 25591 12542 25611
rect 12588 25591 12590 25611
rect 12636 25591 12638 25611
rect 12732 25591 12734 25611
rect 12756 25591 12758 25611
rect 12804 25591 12806 25611
rect 12828 25591 12830 25611
rect 12852 25591 12854 25611
rect 12948 25591 12950 25611
rect 12972 25591 12974 25611
rect 13044 25591 13046 25611
rect 13068 25591 13070 25611
rect 13116 25591 13118 25611
rect 13284 25591 13286 25611
rect 13332 25591 13334 25611
rect 13572 25591 13574 25611
rect 13620 25591 13622 25611
rect 13668 25591 13670 25611
rect 13716 25591 13718 25611
rect 13764 25591 13766 25611
rect 13860 25591 13862 25611
rect 13956 25591 13958 25611
rect 14004 25591 14006 25611
rect 14100 25591 14102 25611
rect 14185 25606 14188 25611
rect 14196 25606 14198 25611
rect 14195 25592 14198 25606
rect 14292 25608 14294 25611
rect 14292 25591 14295 25608
rect 15180 25591 15182 25611
rect 15276 25591 15278 25611
rect 15420 25591 15422 25611
rect 15492 25591 15494 25611
rect 15660 25591 15662 25611
rect 15708 25591 15710 25611
rect 15732 25591 15734 25611
rect 15756 25591 15758 25611
rect 15804 25591 15806 25611
rect 15828 25591 15830 25611
rect 15852 25591 15854 25611
rect 15900 25591 15902 25611
rect 15948 25591 15950 25611
rect 16044 25591 16046 25611
rect 16068 25591 16070 25611
rect 16164 25591 16166 25611
rect 16260 25591 16262 25611
rect 16308 25591 16310 25611
rect 16332 25591 16334 25611
rect 16356 25591 16358 25611
rect 16404 25591 16406 25611
rect 16452 25591 16454 25611
rect 16548 25591 16550 25611
rect 16572 25591 16574 25611
rect 16620 25591 16622 25611
rect 16668 25591 16670 25611
rect 16716 25591 16718 25611
rect 16764 25591 16766 25611
rect 16812 25591 16814 25611
rect 16884 25591 16886 25611
rect 16908 25591 16910 25611
rect 16980 25591 16982 25611
rect 17052 25591 17054 25611
rect 17196 25591 17198 25611
rect 17220 25591 17222 25611
rect 17292 25591 17294 25611
rect 17316 25591 17318 25611
rect 18084 25591 18086 25611
rect 18132 25591 18134 25611
rect 18228 25591 18230 25611
rect 18396 25591 18398 25611
rect 18492 25591 18494 25611
rect 18516 25591 18518 25611
rect 18564 25591 18566 25611
rect 18612 25591 18614 25611
rect 18660 25591 18662 25611
rect 18697 25606 18700 25611
rect 18708 25606 18710 25611
rect 18707 25592 18710 25606
rect 18756 25591 18758 25611
rect 18804 25608 18806 25611
rect 18804 25591 18807 25608
rect 18852 25591 18854 25611
rect 18900 25591 18902 25611
rect 18996 25591 18998 25611
rect 19020 25591 19022 25611
rect 19092 25591 19094 25611
rect 19116 25591 19118 25611
rect 19140 25591 19142 25611
rect 19188 25591 19190 25611
rect 19236 25591 19238 25611
rect 19332 25591 19334 25611
rect 19476 25591 19478 25611
rect 19788 25591 19790 25611
rect 19836 25591 19838 25611
rect 19860 25591 19862 25611
rect 19884 25591 19886 25611
rect 19932 25591 19934 25611
rect 19956 25591 19958 25611
rect 19980 25591 19982 25611
rect 20028 25591 20030 25611
rect 20052 25591 20054 25611
rect 20076 25591 20078 25611
rect 20148 25591 20150 25611
rect 20172 25591 20174 25611
rect 20196 25591 20198 25611
rect 20268 25591 20270 25611
rect 20292 25591 20294 25611
rect 20388 25591 20390 25611
rect 20412 25591 20414 25611
rect 20508 25591 20510 25611
rect 20556 25591 20558 25611
rect 20604 25591 20606 25611
rect 20916 25591 20918 25611
rect 20964 25591 20966 25611
rect 21012 25591 21014 25611
rect 21060 25591 21062 25611
rect 21108 25591 21110 25611
rect 21204 25591 21206 25611
rect 21300 25591 21302 25611
rect 21324 25591 21326 25611
rect 21444 25591 21446 25611
rect 21468 25591 21470 25611
rect 21564 25591 21566 25611
rect 21588 25591 21590 25611
rect 21684 25591 21686 25611
rect 21708 25591 21710 25611
rect 21828 25591 21830 25611
rect 21924 25591 21926 25611
rect 22068 25591 22070 25611
rect 22188 25591 22190 25611
rect 22212 25591 22214 25611
rect 22884 25591 22886 25611
rect 22980 25591 22982 25611
rect 23076 25591 23078 25611
rect 23100 25591 23102 25611
rect 23124 25591 23126 25611
rect 23244 25591 23246 25611
rect 23340 25591 23342 25611
rect 23353 25591 23411 25592
rect 23412 25591 23414 25611
rect 23508 25591 23510 25611
rect 23556 25591 23558 25611
rect 23604 25591 23606 25611
rect 23652 25591 23654 25611
rect 23676 25591 23678 25611
rect 23772 25591 23774 25611
rect 23820 25591 23822 25611
rect 23916 25591 23918 25611
rect 24012 25591 24014 25611
rect 24060 25591 24062 25611
rect 24156 25591 24158 25611
rect 24492 25591 24494 25611
rect 24516 25591 24518 25611
rect 24588 25591 24590 25611
rect 24612 25591 24614 25611
rect 24684 25591 24686 25611
rect 24732 25591 24734 25611
rect 24756 25591 24758 25611
rect 24780 25591 24782 25611
rect 24852 25591 24854 25611
rect 24876 25591 24878 25611
rect 24972 25591 24974 25611
rect 25068 25591 25070 25611
rect 25164 25591 25166 25611
rect 25260 25591 25262 25611
rect 25284 25591 25286 25611
rect 25356 25591 25358 25611
rect 25380 25591 25382 25611
rect 25404 25591 25406 25611
rect 25500 25591 25502 25611
rect 25596 25591 25598 25611
rect 26185 25591 26219 25592
rect -16233 25587 -13435 25591
rect -16233 25584 -16219 25587
rect -15324 25584 -15322 25587
rect -15324 25567 -15321 25584
rect -15108 25567 -15106 25587
rect -14892 25567 -14890 25587
rect -14831 25567 -14797 25568
rect -14676 25567 -14674 25587
rect -14340 25567 -14338 25587
rect -13788 25567 -13786 25587
rect -13449 25584 -13435 25587
rect -13428 25587 14261 25591
rect -13428 25584 -13411 25587
rect -13428 25567 -13426 25584
rect -12756 25567 -12754 25587
rect -12660 25567 -12658 25587
rect -12492 25567 -12490 25587
rect -12396 25567 -12394 25587
rect -12348 25567 -12346 25587
rect -12252 25567 -12250 25587
rect -12156 25567 -12154 25587
rect -12060 25567 -12058 25587
rect -11844 25567 -11842 25587
rect -11676 25567 -11674 25587
rect -11508 25567 -11506 25587
rect -11436 25567 -11434 25587
rect -11412 25567 -11410 25587
rect -11340 25567 -11338 25587
rect -11196 25567 -11194 25587
rect -11100 25567 -11098 25587
rect -10740 25567 -10738 25587
rect -10644 25567 -10642 25587
rect -9996 25567 -9994 25587
rect -9900 25567 -9898 25587
rect -9828 25584 -9826 25587
rect -9828 25567 -9825 25584
rect -9732 25567 -9730 25587
rect -9516 25567 -9514 25587
rect -9468 25567 -9466 25587
rect -9348 25567 -9346 25587
rect -9180 25567 -9178 25587
rect -8604 25567 -8602 25587
rect -8484 25568 -8482 25587
rect -8495 25567 -8461 25568
rect -8436 25567 -8434 25587
rect -8388 25567 -8386 25587
rect -8364 25567 -8362 25587
rect -8340 25567 -8338 25587
rect -8268 25567 -8266 25587
rect -8100 25567 -8098 25587
rect -8052 25567 -8050 25587
rect -8004 25567 -8002 25587
rect -7932 25567 -7930 25587
rect -7692 25567 -7690 25587
rect -7620 25567 -7618 25587
rect -7524 25567 -7522 25587
rect -7356 25567 -7354 25587
rect -7308 25567 -7306 25587
rect -7212 25567 -7210 25587
rect -7127 25582 -7124 25587
rect -7116 25582 -7114 25587
rect -7117 25568 -7114 25582
rect -7044 25567 -7041 25584
rect -6972 25567 -6970 25587
rect -6948 25567 -6946 25587
rect -6876 25567 -6874 25587
rect -6852 25567 -6850 25587
rect -6780 25567 -6778 25587
rect -6756 25567 -6754 25587
rect -6660 25567 -6658 25587
rect -6612 25567 -6610 25587
rect -6516 25567 -6514 25587
rect -6372 25567 -6370 25587
rect -6156 25567 -6154 25587
rect -6060 25567 -6058 25587
rect -6036 25567 -6034 25587
rect -5892 25567 -5890 25587
rect -5268 25567 -5266 25587
rect -5196 25567 -5194 25587
rect -5172 25567 -5170 25587
rect -5100 25567 -5098 25587
rect -5076 25567 -5074 25587
rect -4980 25567 -4978 25587
rect -4956 25567 -4954 25587
rect -4860 25567 -4858 25587
rect -4644 25567 -4642 25587
rect -4548 25568 -4546 25587
rect -4559 25567 -4525 25568
rect -4500 25567 -4498 25587
rect -4404 25567 -4402 25587
rect -4308 25567 -4306 25587
rect -4260 25567 -4258 25587
rect -4164 25567 -4162 25587
rect -4020 25567 -4018 25587
rect -3876 25567 -3874 25587
rect -3732 25567 -3730 25587
rect -3588 25567 -3586 25587
rect -3564 25567 -3562 25587
rect -3516 25567 -3514 25587
rect -3492 25567 -3490 25587
rect -3468 25567 -3466 25587
rect -3420 25567 -3418 25587
rect -3324 25567 -3322 25587
rect -3228 25567 -3226 25587
rect -3132 25567 -3130 25587
rect -3012 25567 -3010 25587
rect -2964 25567 -2962 25587
rect -2916 25567 -2914 25587
rect -2892 25567 -2890 25587
rect -2868 25567 -2866 25587
rect -2820 25567 -2818 25587
rect -2796 25567 -2794 25587
rect -2772 25567 -2770 25587
rect -2676 25567 -2674 25587
rect -2580 25567 -2578 25587
rect -2364 25567 -2362 25587
rect -2316 25567 -2314 25587
rect -2268 25567 -2266 25587
rect -2244 25567 -2242 25587
rect -2172 25567 -2170 25587
rect -2148 25567 -2146 25587
rect -2076 25567 -2074 25587
rect -2052 25567 -2050 25587
rect -1980 25567 -1978 25587
rect -1884 25567 -1882 25587
rect -1572 25567 -1570 25587
rect -1476 25567 -1474 25587
rect -1380 25567 -1378 25587
rect -1356 25567 -1354 25587
rect -1308 25567 -1306 25587
rect -1260 25567 -1258 25587
rect -1140 25567 -1138 25587
rect -708 25567 -706 25587
rect -612 25567 -610 25587
rect -588 25567 -586 25587
rect -540 25567 -538 25587
rect -492 25567 -490 25587
rect -444 25567 -442 25587
rect -396 25567 -394 25587
rect -300 25567 -298 25587
rect -276 25567 -274 25587
rect -228 25567 -226 25587
rect -12 25567 -10 25587
rect 156 25567 158 25587
rect 204 25567 206 25587
rect 252 25567 254 25587
rect 348 25567 350 25587
rect 468 25567 470 25587
rect 492 25567 494 25587
rect 564 25567 566 25587
rect 588 25567 590 25587
rect 636 25567 638 25587
rect 660 25567 662 25587
rect 732 25567 734 25587
rect 1092 25567 1094 25587
rect 1308 25567 1310 25587
rect 1332 25567 1334 25587
rect 1380 25567 1382 25587
rect 1428 25567 1430 25587
rect 1476 25567 1478 25587
rect 1644 25567 1646 25587
rect 1692 25567 1694 25587
rect 1740 25567 1742 25587
rect 1788 25567 1790 25587
rect 2028 25567 2030 25587
rect 2076 25567 2078 25587
rect 2100 25567 2102 25587
rect 2124 25567 2126 25587
rect 2172 25567 2174 25587
rect 2220 25567 2222 25587
rect 2316 25567 2318 25587
rect 2412 25567 2414 25587
rect 2460 25567 2462 25587
rect 2508 25567 2510 25587
rect 2580 25567 2582 25587
rect 2604 25567 2606 25587
rect 2676 25567 2678 25587
rect 2700 25567 2702 25587
rect 2748 25567 2750 25587
rect 2772 25567 2774 25587
rect 2796 25567 2798 25587
rect 2844 25567 2846 25587
rect 2868 25567 2870 25587
rect 2892 25567 2894 25587
rect 2940 25567 2942 25587
rect 3012 25567 3014 25587
rect 3108 25567 3110 25587
rect 3252 25567 3254 25587
rect 3348 25567 3350 25587
rect 3396 25567 3398 25587
rect 3564 25567 3566 25587
rect 3636 25567 3638 25587
rect 3660 25567 3662 25587
rect 3732 25567 3734 25587
rect 3828 25567 3830 25587
rect 3924 25567 3926 25587
rect 4020 25567 4022 25587
rect 4044 25567 4046 25587
rect 4092 25567 4094 25587
rect 4116 25567 4118 25587
rect 4140 25567 4142 25587
rect 4188 25567 4190 25587
rect 4212 25567 4214 25587
rect 4236 25567 4238 25587
rect 4308 25567 4310 25587
rect 4332 25567 4334 25587
rect 4404 25567 4406 25587
rect 4500 25567 4502 25587
rect 4596 25567 4598 25587
rect 4692 25567 4694 25587
rect 4860 25567 4862 25587
rect 4956 25567 4958 25587
rect 4980 25567 4982 25587
rect 5004 25567 5006 25587
rect 5052 25567 5054 25587
rect 5100 25567 5102 25587
rect 5124 25567 5126 25587
rect 5220 25567 5222 25587
rect 5268 25567 5270 25587
rect 5388 25567 5390 25587
rect 5484 25567 5486 25587
rect 5508 25567 5510 25587
rect 5532 25567 5534 25587
rect 5628 25567 5630 25587
rect 5652 25567 5654 25587
rect 5748 25567 5750 25587
rect 5796 25567 5798 25587
rect 5844 25567 5846 25587
rect 5892 25567 5894 25587
rect 6132 25567 6134 25587
rect 6180 25567 6182 25587
rect 6228 25567 6230 25587
rect 6252 25567 6254 25587
rect 6276 25567 6278 25587
rect 6324 25567 6326 25587
rect 6372 25567 6374 25587
rect 6492 25567 6494 25587
rect 6588 25567 6590 25587
rect 6612 25567 6614 25587
rect 6660 25567 6662 25587
rect 6684 25567 6686 25587
rect 6708 25567 6710 25587
rect 6780 25567 6782 25587
rect 6804 25567 6806 25587
rect 6900 25567 6902 25587
rect 6924 25567 6926 25587
rect 7020 25567 7022 25587
rect 7068 25567 7070 25587
rect 7164 25567 7166 25587
rect 7236 25567 7238 25587
rect 7332 25567 7334 25587
rect 7380 25567 7382 25587
rect 7428 25567 7430 25587
rect 7452 25567 7454 25587
rect 7476 25567 7478 25587
rect 7524 25567 7526 25587
rect 7548 25567 7550 25587
rect 7572 25567 7574 25587
rect 7620 25567 7622 25587
rect 7644 25567 7646 25587
rect 7668 25567 7670 25587
rect 7788 25567 7790 25587
rect 7884 25567 7886 25587
rect 7956 25567 7958 25587
rect 7980 25567 7982 25587
rect 8028 25567 8030 25587
rect 8196 25567 8198 25587
rect 8244 25567 8246 25587
rect 8268 25567 8270 25587
rect 8292 25567 8294 25587
rect 8340 25567 8342 25587
rect 8364 25567 8366 25587
rect 8388 25567 8390 25587
rect 8436 25567 8438 25587
rect 8497 25567 8531 25568
rect 8604 25567 8606 25587
rect 8617 25567 8651 25568
rect 8652 25567 8654 25587
rect 8700 25567 8702 25587
rect 8724 25567 8726 25587
rect 8748 25567 8750 25587
rect 8820 25567 8822 25587
rect 8844 25567 8846 25587
rect 8868 25567 8870 25587
rect 9516 25567 9518 25587
rect 9612 25567 9614 25587
rect 9660 25567 9662 25587
rect 9684 25567 9686 25587
rect 9708 25567 9710 25587
rect 9756 25567 9758 25587
rect 9780 25567 9782 25587
rect 9804 25567 9806 25587
rect 9852 25567 9854 25587
rect 9900 25567 9902 25587
rect 9948 25567 9950 25587
rect 9996 25567 9998 25587
rect 10068 25567 10070 25587
rect 10092 25567 10094 25587
rect 10116 25567 10118 25587
rect 10164 25567 10166 25587
rect 10188 25567 10190 25587
rect 10212 25567 10214 25587
rect 10284 25567 10286 25587
rect 10308 25567 10310 25587
rect 10332 25567 10334 25587
rect 10380 25567 10382 25587
rect 10404 25567 10406 25587
rect 10428 25567 10430 25587
rect 10476 25567 10478 25587
rect 10500 25567 10502 25587
rect 10524 25567 10526 25587
rect 10572 25567 10574 25587
rect 10596 25567 10598 25587
rect 10620 25567 10622 25587
rect 10668 25567 10670 25587
rect 10692 25567 10694 25587
rect 10716 25567 10718 25587
rect 10729 25567 10763 25568
rect 10788 25567 10790 25587
rect 10836 25567 10838 25587
rect 10956 25567 10958 25587
rect 11004 25567 11006 25587
rect 11052 25567 11054 25587
rect 11100 25567 11102 25587
rect 11172 25567 11174 25587
rect 11220 25567 11222 25587
rect 11340 25567 11342 25587
rect 11436 25567 11438 25587
rect 11532 25567 11534 25587
rect 11580 25567 11582 25587
rect 11628 25567 11630 25587
rect 11676 25567 11678 25587
rect 11724 25567 11726 25587
rect 11772 25567 11774 25587
rect 11796 25567 11798 25587
rect 11892 25567 11894 25587
rect 11988 25567 11990 25587
rect 12060 25567 12062 25587
rect 12132 25567 12134 25587
rect 12228 25567 12230 25587
rect 12276 25567 12278 25587
rect 12324 25567 12326 25587
rect 12420 25567 12422 25587
rect 12444 25567 12446 25587
rect 12492 25567 12494 25587
rect 12516 25567 12518 25587
rect 12540 25567 12542 25587
rect 12588 25567 12590 25587
rect 12636 25567 12638 25587
rect 12732 25567 12734 25587
rect 12756 25567 12758 25587
rect 12804 25567 12806 25587
rect 12828 25567 12830 25587
rect 12852 25567 12854 25587
rect 12948 25567 12950 25587
rect 12972 25567 12974 25587
rect 13044 25567 13046 25587
rect 13068 25567 13070 25587
rect 13116 25567 13118 25587
rect 13284 25567 13286 25587
rect 13332 25567 13334 25587
rect 13572 25567 13574 25587
rect 13620 25567 13622 25587
rect 13668 25567 13670 25587
rect 13716 25567 13718 25587
rect 13764 25567 13766 25587
rect 13860 25567 13862 25587
rect 13956 25567 13958 25587
rect 14004 25567 14006 25587
rect 14100 25567 14102 25587
rect 14247 25584 14261 25587
rect 14271 25587 18773 25591
rect 14271 25584 14285 25587
rect 14292 25584 14295 25587
rect 15180 25567 15182 25587
rect 15276 25567 15278 25587
rect 15420 25567 15422 25587
rect 15492 25567 15494 25587
rect 15660 25567 15662 25587
rect 15708 25567 15710 25587
rect 15732 25567 15734 25587
rect 15756 25567 15758 25587
rect 15804 25567 15806 25587
rect 15828 25567 15830 25587
rect 15852 25567 15854 25587
rect 15900 25567 15902 25587
rect 15948 25567 15950 25587
rect 16044 25567 16046 25587
rect 16068 25567 16070 25587
rect 16164 25567 16166 25587
rect 16260 25567 16262 25587
rect 16308 25567 16310 25587
rect 16332 25567 16334 25587
rect 16356 25567 16358 25587
rect 16404 25567 16406 25587
rect 16452 25567 16454 25587
rect 16548 25567 16550 25587
rect 16572 25567 16574 25587
rect 16620 25567 16622 25587
rect 16668 25567 16670 25587
rect 16716 25567 16718 25587
rect 16764 25567 16766 25587
rect 16812 25567 16814 25587
rect 16884 25567 16886 25587
rect 16908 25567 16910 25587
rect 16980 25567 16982 25587
rect 17052 25567 17054 25587
rect 17196 25567 17198 25587
rect 17220 25567 17222 25587
rect 17292 25567 17294 25587
rect 17316 25567 17318 25587
rect 18084 25567 18086 25587
rect 18132 25567 18134 25587
rect 18228 25567 18230 25587
rect 18396 25567 18398 25587
rect 18492 25567 18494 25587
rect 18516 25567 18518 25587
rect 18564 25567 18566 25587
rect 18612 25567 18614 25587
rect 18660 25567 18662 25587
rect 18756 25567 18758 25587
rect 18759 25584 18773 25587
rect 18783 25587 26219 25591
rect 18783 25584 18797 25587
rect 18804 25584 18807 25587
rect 18852 25567 18854 25587
rect 18900 25567 18902 25587
rect 18996 25567 18998 25587
rect 19020 25567 19022 25587
rect 19092 25567 19094 25587
rect 19116 25567 19118 25587
rect 19140 25567 19142 25587
rect 19188 25567 19190 25587
rect 19236 25567 19238 25587
rect 19332 25567 19334 25587
rect 19476 25567 19478 25587
rect 19788 25567 19790 25587
rect 19836 25567 19838 25587
rect 19860 25567 19862 25587
rect 19884 25567 19886 25587
rect 19932 25567 19934 25587
rect 19956 25567 19958 25587
rect 19980 25567 19982 25587
rect 20028 25567 20030 25587
rect 20052 25567 20054 25587
rect 20076 25567 20078 25587
rect 20148 25567 20150 25587
rect 20172 25567 20174 25587
rect 20196 25567 20198 25587
rect 20268 25567 20270 25587
rect 20292 25567 20294 25587
rect 20388 25567 20390 25587
rect 20412 25567 20414 25587
rect 20508 25567 20510 25587
rect 20556 25567 20558 25587
rect 20604 25567 20606 25587
rect 20916 25567 20918 25587
rect 20964 25567 20966 25587
rect 21012 25567 21014 25587
rect 21060 25567 21062 25587
rect 21108 25567 21110 25587
rect 21204 25567 21206 25587
rect 21300 25567 21302 25587
rect 21324 25567 21326 25587
rect 21444 25567 21446 25587
rect 21468 25567 21470 25587
rect 21564 25567 21566 25587
rect 21588 25567 21590 25587
rect 21684 25567 21686 25587
rect 21708 25567 21710 25587
rect 21828 25567 21830 25587
rect 21924 25567 21926 25587
rect 22068 25567 22070 25587
rect 22188 25567 22190 25587
rect 22212 25567 22214 25587
rect 22884 25567 22886 25587
rect 22980 25567 22982 25587
rect 23076 25567 23078 25587
rect 23100 25567 23102 25587
rect 23124 25567 23126 25587
rect 23244 25567 23246 25587
rect 23340 25567 23342 25587
rect 23412 25567 23414 25587
rect 23460 25567 23463 25584
rect 23508 25567 23510 25587
rect 23556 25567 23558 25587
rect 23604 25567 23606 25587
rect 23652 25567 23654 25587
rect 23676 25567 23678 25587
rect 23772 25567 23774 25587
rect 23820 25567 23822 25587
rect 23916 25567 23918 25587
rect 24012 25567 24014 25587
rect 24060 25567 24062 25587
rect 24156 25567 24158 25587
rect 24492 25567 24494 25587
rect 24516 25567 24518 25587
rect 24588 25567 24590 25587
rect 24612 25567 24614 25587
rect 24684 25567 24686 25587
rect 24732 25567 24734 25587
rect 24756 25567 24758 25587
rect 24780 25567 24782 25587
rect 24852 25567 24854 25587
rect 24876 25567 24878 25587
rect 24972 25567 24974 25587
rect 25068 25567 25070 25587
rect 25164 25567 25166 25587
rect 25260 25567 25262 25587
rect 25284 25567 25286 25587
rect 25356 25567 25358 25587
rect 25380 25567 25382 25587
rect 25404 25567 25406 25587
rect 25500 25567 25502 25587
rect 25596 25567 25598 25587
rect 25825 25567 25859 25568
rect -16209 25563 -15355 25567
rect -16209 25560 -16195 25563
rect -15369 25560 -15355 25563
rect -15345 25563 -7051 25567
rect -15345 25560 -15331 25563
rect -15324 25560 -15321 25563
rect -16079 25543 -16045 25544
rect -15647 25543 -15613 25544
rect -16079 25539 -15613 25543
rect -15455 25543 -15421 25544
rect -15108 25543 -15106 25563
rect -14892 25543 -14890 25563
rect -14676 25543 -14674 25563
rect -14340 25543 -14338 25563
rect -13788 25543 -13786 25563
rect -13428 25543 -13426 25563
rect -12921 25560 -12907 25563
rect -12756 25543 -12754 25563
rect -12660 25543 -12658 25563
rect -12599 25543 -12565 25544
rect -12492 25543 -12490 25563
rect -12396 25543 -12394 25563
rect -12348 25543 -12346 25563
rect -12252 25543 -12250 25563
rect -12156 25543 -12154 25563
rect -12060 25543 -12058 25563
rect -11844 25543 -11842 25563
rect -11676 25543 -11674 25563
rect -11508 25543 -11506 25563
rect -11436 25543 -11434 25563
rect -11412 25543 -11410 25563
rect -11340 25543 -11338 25563
rect -11196 25543 -11194 25563
rect -11100 25543 -11098 25563
rect -10740 25543 -10738 25563
rect -10644 25543 -10642 25563
rect -9996 25543 -9994 25563
rect -9900 25543 -9898 25563
rect -9849 25560 -9835 25563
rect -9828 25560 -9825 25563
rect -9732 25543 -9730 25563
rect -9516 25543 -9514 25563
rect -9468 25543 -9466 25563
rect -9348 25543 -9346 25563
rect -9180 25543 -9178 25563
rect -8604 25543 -8602 25563
rect -8495 25558 -8492 25563
rect -8484 25558 -8482 25563
rect -8485 25544 -8482 25558
rect -8436 25543 -8434 25563
rect -8388 25560 -8386 25563
rect -8388 25543 -8385 25560
rect -8364 25543 -8362 25563
rect -8340 25543 -8338 25563
rect -8268 25543 -8266 25563
rect -8100 25543 -8098 25563
rect -8052 25543 -8050 25563
rect -8004 25543 -8002 25563
rect -7932 25543 -7930 25563
rect -7692 25543 -7690 25563
rect -7620 25543 -7618 25563
rect -7524 25543 -7522 25563
rect -7356 25543 -7354 25563
rect -7308 25543 -7306 25563
rect -7212 25543 -7210 25563
rect -7065 25560 -7051 25563
rect -7044 25563 23453 25567
rect -7044 25560 -7027 25563
rect -7044 25543 -7042 25560
rect -6972 25544 -6970 25563
rect -6983 25543 -6949 25544
rect -6948 25543 -6946 25563
rect -6876 25543 -6874 25563
rect -6852 25543 -6850 25563
rect -6780 25543 -6778 25563
rect -6756 25543 -6754 25563
rect -6660 25543 -6658 25563
rect -6612 25543 -6610 25563
rect -6516 25543 -6514 25563
rect -6372 25543 -6370 25563
rect -6156 25543 -6154 25563
rect -6060 25543 -6058 25563
rect -6036 25543 -6034 25563
rect -5892 25543 -5890 25563
rect -5268 25543 -5266 25563
rect -5196 25543 -5194 25563
rect -5172 25543 -5170 25563
rect -5100 25543 -5098 25563
rect -5076 25543 -5074 25563
rect -4980 25543 -4978 25563
rect -4956 25543 -4954 25563
rect -4860 25543 -4858 25563
rect -4644 25543 -4642 25563
rect -4559 25558 -4556 25563
rect -4548 25558 -4546 25563
rect -4549 25544 -4546 25558
rect -4500 25543 -4498 25563
rect -4404 25543 -4402 25563
rect -4308 25543 -4306 25563
rect -4260 25543 -4258 25563
rect -4164 25543 -4162 25563
rect -4020 25543 -4018 25563
rect -3876 25543 -3874 25563
rect -3732 25543 -3730 25563
rect -3588 25544 -3586 25563
rect -3599 25543 -3565 25544
rect -3564 25543 -3562 25563
rect -3516 25543 -3514 25563
rect -3492 25544 -3490 25563
rect -3503 25543 -3469 25544
rect -3468 25543 -3466 25563
rect -3420 25543 -3418 25563
rect -3324 25543 -3322 25563
rect -3228 25543 -3226 25563
rect -3132 25543 -3130 25563
rect -3012 25543 -3010 25563
rect -2964 25543 -2962 25563
rect -2916 25543 -2914 25563
rect -2892 25543 -2890 25563
rect -2868 25543 -2866 25563
rect -2820 25543 -2818 25563
rect -2796 25543 -2794 25563
rect -2772 25543 -2770 25563
rect -2676 25543 -2674 25563
rect -2580 25543 -2578 25563
rect -2364 25543 -2362 25563
rect -2316 25543 -2314 25563
rect -2268 25543 -2266 25563
rect -2244 25543 -2242 25563
rect -2172 25543 -2170 25563
rect -2148 25543 -2146 25563
rect -2076 25543 -2074 25563
rect -2052 25543 -2050 25563
rect -1980 25543 -1978 25563
rect -1884 25543 -1882 25563
rect -1572 25543 -1570 25563
rect -1476 25543 -1474 25563
rect -1380 25543 -1378 25563
rect -1356 25543 -1354 25563
rect -1308 25543 -1306 25563
rect -1260 25543 -1258 25563
rect -1140 25543 -1138 25563
rect -708 25543 -706 25563
rect -612 25543 -610 25563
rect -588 25543 -586 25563
rect -540 25543 -538 25563
rect -492 25543 -490 25563
rect -444 25543 -442 25563
rect -396 25543 -394 25563
rect -300 25543 -298 25563
rect -276 25543 -274 25563
rect -228 25543 -226 25563
rect -12 25543 -10 25563
rect 156 25543 158 25563
rect 204 25543 206 25563
rect 252 25543 254 25563
rect 348 25543 350 25563
rect 468 25543 470 25563
rect 492 25543 494 25563
rect 564 25543 566 25563
rect 588 25543 590 25563
rect 636 25543 638 25563
rect 660 25543 662 25563
rect 732 25543 734 25563
rect 1092 25543 1094 25563
rect 1308 25543 1310 25563
rect 1332 25543 1334 25563
rect 1380 25543 1382 25563
rect 1428 25543 1430 25563
rect 1476 25543 1478 25563
rect 1644 25543 1646 25563
rect 1692 25543 1694 25563
rect 1740 25543 1742 25563
rect 1788 25543 1790 25563
rect 2028 25543 2030 25563
rect 2076 25543 2078 25563
rect 2100 25543 2102 25563
rect 2124 25543 2126 25563
rect 2172 25543 2174 25563
rect 2220 25543 2222 25563
rect 2316 25543 2318 25563
rect 2412 25543 2414 25563
rect 2460 25543 2462 25563
rect 2508 25543 2510 25563
rect 2580 25543 2582 25563
rect 2604 25543 2606 25563
rect 2676 25543 2678 25563
rect 2700 25543 2702 25563
rect 2748 25543 2750 25563
rect 2772 25543 2774 25563
rect 2796 25543 2798 25563
rect 2844 25543 2846 25563
rect 2868 25543 2870 25563
rect 2892 25543 2894 25563
rect 2940 25543 2942 25563
rect 3012 25543 3014 25563
rect 3108 25543 3110 25563
rect 3252 25543 3254 25563
rect 3348 25543 3350 25563
rect 3396 25543 3398 25563
rect 3564 25543 3566 25563
rect 3636 25543 3638 25563
rect 3660 25543 3662 25563
rect 3732 25543 3734 25563
rect 3828 25543 3830 25563
rect 3924 25543 3926 25563
rect 4020 25543 4022 25563
rect 4044 25543 4046 25563
rect 4092 25543 4094 25563
rect 4116 25544 4118 25563
rect 4105 25543 4139 25544
rect 4140 25543 4142 25563
rect 4188 25543 4190 25563
rect 4212 25543 4214 25563
rect 4236 25543 4238 25563
rect 4308 25543 4310 25563
rect 4332 25543 4334 25563
rect 4404 25543 4406 25563
rect 4500 25543 4502 25563
rect 4596 25543 4598 25563
rect 4692 25543 4694 25563
rect 4860 25543 4862 25563
rect 4956 25543 4958 25563
rect 4980 25543 4982 25563
rect 5004 25543 5006 25563
rect 5052 25543 5054 25563
rect 5100 25543 5102 25563
rect 5124 25543 5126 25563
rect 5220 25543 5222 25563
rect 5268 25543 5270 25563
rect 5388 25543 5390 25563
rect 5484 25543 5486 25563
rect 5508 25543 5510 25563
rect 5532 25543 5534 25563
rect 5628 25543 5630 25563
rect 5652 25543 5654 25563
rect 5748 25543 5750 25563
rect 5796 25543 5798 25563
rect 5844 25543 5846 25563
rect 5892 25543 5894 25563
rect 6132 25543 6134 25563
rect 6180 25543 6182 25563
rect 6228 25543 6230 25563
rect 6252 25543 6254 25563
rect 6276 25543 6278 25563
rect 6324 25543 6326 25563
rect 6372 25543 6374 25563
rect 6492 25543 6494 25563
rect 6588 25543 6590 25563
rect 6612 25543 6614 25563
rect 6660 25543 6662 25563
rect 6684 25543 6686 25563
rect 6708 25543 6710 25563
rect 6780 25543 6782 25563
rect 6804 25543 6806 25563
rect 6900 25543 6902 25563
rect 6924 25543 6926 25563
rect 7020 25543 7022 25563
rect 7068 25543 7070 25563
rect 7164 25543 7166 25563
rect 7236 25543 7238 25563
rect 7332 25543 7334 25563
rect 7380 25543 7382 25563
rect 7428 25543 7430 25563
rect 7452 25543 7454 25563
rect 7476 25543 7478 25563
rect 7524 25543 7526 25563
rect 7548 25543 7550 25563
rect 7572 25543 7574 25563
rect 7620 25543 7622 25563
rect 7644 25543 7646 25563
rect 7668 25543 7670 25563
rect 7788 25543 7790 25563
rect 7884 25543 7886 25563
rect 7956 25543 7958 25563
rect 7980 25543 7982 25563
rect 8028 25543 8030 25563
rect 8196 25543 8198 25563
rect 8244 25543 8246 25563
rect 8268 25543 8270 25563
rect 8292 25543 8294 25563
rect 8340 25543 8342 25563
rect 8364 25543 8366 25563
rect 8388 25543 8390 25563
rect 8436 25543 8438 25563
rect 8604 25560 8606 25563
rect 8604 25543 8607 25560
rect 8652 25543 8654 25563
rect 8700 25543 8702 25563
rect 8724 25560 8726 25563
rect 8724 25543 8727 25560
rect 8748 25543 8750 25563
rect 8820 25543 8822 25563
rect 8844 25543 8846 25563
rect 8868 25543 8870 25563
rect 9516 25543 9518 25563
rect 9612 25544 9614 25563
rect 9601 25543 9635 25544
rect 9660 25543 9662 25563
rect 9684 25543 9686 25563
rect 9708 25543 9710 25563
rect 9756 25543 9758 25563
rect 9780 25543 9782 25563
rect 9804 25543 9806 25563
rect 9852 25543 9854 25563
rect 9900 25543 9902 25563
rect 9948 25543 9950 25563
rect 9996 25543 9998 25563
rect 10068 25543 10070 25563
rect 10092 25543 10094 25563
rect 10116 25543 10118 25563
rect 10164 25543 10166 25563
rect 10188 25543 10190 25563
rect 10212 25543 10214 25563
rect 10284 25543 10286 25563
rect 10308 25543 10310 25563
rect 10332 25543 10334 25563
rect 10380 25543 10382 25563
rect 10404 25543 10406 25563
rect 10428 25543 10430 25563
rect 10476 25543 10478 25563
rect 10500 25543 10502 25563
rect 10524 25543 10526 25563
rect 10572 25543 10574 25563
rect 10596 25543 10598 25563
rect 10620 25543 10622 25563
rect 10668 25543 10670 25563
rect 10692 25543 10694 25563
rect 10716 25543 10718 25563
rect 10788 25543 10790 25563
rect 10836 25560 10838 25563
rect 10836 25543 10839 25560
rect 10956 25543 10958 25563
rect 11004 25543 11006 25563
rect 11052 25543 11054 25563
rect 11100 25543 11102 25563
rect 11172 25543 11174 25563
rect 11220 25543 11222 25563
rect 11340 25543 11342 25563
rect 11436 25543 11438 25563
rect 11532 25543 11534 25563
rect 11580 25543 11582 25563
rect 11628 25543 11630 25563
rect 11676 25543 11678 25563
rect 11724 25543 11726 25563
rect 11772 25543 11774 25563
rect 11796 25543 11798 25563
rect 11892 25543 11894 25563
rect 11988 25543 11990 25563
rect 12060 25543 12062 25563
rect 12132 25543 12134 25563
rect 12228 25543 12230 25563
rect 12276 25543 12278 25563
rect 12324 25543 12326 25563
rect 12420 25543 12422 25563
rect 12444 25543 12446 25563
rect 12492 25543 12494 25563
rect 12516 25543 12518 25563
rect 12540 25543 12542 25563
rect 12588 25543 12590 25563
rect 12636 25543 12638 25563
rect 12732 25543 12734 25563
rect 12756 25543 12758 25563
rect 12804 25543 12806 25563
rect 12828 25543 12830 25563
rect 12852 25543 12854 25563
rect 12948 25543 12950 25563
rect 12972 25543 12974 25563
rect 13044 25543 13046 25563
rect 13068 25543 13070 25563
rect 13116 25543 13118 25563
rect 13284 25543 13286 25563
rect 13332 25543 13334 25563
rect 13572 25543 13574 25563
rect 13620 25543 13622 25563
rect 13668 25543 13670 25563
rect 13716 25543 13718 25563
rect 13764 25543 13766 25563
rect 13860 25543 13862 25563
rect 13956 25543 13958 25563
rect 14004 25543 14006 25563
rect 14100 25543 14102 25563
rect 15180 25543 15182 25563
rect 15276 25543 15278 25563
rect 15420 25543 15422 25563
rect 15492 25543 15494 25563
rect 15660 25543 15662 25563
rect 15708 25543 15710 25563
rect 15732 25543 15734 25563
rect 15756 25543 15758 25563
rect 15804 25543 15806 25563
rect 15828 25543 15830 25563
rect 15852 25543 15854 25563
rect 15900 25543 15902 25563
rect 15948 25543 15950 25563
rect 16044 25543 16046 25563
rect 16068 25543 16070 25563
rect 16164 25543 16166 25563
rect 16260 25543 16262 25563
rect 16308 25543 16310 25563
rect 16332 25543 16334 25563
rect 16356 25543 16358 25563
rect 16404 25543 16406 25563
rect 16452 25543 16454 25563
rect 16548 25543 16550 25563
rect 16572 25543 16574 25563
rect 16620 25543 16622 25563
rect 16668 25543 16670 25563
rect 16716 25543 16718 25563
rect 16764 25543 16766 25563
rect 16812 25543 16814 25563
rect 16884 25543 16886 25563
rect 16908 25543 16910 25563
rect 16980 25543 16982 25563
rect 17052 25543 17054 25563
rect 17196 25543 17198 25563
rect 17220 25543 17222 25563
rect 17292 25543 17294 25563
rect 17316 25543 17318 25563
rect 18084 25543 18086 25563
rect 18132 25543 18134 25563
rect 18228 25543 18230 25563
rect 18396 25543 18398 25563
rect 18492 25543 18494 25563
rect 18516 25543 18518 25563
rect 18564 25543 18566 25563
rect 18612 25543 18614 25563
rect 18660 25543 18662 25563
rect 18756 25543 18758 25563
rect 18852 25543 18854 25563
rect 18900 25543 18902 25563
rect 18996 25543 18998 25563
rect 19020 25543 19022 25563
rect 19092 25543 19094 25563
rect 19116 25543 19118 25563
rect 19140 25543 19142 25563
rect 19188 25543 19190 25563
rect 19236 25543 19238 25563
rect 19332 25543 19334 25563
rect 19476 25543 19478 25563
rect 19788 25543 19790 25563
rect 19836 25543 19838 25563
rect 19860 25543 19862 25563
rect 19884 25543 19886 25563
rect 19932 25543 19934 25563
rect 19956 25543 19958 25563
rect 19980 25543 19982 25563
rect 20028 25543 20030 25563
rect 20052 25543 20054 25563
rect 20076 25543 20078 25563
rect 20148 25543 20150 25563
rect 20172 25543 20174 25563
rect 20196 25543 20198 25563
rect 20268 25543 20270 25563
rect 20292 25543 20294 25563
rect 20388 25543 20390 25563
rect 20412 25543 20414 25563
rect 20508 25543 20510 25563
rect 20556 25543 20558 25563
rect 20604 25543 20606 25563
rect 20916 25543 20918 25563
rect 20964 25543 20966 25563
rect 21012 25543 21014 25563
rect 21060 25543 21062 25563
rect 21108 25543 21110 25563
rect 21204 25543 21206 25563
rect 21300 25543 21302 25563
rect 21324 25543 21326 25563
rect 21444 25543 21446 25563
rect 21468 25543 21470 25563
rect 21564 25543 21566 25563
rect 21588 25543 21590 25563
rect 21684 25543 21686 25563
rect 21708 25543 21710 25563
rect 21828 25543 21830 25563
rect 21924 25543 21926 25563
rect 22068 25543 22070 25563
rect 22188 25543 22190 25563
rect 22212 25543 22214 25563
rect 22884 25543 22886 25563
rect 22980 25543 22982 25563
rect 23076 25543 23078 25563
rect 23100 25543 23102 25563
rect 23124 25543 23126 25563
rect 23244 25543 23246 25563
rect 23340 25543 23342 25563
rect 23412 25543 23414 25563
rect 23439 25560 23453 25563
rect 23460 25563 25859 25567
rect 23460 25560 23477 25563
rect 23460 25543 23462 25560
rect 23508 25543 23510 25563
rect 23556 25543 23558 25563
rect 23604 25543 23606 25563
rect 23652 25543 23654 25563
rect 23676 25543 23678 25563
rect 23772 25543 23774 25563
rect 23820 25543 23822 25563
rect 23916 25543 23918 25563
rect 24012 25543 24014 25563
rect 24060 25543 24062 25563
rect 24156 25543 24158 25563
rect 24492 25543 24494 25563
rect 24516 25543 24518 25563
rect 24588 25543 24590 25563
rect 24612 25543 24614 25563
rect 24684 25543 24686 25563
rect 24732 25543 24734 25563
rect 24756 25543 24758 25563
rect 24780 25543 24782 25563
rect 24852 25543 24854 25563
rect 24876 25543 24878 25563
rect 24972 25543 24974 25563
rect 25068 25543 25070 25563
rect 25164 25543 25166 25563
rect 25260 25543 25262 25563
rect 25284 25543 25286 25563
rect 25356 25543 25358 25563
rect 25380 25543 25382 25563
rect 25404 25543 25406 25563
rect 25500 25543 25502 25563
rect 25596 25543 25598 25563
rect 25777 25543 25811 25544
rect -15455 25539 25811 25543
rect -15335 25519 -15301 25520
rect -15108 25519 -15106 25539
rect -14892 25519 -14890 25539
rect -14745 25536 -14731 25539
rect -14676 25519 -14674 25539
rect -14495 25519 -14413 25520
rect -14340 25519 -14338 25539
rect -13788 25519 -13786 25539
rect -13428 25519 -13426 25539
rect -12756 25519 -12754 25539
rect -12660 25519 -12658 25539
rect -12492 25536 -12490 25539
rect -12492 25520 -12489 25536
rect -12527 25519 -12469 25520
rect -12396 25519 -12394 25539
rect -12348 25519 -12346 25539
rect -12252 25519 -12250 25539
rect -12156 25519 -12154 25539
rect -12060 25519 -12058 25539
rect -11844 25519 -11842 25539
rect -11676 25519 -11674 25539
rect -11508 25519 -11506 25539
rect -11436 25519 -11434 25539
rect -11412 25519 -11410 25539
rect -11340 25519 -11338 25539
rect -11196 25519 -11194 25539
rect -11100 25519 -11098 25539
rect -10740 25519 -10738 25539
rect -10644 25519 -10642 25539
rect -9996 25519 -9994 25539
rect -9900 25519 -9898 25539
rect -9732 25519 -9730 25539
rect -9516 25519 -9514 25539
rect -9468 25519 -9466 25539
rect -9348 25519 -9346 25539
rect -9180 25519 -9178 25539
rect -8604 25519 -8602 25539
rect -8436 25519 -8434 25539
rect -8409 25536 -8395 25539
rect -8388 25536 -8385 25539
rect -8364 25519 -8362 25539
rect -8340 25519 -8338 25539
rect -8268 25519 -8266 25539
rect -8100 25519 -8098 25539
rect -8052 25520 -8050 25539
rect -8063 25519 -8029 25520
rect -8004 25519 -8002 25539
rect -7932 25519 -7930 25539
rect -7692 25520 -7690 25539
rect -7703 25519 -7669 25520
rect -7620 25519 -7618 25539
rect -7524 25519 -7522 25539
rect -7356 25519 -7354 25539
rect -7308 25519 -7306 25539
rect -7212 25519 -7210 25539
rect -7079 25519 -7045 25520
rect -7044 25519 -7042 25539
rect -6983 25534 -6980 25539
rect -6972 25534 -6970 25539
rect -6973 25520 -6970 25534
rect -6948 25519 -6946 25539
rect -6876 25536 -6874 25539
rect -6876 25519 -6873 25536
rect -6852 25519 -6850 25539
rect -6780 25519 -6778 25539
rect -6756 25519 -6754 25539
rect -6660 25519 -6658 25539
rect -6612 25519 -6610 25539
rect -6599 25519 -6565 25520
rect -6516 25519 -6514 25539
rect -6372 25519 -6370 25539
rect -6156 25519 -6154 25539
rect -6060 25519 -6058 25539
rect -6036 25519 -6034 25539
rect -5892 25519 -5890 25539
rect -5268 25519 -5266 25539
rect -5196 25519 -5194 25539
rect -5172 25519 -5170 25539
rect -5100 25519 -5098 25539
rect -5076 25519 -5074 25539
rect -4980 25519 -4978 25539
rect -4956 25519 -4954 25539
rect -4860 25519 -4858 25539
rect -4644 25519 -4642 25539
rect -4500 25519 -4498 25539
rect -4473 25536 -4459 25539
rect -4404 25519 -4402 25539
rect -4308 25519 -4306 25539
rect -4260 25519 -4258 25539
rect -4164 25519 -4162 25539
rect -4020 25519 -4018 25539
rect -3876 25519 -3874 25539
rect -3732 25519 -3730 25539
rect -3599 25534 -3596 25539
rect -3588 25534 -3586 25539
rect -3589 25520 -3586 25534
rect -3564 25519 -3562 25539
rect -3516 25519 -3514 25539
rect -3503 25534 -3500 25539
rect -3492 25536 -3490 25539
rect -3492 25534 -3489 25536
rect -3493 25520 -3489 25534
rect -3468 25519 -3466 25539
rect -3420 25519 -3418 25539
rect -3324 25519 -3322 25539
rect -3228 25519 -3226 25539
rect -3132 25519 -3130 25539
rect -3012 25519 -3010 25539
rect -2964 25519 -2962 25539
rect -2916 25519 -2914 25539
rect -2892 25519 -2890 25539
rect -2868 25519 -2866 25539
rect -2820 25519 -2818 25539
rect -2796 25519 -2794 25539
rect -2772 25519 -2770 25539
rect -2676 25519 -2674 25539
rect -2580 25519 -2578 25539
rect -2364 25519 -2362 25539
rect -2316 25519 -2314 25539
rect -2268 25519 -2266 25539
rect -2244 25519 -2242 25539
rect -2172 25519 -2170 25539
rect -2148 25519 -2146 25539
rect -2076 25519 -2074 25539
rect -2052 25519 -2050 25539
rect -1980 25519 -1978 25539
rect -1884 25519 -1882 25539
rect -1572 25519 -1570 25539
rect -1476 25519 -1474 25539
rect -1380 25519 -1378 25539
rect -1356 25519 -1354 25539
rect -1308 25519 -1306 25539
rect -1260 25519 -1258 25539
rect -1140 25519 -1138 25539
rect -708 25519 -706 25539
rect -612 25519 -610 25539
rect -588 25519 -586 25539
rect -540 25519 -538 25539
rect -492 25519 -490 25539
rect -444 25519 -442 25539
rect -396 25519 -394 25539
rect -300 25519 -298 25539
rect -276 25519 -274 25539
rect -228 25519 -226 25539
rect -12 25519 -10 25539
rect 156 25519 158 25539
rect 204 25519 206 25539
rect 252 25519 254 25539
rect 348 25519 350 25539
rect 468 25519 470 25539
rect 492 25519 494 25539
rect 564 25519 566 25539
rect 588 25519 590 25539
rect 636 25519 638 25539
rect 660 25519 662 25539
rect 732 25519 734 25539
rect 1092 25519 1094 25539
rect 1308 25519 1310 25539
rect 1332 25519 1334 25539
rect 1380 25519 1382 25539
rect 1428 25519 1430 25539
rect 1476 25519 1478 25539
rect 1644 25519 1646 25539
rect 1692 25519 1694 25539
rect 1740 25519 1742 25539
rect 1788 25519 1790 25539
rect 2028 25519 2030 25539
rect 2076 25519 2078 25539
rect 2100 25519 2102 25539
rect 2124 25519 2126 25539
rect 2172 25519 2174 25539
rect 2220 25519 2222 25539
rect 2316 25519 2318 25539
rect 2412 25519 2414 25539
rect 2460 25519 2462 25539
rect 2508 25519 2510 25539
rect 2580 25519 2582 25539
rect 2604 25519 2606 25539
rect 2676 25519 2678 25539
rect 2700 25519 2702 25539
rect 2748 25519 2750 25539
rect 2772 25519 2774 25539
rect 2796 25519 2798 25539
rect 2844 25519 2846 25539
rect 2868 25519 2870 25539
rect 2892 25519 2894 25539
rect 2940 25519 2942 25539
rect 3012 25519 3014 25539
rect 3108 25519 3110 25539
rect 3252 25519 3254 25539
rect 3348 25519 3350 25539
rect 3396 25519 3398 25539
rect 3564 25519 3566 25539
rect 3636 25519 3638 25539
rect 3660 25519 3662 25539
rect 3732 25519 3734 25539
rect 3828 25519 3830 25539
rect 3924 25519 3926 25539
rect 4020 25519 4022 25539
rect 4044 25519 4046 25539
rect 4092 25519 4094 25539
rect 4105 25534 4108 25539
rect 4116 25534 4118 25539
rect 4115 25520 4118 25534
rect 4140 25519 4142 25539
rect 4188 25519 4190 25539
rect 4212 25536 4214 25539
rect 4212 25519 4215 25536
rect 4236 25519 4238 25539
rect 4308 25519 4310 25539
rect 4332 25519 4334 25539
rect 4404 25519 4406 25539
rect 4500 25519 4502 25539
rect 4596 25519 4598 25539
rect 4692 25519 4694 25539
rect 4860 25519 4862 25539
rect 4956 25519 4958 25539
rect 4980 25519 4982 25539
rect 5004 25520 5006 25539
rect 4993 25519 5027 25520
rect 5052 25519 5054 25539
rect 5100 25519 5102 25539
rect 5124 25519 5126 25539
rect 5220 25519 5222 25539
rect 5268 25519 5270 25539
rect 5388 25519 5390 25539
rect 5484 25519 5486 25539
rect 5508 25519 5510 25539
rect 5532 25519 5534 25539
rect 5628 25519 5630 25539
rect 5652 25519 5654 25539
rect 5748 25519 5750 25539
rect 5796 25519 5798 25539
rect 5844 25519 5846 25539
rect 5892 25519 5894 25539
rect 6132 25519 6134 25539
rect 6180 25519 6182 25539
rect 6228 25519 6230 25539
rect 6252 25519 6254 25539
rect 6276 25519 6278 25539
rect 6324 25519 6326 25539
rect 6372 25519 6374 25539
rect 6492 25519 6494 25539
rect 6588 25519 6590 25539
rect 6612 25519 6614 25539
rect 6660 25519 6662 25539
rect 6684 25519 6686 25539
rect 6708 25519 6710 25539
rect 6780 25519 6782 25539
rect 6804 25519 6806 25539
rect 6900 25519 6902 25539
rect 6924 25519 6926 25539
rect 7020 25519 7022 25539
rect 7068 25519 7070 25539
rect 7164 25519 7166 25539
rect 7236 25519 7238 25539
rect 7332 25519 7334 25539
rect 7380 25519 7382 25539
rect 7428 25519 7430 25539
rect 7452 25519 7454 25539
rect 7476 25519 7478 25539
rect 7524 25519 7526 25539
rect 7548 25519 7550 25539
rect 7572 25519 7574 25539
rect 7620 25519 7622 25539
rect 7644 25519 7646 25539
rect 7668 25519 7670 25539
rect 7788 25520 7790 25539
rect 7777 25519 7811 25520
rect 7884 25519 7886 25539
rect 7956 25519 7958 25539
rect 7980 25519 7982 25539
rect 8028 25519 8030 25539
rect 8113 25519 8171 25520
rect 8196 25519 8198 25539
rect 8244 25519 8246 25539
rect 8268 25519 8270 25539
rect 8292 25519 8294 25539
rect 8340 25519 8342 25539
rect 8364 25519 8366 25539
rect 8388 25519 8390 25539
rect 8436 25519 8438 25539
rect 8583 25536 8597 25539
rect 8604 25536 8607 25539
rect 8652 25519 8654 25539
rect 8700 25519 8702 25539
rect 8703 25536 8717 25539
rect 8724 25536 8727 25539
rect 8748 25519 8750 25539
rect 8820 25519 8822 25539
rect 8844 25519 8846 25539
rect 8868 25519 8870 25539
rect 9516 25519 9518 25539
rect 9601 25534 9604 25539
rect 9612 25534 9614 25539
rect 9611 25520 9614 25534
rect 9660 25519 9662 25539
rect 9684 25519 9686 25539
rect 9708 25536 9710 25539
rect 9708 25519 9711 25536
rect 9756 25519 9758 25539
rect 9780 25519 9782 25539
rect 9804 25519 9806 25539
rect 9852 25519 9854 25539
rect 9900 25519 9902 25539
rect 9948 25519 9950 25539
rect 9996 25519 9998 25539
rect 10068 25519 10070 25539
rect 10092 25519 10094 25539
rect 10116 25519 10118 25539
rect 10164 25519 10166 25539
rect 10188 25519 10190 25539
rect 10212 25519 10214 25539
rect 10284 25519 10286 25539
rect 10308 25519 10310 25539
rect 10332 25519 10334 25539
rect 10380 25519 10382 25539
rect 10404 25519 10406 25539
rect 10428 25519 10430 25539
rect 10476 25519 10478 25539
rect 10500 25519 10502 25539
rect 10524 25519 10526 25539
rect 10572 25519 10574 25539
rect 10596 25519 10598 25539
rect 10620 25519 10622 25539
rect 10668 25519 10670 25539
rect 10692 25519 10694 25539
rect 10716 25519 10718 25539
rect 10788 25519 10790 25539
rect 10815 25536 10829 25539
rect 10836 25536 10839 25539
rect 10956 25519 10958 25539
rect 11004 25519 11006 25539
rect 11052 25519 11054 25539
rect 11100 25519 11102 25539
rect 11172 25519 11174 25539
rect 11220 25519 11222 25539
rect 11340 25519 11342 25539
rect 11436 25519 11438 25539
rect 11532 25519 11534 25539
rect 11580 25519 11582 25539
rect 11628 25519 11630 25539
rect 11676 25519 11678 25539
rect 11724 25519 11726 25539
rect 11772 25519 11774 25539
rect 11796 25519 11798 25539
rect 11892 25519 11894 25539
rect 11988 25519 11990 25539
rect 12060 25519 12062 25539
rect 12132 25519 12134 25539
rect 12228 25519 12230 25539
rect 12276 25519 12278 25539
rect 12324 25519 12326 25539
rect 12420 25519 12422 25539
rect 12444 25519 12446 25539
rect 12492 25519 12494 25539
rect 12516 25519 12518 25539
rect 12540 25519 12542 25539
rect 12588 25519 12590 25539
rect 12636 25519 12638 25539
rect 12732 25519 12734 25539
rect 12756 25519 12758 25539
rect 12804 25519 12806 25539
rect 12828 25519 12830 25539
rect 12852 25519 12854 25539
rect 12948 25519 12950 25539
rect 12972 25519 12974 25539
rect 13044 25519 13046 25539
rect 13068 25519 13070 25539
rect 13116 25519 13118 25539
rect 13284 25519 13286 25539
rect 13332 25519 13334 25539
rect 13572 25519 13574 25539
rect 13620 25519 13622 25539
rect 13668 25519 13670 25539
rect 13716 25519 13718 25539
rect 13764 25519 13766 25539
rect 13860 25519 13862 25539
rect 13956 25519 13958 25539
rect 14004 25519 14006 25539
rect 14100 25519 14102 25539
rect 15180 25519 15182 25539
rect 15276 25519 15278 25539
rect 15420 25519 15422 25539
rect 15492 25519 15494 25539
rect 15660 25519 15662 25539
rect 15708 25519 15710 25539
rect 15732 25519 15734 25539
rect 15756 25519 15758 25539
rect 15804 25519 15806 25539
rect 15828 25519 15830 25539
rect 15852 25519 15854 25539
rect 15900 25519 15902 25539
rect 15948 25519 15950 25539
rect 16044 25519 16046 25539
rect 16068 25519 16070 25539
rect 16164 25519 16166 25539
rect 16260 25519 16262 25539
rect 16308 25519 16310 25539
rect 16332 25519 16334 25539
rect 16356 25519 16358 25539
rect 16404 25519 16406 25539
rect 16452 25519 16454 25539
rect 16548 25519 16550 25539
rect 16572 25519 16574 25539
rect 16620 25519 16622 25539
rect 16668 25519 16670 25539
rect 16716 25519 16718 25539
rect 16764 25519 16766 25539
rect 16812 25519 16814 25539
rect 16884 25519 16886 25539
rect 16908 25519 16910 25539
rect 16980 25519 16982 25539
rect 17052 25519 17054 25539
rect 17196 25519 17198 25539
rect 17220 25519 17222 25539
rect 17292 25519 17294 25539
rect 17316 25519 17318 25539
rect 18084 25519 18086 25539
rect 18132 25519 18134 25539
rect 18228 25519 18230 25539
rect 18396 25519 18398 25539
rect 18492 25519 18494 25539
rect 18516 25519 18518 25539
rect 18564 25519 18566 25539
rect 18612 25519 18614 25539
rect 18660 25519 18662 25539
rect 18756 25519 18758 25539
rect 18852 25519 18854 25539
rect 18900 25519 18902 25539
rect 18996 25519 18998 25539
rect 19020 25519 19022 25539
rect 19092 25519 19094 25539
rect 19116 25519 19118 25539
rect 19140 25519 19142 25539
rect 19188 25519 19190 25539
rect 19236 25519 19238 25539
rect 19332 25519 19334 25539
rect 19476 25519 19478 25539
rect 19788 25519 19790 25539
rect 19836 25519 19838 25539
rect 19860 25519 19862 25539
rect 19884 25519 19886 25539
rect 19932 25519 19934 25539
rect 19956 25519 19958 25539
rect 19980 25519 19982 25539
rect 20028 25519 20030 25539
rect 20052 25519 20054 25539
rect 20076 25519 20078 25539
rect 20148 25519 20150 25539
rect 20172 25519 20174 25539
rect 20196 25519 20198 25539
rect 20268 25519 20270 25539
rect 20292 25519 20294 25539
rect 20388 25519 20390 25539
rect 20412 25519 20414 25539
rect 20508 25519 20510 25539
rect 20556 25519 20558 25539
rect 20604 25519 20606 25539
rect 20916 25519 20918 25539
rect 20964 25519 20966 25539
rect 21012 25519 21014 25539
rect 21060 25519 21062 25539
rect 21108 25519 21110 25539
rect 21204 25519 21206 25539
rect 21300 25519 21302 25539
rect 21324 25519 21326 25539
rect 21444 25519 21446 25539
rect 21468 25519 21470 25539
rect 21564 25519 21566 25539
rect 21588 25519 21590 25539
rect 21684 25519 21686 25539
rect 21708 25519 21710 25539
rect 21828 25519 21830 25539
rect 21924 25519 21926 25539
rect 22068 25519 22070 25539
rect 22188 25519 22190 25539
rect 22212 25519 22214 25539
rect 22884 25519 22886 25539
rect 22980 25519 22982 25539
rect 23076 25519 23078 25539
rect 23100 25519 23102 25539
rect 23124 25519 23126 25539
rect 23244 25519 23246 25539
rect 23340 25519 23342 25539
rect 23412 25519 23414 25539
rect 23460 25519 23462 25539
rect 23508 25519 23510 25539
rect 23556 25519 23558 25539
rect 23604 25519 23606 25539
rect 23652 25519 23654 25539
rect 23676 25519 23678 25539
rect 23772 25519 23774 25539
rect 23820 25519 23822 25539
rect 23916 25519 23918 25539
rect 24012 25519 24014 25539
rect 24060 25519 24062 25539
rect 24156 25519 24158 25539
rect 24492 25519 24494 25539
rect 24516 25519 24518 25539
rect 24588 25519 24590 25539
rect 24612 25519 24614 25539
rect 24684 25519 24686 25539
rect 24732 25519 24734 25539
rect 24756 25519 24758 25539
rect 24780 25519 24782 25539
rect 24852 25519 24854 25539
rect 24876 25519 24878 25539
rect 24972 25519 24974 25539
rect 25068 25519 25070 25539
rect 25164 25519 25166 25539
rect 25260 25519 25262 25539
rect 25284 25519 25286 25539
rect 25356 25519 25358 25539
rect 25380 25519 25382 25539
rect 25404 25519 25406 25539
rect 25500 25519 25502 25539
rect 25596 25519 25598 25539
rect 25633 25519 25667 25520
rect -15335 25515 25667 25519
rect -15215 25495 -15181 25496
rect -15108 25495 -15106 25515
rect -14892 25495 -14890 25515
rect -14676 25495 -14674 25515
rect -14471 25510 -14468 25515
rect -14340 25512 -14338 25515
rect -14461 25496 -14458 25510
rect -14460 25495 -14458 25496
rect -14340 25495 -14337 25512
rect -13788 25495 -13786 25515
rect -13463 25495 -13429 25496
rect -13428 25495 -13426 25515
rect -12756 25495 -12754 25515
rect -12660 25495 -12658 25515
rect -12513 25512 -12499 25515
rect -12492 25512 -12489 25515
rect -12396 25512 -12394 25515
rect -12396 25495 -12393 25512
rect -12348 25495 -12346 25515
rect -12252 25495 -12250 25515
rect -12156 25495 -12154 25515
rect -12060 25495 -12058 25515
rect -11844 25495 -11842 25515
rect -11676 25495 -11674 25515
rect -11508 25495 -11506 25515
rect -11436 25495 -11434 25515
rect -11412 25495 -11410 25515
rect -11340 25495 -11338 25515
rect -11196 25495 -11194 25515
rect -11100 25495 -11098 25515
rect -10871 25495 -10813 25496
rect -10740 25495 -10738 25515
rect -10644 25495 -10642 25515
rect -9996 25495 -9994 25515
rect -9900 25495 -9898 25515
rect -9732 25495 -9730 25515
rect -9575 25495 -9541 25496
rect -9516 25495 -9514 25515
rect -9468 25495 -9466 25515
rect -9348 25495 -9346 25515
rect -9180 25495 -9178 25515
rect -8735 25495 -8677 25496
rect -8604 25495 -8602 25515
rect -8436 25495 -8434 25515
rect -8364 25495 -8362 25515
rect -8340 25495 -8338 25515
rect -8268 25495 -8266 25515
rect -8100 25495 -8098 25515
rect -8063 25510 -8060 25515
rect -8052 25510 -8050 25515
rect -8053 25496 -8050 25510
rect -8004 25495 -8002 25515
rect -7932 25495 -7930 25515
rect -7703 25510 -7700 25515
rect -7692 25510 -7690 25515
rect -7693 25496 -7690 25510
rect -7620 25495 -7618 25515
rect -7524 25495 -7522 25515
rect -7356 25495 -7354 25515
rect -7308 25495 -7306 25515
rect -7212 25495 -7210 25515
rect -7044 25495 -7042 25515
rect -6948 25495 -6946 25515
rect -6897 25512 -6883 25515
rect -6876 25512 -6873 25515
rect -6852 25495 -6850 25515
rect -6780 25495 -6778 25515
rect -6756 25495 -6754 25515
rect -6660 25495 -6658 25515
rect -6612 25495 -6610 25515
rect -6516 25495 -6514 25515
rect -6372 25495 -6370 25515
rect -6156 25495 -6154 25515
rect -6060 25495 -6058 25515
rect -6036 25495 -6034 25515
rect -5892 25495 -5890 25515
rect -5268 25495 -5266 25515
rect -5196 25495 -5194 25515
rect -5172 25495 -5170 25515
rect -5100 25495 -5098 25515
rect -5076 25495 -5074 25515
rect -4980 25495 -4978 25515
rect -4956 25495 -4954 25515
rect -4860 25495 -4858 25515
rect -4644 25495 -4642 25515
rect -4500 25495 -4498 25515
rect -4404 25495 -4402 25515
rect -4308 25495 -4306 25515
rect -4260 25495 -4258 25515
rect -4164 25495 -4162 25515
rect -4020 25495 -4018 25515
rect -3876 25495 -3874 25515
rect -3732 25495 -3730 25515
rect -3564 25495 -3562 25515
rect -3516 25495 -3514 25515
rect -3513 25512 -3499 25515
rect -3468 25495 -3466 25515
rect -3420 25495 -3418 25515
rect -3417 25512 -3403 25515
rect -3324 25495 -3322 25515
rect -3228 25495 -3226 25515
rect -3132 25495 -3130 25515
rect -3012 25495 -3010 25515
rect -2964 25495 -2962 25515
rect -2916 25495 -2914 25515
rect -2892 25495 -2890 25515
rect -2868 25495 -2866 25515
rect -2820 25495 -2818 25515
rect -2796 25495 -2794 25515
rect -2772 25495 -2770 25515
rect -2676 25495 -2674 25515
rect -2580 25495 -2578 25515
rect -2364 25495 -2362 25515
rect -2316 25495 -2314 25515
rect -2268 25495 -2266 25515
rect -2244 25495 -2242 25515
rect -2172 25495 -2170 25515
rect -2148 25495 -2146 25515
rect -2076 25495 -2074 25515
rect -2052 25495 -2050 25515
rect -1980 25495 -1978 25515
rect -1884 25495 -1882 25515
rect -1572 25495 -1570 25515
rect -1476 25495 -1474 25515
rect -1380 25495 -1378 25515
rect -1356 25495 -1354 25515
rect -1308 25495 -1306 25515
rect -1260 25495 -1258 25515
rect -1140 25495 -1138 25515
rect -708 25495 -706 25515
rect -612 25495 -610 25515
rect -588 25495 -586 25515
rect -540 25495 -538 25515
rect -492 25495 -490 25515
rect -444 25495 -442 25515
rect -396 25495 -394 25515
rect -300 25495 -298 25515
rect -276 25495 -274 25515
rect -228 25495 -226 25515
rect -12 25495 -10 25515
rect 156 25495 158 25515
rect 204 25495 206 25515
rect 252 25495 254 25515
rect 348 25495 350 25515
rect 468 25495 470 25515
rect 492 25495 494 25515
rect 564 25495 566 25515
rect 588 25495 590 25515
rect 636 25495 638 25515
rect 660 25495 662 25515
rect 732 25495 734 25515
rect 1092 25495 1094 25515
rect 1129 25495 1187 25496
rect 1308 25495 1310 25515
rect 1332 25495 1334 25515
rect 1380 25495 1382 25515
rect 1428 25495 1430 25515
rect 1476 25495 1478 25515
rect 1644 25495 1646 25515
rect 1692 25495 1694 25515
rect 1740 25495 1742 25515
rect 1788 25495 1790 25515
rect 2028 25495 2030 25515
rect 2076 25495 2078 25515
rect 2100 25495 2102 25515
rect 2124 25495 2126 25515
rect 2172 25495 2174 25515
rect 2220 25495 2222 25515
rect 2316 25495 2318 25515
rect 2412 25495 2414 25515
rect 2460 25495 2462 25515
rect 2508 25495 2510 25515
rect 2580 25495 2582 25515
rect 2604 25495 2606 25515
rect 2676 25495 2678 25515
rect 2700 25495 2702 25515
rect 2748 25495 2750 25515
rect 2772 25495 2774 25515
rect 2796 25495 2798 25515
rect 2844 25495 2846 25515
rect 2868 25495 2870 25515
rect 2892 25495 2894 25515
rect 2940 25495 2942 25515
rect 3012 25495 3014 25515
rect 3108 25495 3110 25515
rect 3252 25495 3254 25515
rect 3348 25495 3350 25515
rect 3396 25495 3398 25515
rect 3564 25495 3566 25515
rect 3636 25495 3638 25515
rect 3660 25495 3662 25515
rect 3732 25495 3734 25515
rect 3828 25495 3830 25515
rect 3924 25495 3926 25515
rect 4020 25495 4022 25515
rect 4044 25495 4046 25515
rect 4092 25495 4094 25515
rect 4140 25495 4142 25515
rect 4188 25495 4190 25515
rect 4191 25512 4205 25515
rect 4212 25512 4215 25515
rect 4236 25495 4238 25515
rect 4308 25495 4310 25515
rect 4332 25495 4334 25515
rect 4404 25495 4406 25515
rect 4500 25495 4502 25515
rect 4596 25495 4598 25515
rect 4692 25495 4694 25515
rect 4860 25495 4862 25515
rect 4956 25495 4958 25515
rect 4980 25495 4982 25515
rect 4993 25510 4996 25515
rect 5004 25510 5006 25515
rect 5003 25496 5006 25510
rect 5052 25495 5054 25515
rect 5100 25512 5102 25515
rect 5100 25495 5103 25512
rect 5124 25495 5126 25515
rect 5220 25495 5222 25515
rect 5268 25495 5270 25515
rect 5388 25495 5390 25515
rect 5484 25495 5486 25515
rect 5508 25495 5510 25515
rect 5532 25495 5534 25515
rect 5628 25495 5630 25515
rect 5652 25495 5654 25515
rect 5748 25495 5750 25515
rect 5796 25495 5798 25515
rect 5844 25495 5846 25515
rect 5892 25495 5894 25515
rect 6132 25495 6134 25515
rect 6180 25495 6182 25515
rect 6228 25495 6230 25515
rect 6252 25495 6254 25515
rect 6276 25495 6278 25515
rect 6324 25495 6326 25515
rect 6372 25495 6374 25515
rect 6492 25495 6494 25515
rect 6588 25495 6590 25515
rect 6612 25495 6614 25515
rect 6660 25495 6662 25515
rect 6684 25495 6686 25515
rect 6708 25495 6710 25515
rect 6780 25495 6782 25515
rect 6804 25495 6806 25515
rect 6900 25495 6902 25515
rect 6924 25495 6926 25515
rect 7020 25495 7022 25515
rect 7068 25495 7070 25515
rect 7164 25495 7166 25515
rect 7236 25495 7238 25515
rect 7332 25495 7334 25515
rect 7380 25495 7382 25515
rect 7428 25495 7430 25515
rect 7452 25495 7454 25515
rect 7476 25495 7478 25515
rect 7524 25495 7526 25515
rect 7548 25495 7550 25515
rect 7572 25495 7574 25515
rect 7620 25495 7622 25515
rect 7644 25495 7646 25515
rect 7668 25495 7670 25515
rect 7777 25510 7780 25515
rect 7788 25510 7790 25515
rect 7787 25496 7790 25510
rect 7884 25512 7886 25515
rect 7884 25495 7887 25512
rect 7956 25495 7958 25515
rect 7980 25496 7982 25515
rect 7969 25495 8003 25496
rect 8028 25495 8030 25515
rect 8113 25510 8116 25515
rect 8123 25496 8126 25510
rect 8196 25496 8198 25515
rect 8244 25512 8246 25515
rect 8124 25495 8126 25496
rect 8185 25495 8213 25496
rect 8244 25495 8247 25512
rect 8268 25495 8270 25515
rect 8292 25496 8294 25515
rect 8281 25495 8315 25496
rect 8340 25495 8342 25515
rect 8364 25495 8366 25515
rect 8388 25495 8390 25515
rect 8436 25495 8438 25515
rect 8652 25495 8654 25515
rect 8700 25495 8702 25515
rect 8748 25495 8750 25515
rect 8820 25495 8822 25515
rect 8844 25495 8846 25515
rect 8868 25495 8870 25515
rect 9516 25495 9518 25515
rect 9660 25495 9662 25515
rect 9684 25495 9686 25515
rect 9687 25512 9701 25515
rect 9708 25512 9711 25515
rect 9756 25495 9758 25515
rect 9780 25495 9782 25515
rect 9804 25495 9806 25515
rect 9852 25495 9854 25515
rect 9900 25495 9902 25515
rect 9948 25495 9950 25515
rect 9996 25496 9998 25515
rect 9985 25495 10019 25496
rect 10068 25495 10070 25515
rect 10092 25495 10094 25515
rect 10116 25495 10118 25515
rect 10164 25495 10166 25515
rect 10188 25495 10190 25515
rect 10212 25495 10214 25515
rect 10284 25495 10286 25515
rect 10308 25496 10310 25515
rect 10297 25495 10331 25496
rect 10332 25495 10334 25515
rect 10380 25495 10382 25515
rect 10404 25495 10406 25515
rect 10428 25495 10430 25515
rect 10476 25495 10478 25515
rect 10500 25495 10502 25515
rect 10524 25495 10526 25515
rect 10572 25495 10574 25515
rect 10596 25495 10598 25515
rect 10620 25495 10622 25515
rect 10668 25496 10670 25515
rect 10633 25495 10691 25496
rect 10692 25495 10694 25515
rect 10716 25495 10718 25515
rect 10788 25495 10790 25515
rect 10956 25495 10958 25515
rect 11004 25495 11006 25515
rect 11052 25495 11054 25515
rect 11100 25495 11102 25515
rect 11172 25495 11174 25515
rect 11220 25495 11222 25515
rect 11340 25495 11342 25515
rect 11436 25495 11438 25515
rect 11532 25495 11534 25515
rect 11580 25495 11582 25515
rect 11628 25495 11630 25515
rect 11676 25495 11678 25515
rect 11724 25495 11726 25515
rect 11772 25495 11774 25515
rect 11796 25495 11798 25515
rect 11892 25495 11894 25515
rect 11988 25495 11990 25515
rect 12060 25495 12062 25515
rect 12132 25495 12134 25515
rect 12228 25495 12230 25515
rect 12276 25495 12278 25515
rect 12324 25495 12326 25515
rect 12420 25495 12422 25515
rect 12444 25495 12446 25515
rect 12492 25495 12494 25515
rect 12516 25495 12518 25515
rect 12540 25495 12542 25515
rect 12588 25495 12590 25515
rect 12636 25495 12638 25515
rect 12732 25495 12734 25515
rect 12756 25495 12758 25515
rect 12804 25495 12806 25515
rect 12828 25495 12830 25515
rect 12852 25495 12854 25515
rect 12948 25495 12950 25515
rect 12972 25495 12974 25515
rect 13044 25495 13046 25515
rect 13068 25495 13070 25515
rect 13116 25495 13118 25515
rect 13284 25495 13286 25515
rect 13332 25495 13334 25515
rect 13572 25495 13574 25515
rect 13620 25495 13622 25515
rect 13668 25495 13670 25515
rect 13716 25495 13718 25515
rect 13764 25495 13766 25515
rect 13860 25495 13862 25515
rect 13956 25495 13958 25515
rect 14004 25495 14006 25515
rect 14100 25495 14102 25515
rect 15180 25495 15182 25515
rect 15276 25495 15278 25515
rect 15420 25495 15422 25515
rect 15492 25495 15494 25515
rect 15660 25495 15662 25515
rect 15708 25495 15710 25515
rect 15732 25495 15734 25515
rect 15756 25495 15758 25515
rect 15804 25495 15806 25515
rect 15828 25495 15830 25515
rect 15852 25495 15854 25515
rect 15900 25495 15902 25515
rect 15948 25495 15950 25515
rect 16044 25495 16046 25515
rect 16068 25495 16070 25515
rect 16164 25495 16166 25515
rect 16260 25495 16262 25515
rect 16308 25495 16310 25515
rect 16332 25495 16334 25515
rect 16356 25495 16358 25515
rect 16404 25495 16406 25515
rect 16452 25495 16454 25515
rect 16548 25495 16550 25515
rect 16572 25495 16574 25515
rect 16620 25495 16622 25515
rect 16668 25495 16670 25515
rect 16716 25495 16718 25515
rect 16764 25495 16766 25515
rect 16812 25495 16814 25515
rect 16884 25495 16886 25515
rect 16908 25495 16910 25515
rect 16980 25495 16982 25515
rect 17052 25495 17054 25515
rect 17196 25495 17198 25515
rect 17220 25495 17222 25515
rect 17292 25495 17294 25515
rect 17316 25495 17318 25515
rect 18084 25495 18086 25515
rect 18132 25495 18134 25515
rect 18228 25495 18230 25515
rect 18396 25495 18398 25515
rect 18492 25495 18494 25515
rect 18516 25495 18518 25515
rect 18564 25495 18566 25515
rect 18612 25495 18614 25515
rect 18660 25495 18662 25515
rect 18756 25495 18758 25515
rect 18852 25495 18854 25515
rect 18900 25495 18902 25515
rect 18996 25495 18998 25515
rect 19020 25495 19022 25515
rect 19092 25495 19094 25515
rect 19116 25495 19118 25515
rect 19140 25495 19142 25515
rect 19188 25495 19190 25515
rect 19236 25495 19238 25515
rect 19332 25495 19334 25515
rect 19476 25495 19478 25515
rect 19788 25495 19790 25515
rect 19836 25495 19838 25515
rect 19860 25495 19862 25515
rect 19884 25495 19886 25515
rect 19932 25495 19934 25515
rect 19956 25495 19958 25515
rect 19980 25495 19982 25515
rect 20028 25495 20030 25515
rect 20052 25495 20054 25515
rect 20076 25495 20078 25515
rect 20148 25495 20150 25515
rect 20172 25495 20174 25515
rect 20196 25495 20198 25515
rect 20268 25495 20270 25515
rect 20292 25495 20294 25515
rect 20388 25495 20390 25515
rect 20412 25495 20414 25515
rect 20508 25495 20510 25515
rect 20556 25495 20558 25515
rect 20604 25495 20606 25515
rect 20916 25495 20918 25515
rect 20964 25495 20966 25515
rect 21012 25495 21014 25515
rect 21060 25495 21062 25515
rect 21108 25495 21110 25515
rect 21204 25495 21206 25515
rect 21300 25495 21302 25515
rect 21324 25495 21326 25515
rect 21444 25495 21446 25515
rect 21468 25495 21470 25515
rect 21564 25495 21566 25515
rect 21588 25495 21590 25515
rect 21684 25495 21686 25515
rect 21708 25495 21710 25515
rect 21828 25495 21830 25515
rect 21924 25495 21926 25515
rect 22068 25495 22070 25515
rect 22188 25495 22190 25515
rect 22212 25495 22214 25515
rect 22884 25495 22886 25515
rect 22980 25495 22982 25515
rect 23076 25495 23078 25515
rect 23100 25495 23102 25515
rect 23124 25495 23126 25515
rect 23244 25495 23246 25515
rect 23340 25495 23342 25515
rect 23412 25495 23414 25515
rect 23460 25495 23462 25515
rect 23508 25495 23510 25515
rect 23556 25495 23558 25515
rect 23604 25495 23606 25515
rect 23652 25495 23654 25515
rect 23676 25495 23678 25515
rect 23772 25495 23774 25515
rect 23820 25495 23822 25515
rect 23916 25495 23918 25515
rect 24012 25495 24014 25515
rect 24060 25495 24062 25515
rect 24156 25495 24158 25515
rect 24492 25495 24494 25515
rect 24516 25495 24518 25515
rect 24588 25495 24590 25515
rect 24612 25495 24614 25515
rect 24684 25495 24686 25515
rect 24732 25495 24734 25515
rect 24756 25495 24758 25515
rect 24780 25495 24782 25515
rect 24852 25495 24854 25515
rect 24876 25495 24878 25515
rect 24972 25495 24974 25515
rect 25068 25495 25070 25515
rect 25164 25495 25166 25515
rect 25260 25495 25262 25515
rect 25284 25495 25286 25515
rect 25356 25495 25358 25515
rect 25380 25495 25382 25515
rect 25404 25495 25406 25515
rect 25500 25495 25502 25515
rect 25596 25495 25598 25515
rect 25609 25495 25643 25496
rect -15215 25491 -14371 25495
rect -15108 25488 -15106 25491
rect -15108 25472 -15105 25488
rect -15119 25471 -15085 25472
rect -14892 25471 -14890 25491
rect -14676 25471 -14674 25491
rect -14460 25471 -14458 25491
rect -14409 25488 -14395 25491
rect -14385 25488 -14371 25491
rect -14361 25491 -12427 25495
rect -14361 25488 -14347 25491
rect -14340 25488 -14337 25491
rect -14111 25471 -14053 25472
rect -13788 25471 -13786 25491
rect -13428 25471 -13426 25491
rect -12756 25471 -12754 25491
rect -12660 25471 -12658 25491
rect -12441 25488 -12427 25491
rect -12417 25491 8213 25495
rect -12417 25488 -12403 25491
rect -12396 25488 -12393 25491
rect -12348 25471 -12346 25491
rect -12252 25471 -12250 25491
rect -12156 25471 -12154 25491
rect -12060 25471 -12058 25491
rect -11844 25471 -11842 25491
rect -11676 25471 -11674 25491
rect -11508 25471 -11506 25491
rect -11436 25471 -11434 25491
rect -11412 25471 -11410 25491
rect -11340 25471 -11338 25491
rect -11231 25471 -11197 25472
rect -11196 25471 -11194 25491
rect -11100 25471 -11098 25491
rect -10740 25488 -10738 25491
rect -10764 25471 -10761 25488
rect -10740 25471 -10737 25488
rect -10644 25471 -10642 25491
rect -9996 25471 -9994 25491
rect -9900 25471 -9898 25491
rect -9732 25471 -9730 25491
rect -9516 25471 -9514 25491
rect -9468 25488 -9466 25491
rect -9468 25471 -9465 25488
rect -9348 25471 -9346 25491
rect -9180 25471 -9178 25491
rect -8604 25488 -8602 25491
rect -8604 25471 -8601 25488
rect -8436 25471 -8434 25491
rect -8364 25471 -8362 25491
rect -8340 25471 -8338 25491
rect -8268 25471 -8266 25491
rect -8231 25471 -8173 25472
rect -8100 25471 -8098 25491
rect -8004 25471 -8002 25491
rect -7977 25488 -7963 25491
rect -7932 25471 -7930 25491
rect -7620 25471 -7618 25491
rect -7617 25488 -7603 25491
rect -7524 25471 -7522 25491
rect -7356 25471 -7354 25491
rect -7308 25471 -7306 25491
rect -7212 25471 -7210 25491
rect -7044 25471 -7042 25491
rect -6993 25488 -6979 25491
rect -6948 25471 -6946 25491
rect -6852 25471 -6850 25491
rect -6780 25471 -6778 25491
rect -6756 25471 -6754 25491
rect -6660 25471 -6658 25491
rect -6612 25471 -6610 25491
rect -6516 25471 -6514 25491
rect -6513 25488 -6499 25491
rect -6372 25471 -6370 25491
rect -6156 25471 -6154 25491
rect -6060 25471 -6058 25491
rect -6036 25471 -6034 25491
rect -5892 25471 -5890 25491
rect -5268 25472 -5266 25491
rect -5279 25471 -5245 25472
rect -5196 25471 -5194 25491
rect -5172 25471 -5170 25491
rect -5100 25471 -5098 25491
rect -5076 25472 -5074 25491
rect -5087 25471 -5053 25472
rect -4980 25471 -4978 25491
rect -4956 25472 -4954 25491
rect -4860 25472 -4858 25491
rect -4644 25472 -4642 25491
rect -4967 25471 -4933 25472
rect -4871 25471 -4837 25472
rect -4655 25471 -4621 25472
rect -4535 25471 -4501 25472
rect -4500 25471 -4498 25491
rect -4404 25471 -4402 25491
rect -4391 25471 -4333 25472
rect -4308 25471 -4306 25491
rect -4260 25471 -4258 25491
rect -4164 25471 -4162 25491
rect -4020 25471 -4018 25491
rect -3876 25471 -3874 25491
rect -3732 25471 -3730 25491
rect -3564 25471 -3562 25491
rect -3516 25471 -3514 25491
rect -3468 25471 -3466 25491
rect -3420 25471 -3418 25491
rect -3324 25471 -3322 25491
rect -3228 25471 -3226 25491
rect -3132 25471 -3130 25491
rect -3012 25471 -3010 25491
rect -2964 25471 -2962 25491
rect -2916 25471 -2914 25491
rect -2892 25471 -2890 25491
rect -2868 25471 -2866 25491
rect -2820 25471 -2818 25491
rect -2796 25471 -2794 25491
rect -2772 25471 -2770 25491
rect -2676 25471 -2674 25491
rect -2580 25471 -2578 25491
rect -2364 25471 -2362 25491
rect -2316 25471 -2314 25491
rect -2268 25471 -2266 25491
rect -2244 25471 -2242 25491
rect -2172 25471 -2170 25491
rect -2148 25471 -2146 25491
rect -2076 25471 -2074 25491
rect -2052 25471 -2050 25491
rect -1980 25471 -1978 25491
rect -1884 25471 -1882 25491
rect -1572 25471 -1570 25491
rect -1476 25471 -1474 25491
rect -1380 25471 -1378 25491
rect -1356 25471 -1354 25491
rect -1308 25471 -1306 25491
rect -1260 25471 -1258 25491
rect -1140 25471 -1138 25491
rect -708 25471 -706 25491
rect -612 25471 -610 25491
rect -588 25471 -586 25491
rect -540 25471 -538 25491
rect -492 25471 -490 25491
rect -444 25471 -442 25491
rect -396 25471 -394 25491
rect -300 25471 -298 25491
rect -276 25471 -274 25491
rect -228 25471 -226 25491
rect -12 25471 -10 25491
rect 156 25471 158 25491
rect 204 25471 206 25491
rect 252 25471 254 25491
rect 348 25471 350 25491
rect 468 25471 470 25491
rect 492 25471 494 25491
rect 564 25471 566 25491
rect 588 25471 590 25491
rect 636 25471 638 25491
rect 660 25471 662 25491
rect 732 25471 734 25491
rect 1092 25471 1094 25491
rect 1129 25486 1132 25491
rect 1139 25472 1142 25486
rect 1140 25471 1142 25472
rect 1236 25471 1239 25488
rect 1308 25471 1310 25491
rect 1332 25471 1334 25491
rect 1380 25471 1382 25491
rect 1428 25471 1430 25491
rect 1476 25471 1478 25491
rect 1644 25471 1646 25491
rect 1692 25471 1694 25491
rect 1740 25471 1742 25491
rect 1788 25471 1790 25491
rect 2028 25471 2030 25491
rect 2076 25471 2078 25491
rect 2100 25471 2102 25491
rect 2124 25471 2126 25491
rect 2172 25471 2174 25491
rect 2220 25471 2222 25491
rect 2316 25471 2318 25491
rect 2412 25471 2414 25491
rect 2460 25471 2462 25491
rect 2508 25471 2510 25491
rect 2580 25471 2582 25491
rect 2604 25471 2606 25491
rect 2676 25471 2678 25491
rect 2700 25471 2702 25491
rect 2748 25471 2750 25491
rect 2772 25471 2774 25491
rect 2796 25471 2798 25491
rect 2844 25471 2846 25491
rect 2868 25471 2870 25491
rect 2892 25471 2894 25491
rect 2940 25471 2942 25491
rect 3012 25471 3014 25491
rect 3108 25471 3110 25491
rect 3252 25471 3254 25491
rect 3348 25471 3350 25491
rect 3396 25471 3398 25491
rect 3564 25471 3566 25491
rect 3636 25471 3638 25491
rect 3660 25471 3662 25491
rect 3732 25471 3734 25491
rect 3828 25471 3830 25491
rect 3924 25471 3926 25491
rect 4020 25471 4022 25491
rect 4044 25471 4046 25491
rect 4092 25471 4094 25491
rect 4140 25471 4142 25491
rect 4188 25471 4190 25491
rect 4236 25471 4238 25491
rect 4308 25471 4310 25491
rect 4332 25471 4334 25491
rect 4404 25471 4406 25491
rect 4500 25471 4502 25491
rect 4596 25471 4598 25491
rect 4692 25471 4694 25491
rect 4860 25471 4862 25491
rect 4956 25471 4958 25491
rect 4980 25471 4982 25491
rect 5052 25471 5054 25491
rect 5079 25488 5093 25491
rect 5100 25488 5103 25491
rect 5124 25471 5126 25491
rect 5220 25471 5222 25491
rect 5268 25471 5270 25491
rect 5388 25471 5390 25491
rect 5484 25471 5486 25491
rect 5508 25471 5510 25491
rect 5532 25471 5534 25491
rect 5628 25471 5630 25491
rect 5652 25471 5654 25491
rect 5748 25471 5750 25491
rect 5796 25471 5798 25491
rect 5844 25471 5846 25491
rect 5892 25471 5894 25491
rect 6132 25471 6134 25491
rect 6180 25471 6182 25491
rect 6228 25471 6230 25491
rect 6252 25471 6254 25491
rect 6276 25471 6278 25491
rect 6324 25471 6326 25491
rect 6372 25471 6374 25491
rect 6492 25471 6494 25491
rect 6588 25471 6590 25491
rect 6612 25471 6614 25491
rect 6660 25471 6662 25491
rect 6684 25471 6686 25491
rect 6708 25471 6710 25491
rect 6780 25471 6782 25491
rect 6804 25471 6806 25491
rect 6900 25471 6902 25491
rect 6924 25471 6926 25491
rect 7020 25471 7022 25491
rect 7068 25471 7070 25491
rect 7164 25471 7166 25491
rect 7236 25471 7238 25491
rect 7332 25471 7334 25491
rect 7380 25471 7382 25491
rect 7428 25471 7430 25491
rect 7452 25471 7454 25491
rect 7476 25471 7478 25491
rect 7524 25471 7526 25491
rect 7548 25471 7550 25491
rect 7572 25471 7574 25491
rect 7620 25471 7622 25491
rect 7644 25471 7646 25491
rect 7668 25471 7670 25491
rect 7863 25488 7877 25491
rect 7884 25488 7887 25491
rect 7956 25471 7958 25491
rect 7969 25486 7972 25491
rect 7980 25486 7982 25491
rect 7979 25472 7982 25486
rect 8028 25471 8030 25491
rect 8124 25471 8126 25491
rect 8185 25486 8188 25491
rect 8196 25486 8198 25491
rect 8199 25488 8213 25491
rect 8223 25491 25643 25495
rect 8223 25488 8237 25491
rect 8244 25488 8247 25491
rect 8195 25472 8198 25486
rect 8268 25471 8270 25491
rect 8281 25486 8284 25491
rect 8292 25488 8294 25491
rect 8292 25486 8295 25488
rect 8291 25472 8295 25486
rect 8340 25471 8342 25491
rect 8364 25471 8366 25491
rect 8388 25488 8390 25491
rect 8388 25471 8391 25488
rect 8436 25471 8438 25491
rect 8652 25471 8654 25491
rect 8700 25471 8702 25491
rect 8748 25471 8750 25491
rect 8820 25471 8822 25491
rect 8844 25471 8846 25491
rect 8868 25471 8870 25491
rect 9516 25471 9518 25491
rect 9660 25471 9662 25491
rect 9684 25471 9686 25491
rect 9756 25471 9758 25491
rect 9780 25471 9782 25491
rect 9804 25471 9806 25491
rect 9852 25471 9854 25491
rect 9900 25471 9902 25491
rect 9948 25471 9950 25491
rect 9985 25486 9988 25491
rect 9996 25486 9998 25491
rect 9995 25472 9998 25486
rect 10068 25471 10070 25491
rect 10092 25488 10094 25491
rect 10092 25471 10095 25488
rect 10116 25471 10118 25491
rect 10164 25471 10166 25491
rect 10188 25471 10190 25491
rect 10212 25471 10214 25491
rect 10284 25471 10286 25491
rect 10297 25486 10300 25491
rect 10308 25486 10310 25491
rect 10307 25472 10310 25486
rect 10332 25471 10334 25491
rect 10380 25471 10382 25491
rect 10404 25488 10406 25491
rect 10404 25471 10407 25488
rect 10428 25471 10430 25491
rect 10476 25471 10478 25491
rect 10500 25471 10502 25491
rect 10524 25471 10526 25491
rect 10572 25471 10574 25491
rect 10596 25471 10598 25491
rect 10620 25471 10622 25491
rect 10657 25486 10660 25491
rect 10668 25486 10670 25491
rect 10667 25472 10670 25486
rect 10692 25471 10694 25491
rect 10716 25471 10718 25491
rect 10788 25471 10790 25491
rect 10956 25471 10958 25491
rect 11004 25471 11006 25491
rect 11052 25471 11054 25491
rect 11100 25471 11102 25491
rect 11172 25471 11174 25491
rect 11220 25471 11222 25491
rect 11340 25471 11342 25491
rect 11436 25471 11438 25491
rect 11532 25471 11534 25491
rect 11580 25471 11582 25491
rect 11628 25471 11630 25491
rect 11676 25471 11678 25491
rect 11724 25471 11726 25491
rect 11772 25471 11774 25491
rect 11796 25471 11798 25491
rect 11892 25471 11894 25491
rect 11988 25471 11990 25491
rect 12060 25471 12062 25491
rect 12132 25471 12134 25491
rect 12228 25471 12230 25491
rect 12276 25471 12278 25491
rect 12324 25471 12326 25491
rect 12420 25471 12422 25491
rect 12444 25471 12446 25491
rect 12492 25471 12494 25491
rect 12516 25471 12518 25491
rect 12540 25471 12542 25491
rect 12588 25471 12590 25491
rect 12636 25471 12638 25491
rect 12732 25471 12734 25491
rect 12756 25471 12758 25491
rect 12804 25471 12806 25491
rect 12828 25471 12830 25491
rect 12852 25471 12854 25491
rect 12948 25471 12950 25491
rect 12972 25471 12974 25491
rect 13044 25471 13046 25491
rect 13068 25471 13070 25491
rect 13116 25471 13118 25491
rect 13284 25471 13286 25491
rect 13332 25471 13334 25491
rect 13572 25471 13574 25491
rect 13620 25471 13622 25491
rect 13668 25471 13670 25491
rect 13716 25471 13718 25491
rect 13764 25471 13766 25491
rect 13860 25471 13862 25491
rect 13956 25471 13958 25491
rect 14004 25471 14006 25491
rect 14100 25471 14102 25491
rect 15180 25471 15182 25491
rect 15276 25471 15278 25491
rect 15420 25471 15422 25491
rect 15492 25471 15494 25491
rect 15660 25471 15662 25491
rect 15708 25471 15710 25491
rect 15732 25471 15734 25491
rect 15756 25471 15758 25491
rect 15804 25471 15806 25491
rect 15828 25471 15830 25491
rect 15852 25471 15854 25491
rect 15900 25471 15902 25491
rect 15948 25471 15950 25491
rect 16044 25471 16046 25491
rect 16068 25471 16070 25491
rect 16164 25471 16166 25491
rect 16260 25471 16262 25491
rect 16308 25471 16310 25491
rect 16332 25471 16334 25491
rect 16356 25471 16358 25491
rect 16404 25471 16406 25491
rect 16452 25471 16454 25491
rect 16548 25471 16550 25491
rect 16572 25471 16574 25491
rect 16620 25471 16622 25491
rect 16668 25471 16670 25491
rect 16716 25471 16718 25491
rect 16764 25471 16766 25491
rect 16812 25471 16814 25491
rect 16884 25471 16886 25491
rect 16908 25471 16910 25491
rect 16980 25471 16982 25491
rect 17052 25471 17054 25491
rect 17196 25471 17198 25491
rect 17220 25471 17222 25491
rect 17292 25471 17294 25491
rect 17316 25471 17318 25491
rect 18084 25471 18086 25491
rect 18132 25471 18134 25491
rect 18228 25471 18230 25491
rect 18396 25471 18398 25491
rect 18492 25471 18494 25491
rect 18516 25471 18518 25491
rect 18564 25471 18566 25491
rect 18612 25471 18614 25491
rect 18660 25471 18662 25491
rect 18756 25471 18758 25491
rect 18852 25472 18854 25491
rect 18817 25471 18875 25472
rect 18900 25471 18902 25491
rect 18996 25471 18998 25491
rect 19020 25471 19022 25491
rect 19092 25471 19094 25491
rect 19116 25471 19118 25491
rect 19140 25471 19142 25491
rect 19188 25471 19190 25491
rect 19236 25471 19238 25491
rect 19332 25471 19334 25491
rect 19476 25471 19478 25491
rect 19788 25471 19790 25491
rect 19836 25471 19838 25491
rect 19860 25471 19862 25491
rect 19884 25471 19886 25491
rect 19932 25471 19934 25491
rect 19956 25471 19958 25491
rect 19980 25471 19982 25491
rect 20028 25471 20030 25491
rect 20052 25471 20054 25491
rect 20076 25471 20078 25491
rect 20148 25471 20150 25491
rect 20172 25471 20174 25491
rect 20196 25471 20198 25491
rect 20268 25471 20270 25491
rect 20292 25471 20294 25491
rect 20388 25471 20390 25491
rect 20412 25471 20414 25491
rect 20508 25471 20510 25491
rect 20556 25471 20558 25491
rect 20604 25471 20606 25491
rect 20785 25471 20843 25472
rect 20916 25471 20918 25491
rect 20964 25471 20966 25491
rect 21012 25471 21014 25491
rect 21060 25471 21062 25491
rect 21108 25471 21110 25491
rect 21204 25471 21206 25491
rect 21300 25471 21302 25491
rect 21324 25471 21326 25491
rect 21444 25471 21446 25491
rect 21468 25471 21470 25491
rect 21564 25471 21566 25491
rect 21588 25471 21590 25491
rect 21684 25471 21686 25491
rect 21708 25471 21710 25491
rect 21828 25471 21830 25491
rect 21924 25471 21926 25491
rect 22068 25471 22070 25491
rect 22188 25471 22190 25491
rect 22212 25471 22214 25491
rect 22884 25471 22886 25491
rect 22980 25471 22982 25491
rect 23076 25471 23078 25491
rect 23100 25471 23102 25491
rect 23124 25471 23126 25491
rect 23244 25471 23246 25491
rect 23340 25471 23342 25491
rect 23412 25471 23414 25491
rect 23460 25471 23462 25491
rect 23508 25471 23510 25491
rect 23556 25471 23558 25491
rect 23604 25471 23606 25491
rect 23652 25471 23654 25491
rect 23676 25471 23678 25491
rect 23772 25471 23774 25491
rect 23820 25471 23822 25491
rect 23916 25471 23918 25491
rect 24012 25471 24014 25491
rect 24060 25471 24062 25491
rect 24156 25471 24158 25491
rect 24492 25471 24494 25491
rect 24516 25471 24518 25491
rect 24588 25471 24590 25491
rect 24612 25471 24614 25491
rect 24684 25471 24686 25491
rect 24732 25471 24734 25491
rect 24756 25471 24758 25491
rect 24780 25471 24782 25491
rect 24852 25471 24854 25491
rect 24876 25471 24878 25491
rect 24972 25471 24974 25491
rect 25068 25471 25070 25491
rect 25164 25471 25166 25491
rect 25260 25471 25262 25491
rect 25284 25471 25286 25491
rect 25356 25471 25358 25491
rect 25380 25471 25382 25491
rect 25404 25471 25406 25491
rect 25500 25471 25502 25491
rect 25596 25472 25598 25491
rect 25585 25471 25619 25472
rect -15119 25467 -10771 25471
rect -15119 25464 -15115 25467
rect -15108 25464 -15105 25467
rect -14999 25447 -14965 25448
rect -14892 25447 -14890 25467
rect -14676 25447 -14674 25467
rect -14460 25447 -14458 25467
rect -14111 25462 -14108 25467
rect -14101 25448 -14098 25462
rect -14100 25447 -14098 25448
rect -14004 25447 -14001 25464
rect -13788 25447 -13786 25467
rect -13428 25447 -13426 25467
rect -13377 25464 -13363 25467
rect -12756 25447 -12754 25467
rect -12660 25447 -12658 25467
rect -12348 25447 -12346 25467
rect -12252 25447 -12250 25467
rect -12156 25447 -12154 25467
rect -12060 25447 -12058 25467
rect -11844 25448 -11842 25467
rect -11879 25447 -11821 25448
rect -11676 25447 -11674 25467
rect -11508 25447 -11506 25467
rect -11436 25447 -11434 25467
rect -11412 25447 -11410 25467
rect -11340 25447 -11338 25467
rect -11196 25447 -11194 25467
rect -11100 25447 -11098 25467
rect -10785 25464 -10771 25467
rect -10764 25467 -8635 25471
rect -10764 25464 -10747 25467
rect -10740 25464 -10737 25467
rect -10764 25447 -10762 25464
rect -10644 25447 -10642 25467
rect -9996 25447 -9994 25467
rect -9900 25447 -9898 25467
rect -9732 25447 -9730 25467
rect -9516 25447 -9514 25467
rect -9489 25464 -9475 25467
rect -9468 25464 -9465 25467
rect -9348 25447 -9346 25467
rect -9180 25447 -9178 25467
rect -8649 25464 -8635 25467
rect -8625 25467 1229 25471
rect -8625 25464 -8611 25467
rect -8604 25464 -8601 25467
rect -8663 25447 -8629 25448
rect -8436 25447 -8434 25467
rect -8364 25447 -8362 25467
rect -8340 25447 -8338 25467
rect -8268 25447 -8266 25467
rect -8100 25464 -8098 25467
rect -8100 25447 -8097 25464
rect -8004 25447 -8002 25467
rect -7932 25447 -7930 25467
rect -7620 25447 -7618 25467
rect -7524 25447 -7522 25467
rect -7356 25447 -7354 25467
rect -7308 25447 -7306 25467
rect -7212 25447 -7210 25467
rect -7044 25447 -7042 25467
rect -6948 25447 -6946 25467
rect -6852 25447 -6850 25467
rect -6780 25447 -6778 25467
rect -6756 25447 -6754 25467
rect -6660 25447 -6658 25467
rect -6612 25447 -6610 25467
rect -6516 25447 -6514 25467
rect -6372 25447 -6370 25467
rect -6156 25448 -6154 25467
rect -6167 25447 -6133 25448
rect -6060 25447 -6058 25467
rect -6036 25447 -6034 25467
rect -5892 25447 -5890 25467
rect -5279 25462 -5276 25467
rect -5268 25462 -5266 25467
rect -5269 25448 -5266 25462
rect -5196 25447 -5194 25467
rect -5172 25464 -5170 25467
rect -5172 25447 -5169 25464
rect -5100 25447 -5098 25467
rect -5087 25462 -5084 25467
rect -5076 25462 -5074 25467
rect -5077 25448 -5074 25462
rect -4980 25464 -4978 25467
rect -4980 25447 -4977 25464
rect -4967 25462 -4964 25467
rect -4956 25462 -4954 25467
rect -4871 25462 -4868 25467
rect -4860 25464 -4858 25467
rect -4860 25462 -4857 25464
rect -4655 25462 -4652 25467
rect -4644 25462 -4642 25467
rect -4957 25448 -4954 25462
rect -4861 25448 -4857 25462
rect -4645 25448 -4642 25462
rect -4500 25447 -4498 25467
rect -4404 25447 -4402 25467
rect -4308 25447 -4306 25467
rect -4260 25464 -4258 25467
rect -4260 25447 -4257 25464
rect -4164 25447 -4162 25467
rect -4020 25447 -4018 25467
rect -3876 25447 -3874 25467
rect -3732 25447 -3730 25467
rect -3564 25447 -3562 25467
rect -3516 25447 -3514 25467
rect -3468 25447 -3466 25467
rect -3420 25447 -3418 25467
rect -3324 25447 -3322 25467
rect -3228 25447 -3226 25467
rect -3215 25447 -3157 25448
rect -3132 25447 -3130 25467
rect -3012 25447 -3010 25467
rect -2964 25447 -2962 25467
rect -2916 25447 -2914 25467
rect -2892 25447 -2890 25467
rect -2868 25447 -2866 25467
rect -2820 25447 -2818 25467
rect -2796 25447 -2794 25467
rect -2772 25447 -2770 25467
rect -2676 25447 -2674 25467
rect -2580 25447 -2578 25467
rect -2364 25447 -2362 25467
rect -2316 25447 -2314 25467
rect -2268 25447 -2266 25467
rect -2244 25447 -2242 25467
rect -2172 25447 -2170 25467
rect -2148 25447 -2146 25467
rect -2076 25447 -2074 25467
rect -2052 25447 -2050 25467
rect -1980 25447 -1978 25467
rect -1943 25447 -1909 25448
rect -1884 25447 -1882 25467
rect -1572 25447 -1570 25467
rect -1476 25447 -1474 25467
rect -1380 25447 -1378 25467
rect -1356 25447 -1354 25467
rect -1308 25447 -1306 25467
rect -1260 25447 -1258 25467
rect -1140 25447 -1138 25467
rect -708 25447 -706 25467
rect -612 25447 -610 25467
rect -588 25447 -586 25467
rect -540 25447 -538 25467
rect -492 25447 -490 25467
rect -444 25447 -442 25467
rect -396 25447 -394 25467
rect -359 25447 -301 25448
rect -300 25447 -298 25467
rect -276 25447 -274 25467
rect -228 25447 -226 25467
rect -12 25447 -10 25467
rect 156 25447 158 25467
rect 204 25447 206 25467
rect 252 25447 254 25467
rect 348 25447 350 25467
rect 468 25447 470 25467
rect 492 25447 494 25467
rect 564 25447 566 25467
rect 588 25447 590 25467
rect 636 25447 638 25467
rect 660 25447 662 25467
rect 732 25447 734 25467
rect 1092 25447 1094 25467
rect 1140 25447 1142 25467
rect 1215 25464 1229 25467
rect 1236 25467 10733 25471
rect 1236 25464 1253 25467
rect 1236 25447 1238 25464
rect 1308 25447 1310 25467
rect 1332 25447 1334 25467
rect 1380 25447 1382 25467
rect 1428 25447 1430 25467
rect 1476 25447 1478 25467
rect 1644 25447 1646 25467
rect 1692 25447 1694 25467
rect 1740 25447 1742 25467
rect 1788 25447 1790 25467
rect 2028 25447 2030 25467
rect 2076 25447 2078 25467
rect 2100 25447 2102 25467
rect 2124 25447 2126 25467
rect 2172 25447 2174 25467
rect 2220 25447 2222 25467
rect 2316 25447 2318 25467
rect 2412 25447 2414 25467
rect 2460 25447 2462 25467
rect 2508 25447 2510 25467
rect 2580 25447 2582 25467
rect 2604 25447 2606 25467
rect 2676 25447 2678 25467
rect 2700 25447 2702 25467
rect 2748 25447 2750 25467
rect 2772 25447 2774 25467
rect 2796 25447 2798 25467
rect 2844 25447 2846 25467
rect 2868 25447 2870 25467
rect 2892 25447 2894 25467
rect 2940 25447 2942 25467
rect 3012 25447 3014 25467
rect 3108 25447 3110 25467
rect 3252 25447 3254 25467
rect 3348 25447 3350 25467
rect 3396 25447 3398 25467
rect 3564 25447 3566 25467
rect 3636 25447 3638 25467
rect 3660 25447 3662 25467
rect 3673 25447 3731 25448
rect 3732 25447 3734 25467
rect 3828 25447 3830 25467
rect 3924 25447 3926 25467
rect 4020 25447 4022 25467
rect 4044 25447 4046 25467
rect 4092 25447 4094 25467
rect 4140 25447 4142 25467
rect 4188 25447 4190 25467
rect 4236 25447 4238 25467
rect 4308 25447 4310 25467
rect 4332 25447 4334 25467
rect 4404 25447 4406 25467
rect 4500 25447 4502 25467
rect 4596 25447 4598 25467
rect 4692 25447 4694 25467
rect 4860 25447 4862 25467
rect 4956 25447 4958 25467
rect 4980 25447 4982 25467
rect 5052 25447 5054 25467
rect 5124 25447 5126 25467
rect 5220 25447 5222 25467
rect 5268 25447 5270 25467
rect 5388 25447 5390 25467
rect 5484 25447 5486 25467
rect 5508 25447 5510 25467
rect 5532 25447 5534 25467
rect 5628 25447 5630 25467
rect 5652 25447 5654 25467
rect 5748 25447 5750 25467
rect 5796 25447 5798 25467
rect 5844 25447 5846 25467
rect 5892 25447 5894 25467
rect 6132 25447 6134 25467
rect 6180 25447 6182 25467
rect 6228 25447 6230 25467
rect 6252 25447 6254 25467
rect 6276 25447 6278 25467
rect 6324 25447 6326 25467
rect 6372 25447 6374 25467
rect 6492 25447 6494 25467
rect 6588 25447 6590 25467
rect 6612 25447 6614 25467
rect 6660 25447 6662 25467
rect 6684 25447 6686 25467
rect 6708 25447 6710 25467
rect 6780 25447 6782 25467
rect 6804 25447 6806 25467
rect 6900 25447 6902 25467
rect 6924 25447 6926 25467
rect 7020 25447 7022 25467
rect 7068 25447 7070 25467
rect 7164 25447 7166 25467
rect 7236 25447 7238 25467
rect 7332 25447 7334 25467
rect 7380 25447 7382 25467
rect 7428 25447 7430 25467
rect 7452 25447 7454 25467
rect 7476 25447 7478 25467
rect 7524 25447 7526 25467
rect 7548 25447 7550 25467
rect 7572 25447 7574 25467
rect 7620 25447 7622 25467
rect 7644 25447 7646 25467
rect 7668 25447 7670 25467
rect 7956 25447 7958 25467
rect 8028 25447 8030 25467
rect 8055 25464 8069 25467
rect 8124 25447 8126 25467
rect 8268 25447 8270 25467
rect 8271 25464 8285 25467
rect 8340 25447 8342 25467
rect 8364 25447 8366 25467
rect 8367 25464 8381 25467
rect 8388 25464 8391 25467
rect 8436 25447 8438 25467
rect 8652 25447 8654 25467
rect 8700 25447 8702 25467
rect 8748 25447 8750 25467
rect 8820 25447 8822 25467
rect 8844 25447 8846 25467
rect 8868 25447 8870 25467
rect 9516 25447 9518 25467
rect 9660 25447 9662 25467
rect 9684 25447 9686 25467
rect 9756 25447 9758 25467
rect 9780 25447 9782 25467
rect 9804 25447 9806 25467
rect 9852 25447 9854 25467
rect 9900 25447 9902 25467
rect 9948 25447 9950 25467
rect 10068 25447 10070 25467
rect 10071 25464 10085 25467
rect 10092 25464 10095 25467
rect 10116 25447 10118 25467
rect 10164 25447 10166 25467
rect 10188 25447 10190 25467
rect 10212 25447 10214 25467
rect 10284 25447 10286 25467
rect 10332 25447 10334 25467
rect 10380 25447 10382 25467
rect 10383 25464 10397 25467
rect 10404 25464 10407 25467
rect 10428 25447 10430 25467
rect 10476 25447 10478 25467
rect 10500 25447 10502 25467
rect 10524 25447 10526 25467
rect 10572 25447 10574 25467
rect 10596 25447 10598 25467
rect 10620 25447 10622 25467
rect 10692 25447 10694 25467
rect 10716 25447 10718 25467
rect 10719 25464 10733 25467
rect 10743 25467 25619 25471
rect 10743 25464 10757 25467
rect 10788 25447 10790 25467
rect 10956 25447 10958 25467
rect 11004 25447 11006 25467
rect 11052 25447 11054 25467
rect 11100 25447 11102 25467
rect 11172 25447 11174 25467
rect 11220 25447 11222 25467
rect 11340 25447 11342 25467
rect 11436 25447 11438 25467
rect 11532 25447 11534 25467
rect 11580 25447 11582 25467
rect 11628 25447 11630 25467
rect 11676 25447 11678 25467
rect 11724 25447 11726 25467
rect 11772 25447 11774 25467
rect 11796 25447 11798 25467
rect 11892 25447 11894 25467
rect 11988 25447 11990 25467
rect 12060 25447 12062 25467
rect 12132 25447 12134 25467
rect 12228 25447 12230 25467
rect 12276 25447 12278 25467
rect 12324 25447 12326 25467
rect 12420 25447 12422 25467
rect 12444 25447 12446 25467
rect 12492 25447 12494 25467
rect 12516 25447 12518 25467
rect 12540 25447 12542 25467
rect 12588 25447 12590 25467
rect 12636 25447 12638 25467
rect 12732 25447 12734 25467
rect 12756 25447 12758 25467
rect 12804 25447 12806 25467
rect 12828 25447 12830 25467
rect 12852 25447 12854 25467
rect 12948 25447 12950 25467
rect 12972 25447 12974 25467
rect 13044 25447 13046 25467
rect 13068 25447 13070 25467
rect 13116 25447 13118 25467
rect 13284 25447 13286 25467
rect 13332 25447 13334 25467
rect 13572 25447 13574 25467
rect 13620 25447 13622 25467
rect 13668 25447 13670 25467
rect 13716 25447 13718 25467
rect 13764 25447 13766 25467
rect 13860 25447 13862 25467
rect 13956 25447 13958 25467
rect 14004 25447 14006 25467
rect 14100 25447 14102 25467
rect 15180 25447 15182 25467
rect 15276 25447 15278 25467
rect 15420 25447 15422 25467
rect 15492 25447 15494 25467
rect 15660 25447 15662 25467
rect 15708 25447 15710 25467
rect 15732 25447 15734 25467
rect 15756 25447 15758 25467
rect 15804 25447 15806 25467
rect 15828 25447 15830 25467
rect 15852 25447 15854 25467
rect 15900 25447 15902 25467
rect 15948 25447 15950 25467
rect 16044 25447 16046 25467
rect 16068 25447 16070 25467
rect 16164 25447 16166 25467
rect 16260 25447 16262 25467
rect 16308 25447 16310 25467
rect 16332 25447 16334 25467
rect 16356 25447 16358 25467
rect 16404 25447 16406 25467
rect 16452 25447 16454 25467
rect 16548 25447 16550 25467
rect 16572 25447 16574 25467
rect 16620 25447 16622 25467
rect 16668 25447 16670 25467
rect 16716 25447 16718 25467
rect 16764 25447 16766 25467
rect 16812 25447 16814 25467
rect 16884 25447 16886 25467
rect 16908 25447 16910 25467
rect 16980 25447 16982 25467
rect 17052 25447 17054 25467
rect 17196 25447 17198 25467
rect 17220 25447 17222 25467
rect 17292 25447 17294 25467
rect 17316 25447 17318 25467
rect 18084 25447 18086 25467
rect 18132 25447 18134 25467
rect 18228 25447 18230 25467
rect 18396 25447 18398 25467
rect 18492 25447 18494 25467
rect 18516 25447 18518 25467
rect 18564 25447 18566 25467
rect 18612 25447 18614 25467
rect 18660 25447 18662 25467
rect 18756 25447 18758 25467
rect 18841 25462 18844 25467
rect 18852 25462 18854 25467
rect 18851 25448 18854 25462
rect 18900 25447 18902 25467
rect 18924 25447 18927 25464
rect 18996 25447 18998 25467
rect 19020 25447 19022 25467
rect 19092 25447 19094 25467
rect 19116 25447 19118 25467
rect 19140 25447 19142 25467
rect 19188 25447 19190 25467
rect 19236 25447 19238 25467
rect 19332 25447 19334 25467
rect 19476 25447 19478 25467
rect 19788 25447 19790 25467
rect 19836 25447 19838 25467
rect 19860 25447 19862 25467
rect 19884 25447 19886 25467
rect 19932 25447 19934 25467
rect 19956 25447 19958 25467
rect 19980 25447 19982 25467
rect 20028 25447 20030 25467
rect 20052 25447 20054 25467
rect 20076 25447 20078 25467
rect 20148 25447 20150 25467
rect 20172 25447 20174 25467
rect 20196 25447 20198 25467
rect 20268 25447 20270 25467
rect 20292 25447 20294 25467
rect 20388 25447 20390 25467
rect 20412 25447 20414 25467
rect 20508 25447 20510 25467
rect 20556 25447 20558 25467
rect 20604 25447 20606 25467
rect 20916 25464 20918 25467
rect 20916 25447 20919 25464
rect 20964 25447 20966 25467
rect 21012 25447 21014 25467
rect 21060 25447 21062 25467
rect 21108 25447 21110 25467
rect 21204 25447 21206 25467
rect 21300 25447 21302 25467
rect 21324 25447 21326 25467
rect 21444 25447 21446 25467
rect 21468 25447 21470 25467
rect 21564 25447 21566 25467
rect 21588 25447 21590 25467
rect 21684 25447 21686 25467
rect 21708 25447 21710 25467
rect 21828 25447 21830 25467
rect 21924 25447 21926 25467
rect 22068 25447 22070 25467
rect 22188 25447 22190 25467
rect 22212 25447 22214 25467
rect 22884 25447 22886 25467
rect 22980 25447 22982 25467
rect 23076 25447 23078 25467
rect 23100 25447 23102 25467
rect 23124 25447 23126 25467
rect 23244 25447 23246 25467
rect 23340 25447 23342 25467
rect 23412 25447 23414 25467
rect 23460 25447 23462 25467
rect 23508 25447 23510 25467
rect 23556 25447 23558 25467
rect 23604 25447 23606 25467
rect 23652 25447 23654 25467
rect 23676 25447 23678 25467
rect 23772 25447 23774 25467
rect 23820 25447 23822 25467
rect 23916 25447 23918 25467
rect 24012 25447 24014 25467
rect 24060 25447 24062 25467
rect 24156 25447 24158 25467
rect 24492 25447 24494 25467
rect 24516 25447 24518 25467
rect 24588 25447 24590 25467
rect 24612 25447 24614 25467
rect 24684 25447 24686 25467
rect 24732 25447 24734 25467
rect 24756 25447 24758 25467
rect 24780 25447 24782 25467
rect 24852 25447 24854 25467
rect 24876 25447 24878 25467
rect 24972 25447 24974 25467
rect 25068 25447 25070 25467
rect 25164 25447 25166 25467
rect 25260 25447 25262 25467
rect 25284 25447 25286 25467
rect 25356 25447 25358 25467
rect 25380 25447 25382 25467
rect 25404 25447 25406 25467
rect 25500 25447 25502 25467
rect 25585 25462 25588 25467
rect 25596 25462 25598 25467
rect 25595 25448 25598 25462
rect 25561 25447 25595 25448
rect -14999 25443 -14011 25447
rect -14892 25440 -14890 25443
rect -14892 25424 -14889 25440
rect -14903 25423 -14869 25424
rect -14676 25423 -14674 25443
rect -14460 25423 -14458 25443
rect -14100 25423 -14098 25443
rect -14025 25440 -14011 25443
rect -14004 25443 -8131 25447
rect -14004 25440 -13987 25443
rect -14004 25423 -14002 25440
rect -13788 25423 -13786 25443
rect -13751 25423 -13717 25424
rect -13428 25423 -13426 25443
rect -12756 25423 -12754 25443
rect -12660 25423 -12658 25443
rect -12348 25423 -12346 25443
rect -12252 25423 -12250 25443
rect -12156 25423 -12154 25443
rect -12060 25423 -12058 25443
rect -11855 25438 -11852 25443
rect -11844 25438 -11842 25443
rect -11845 25424 -11842 25438
rect -11772 25423 -11769 25440
rect -11676 25423 -11674 25443
rect -11508 25423 -11506 25443
rect -11436 25423 -11434 25443
rect -11412 25423 -11410 25443
rect -11340 25423 -11338 25443
rect -11196 25423 -11194 25443
rect -11145 25440 -11131 25443
rect -11100 25423 -11098 25443
rect -10764 25423 -10762 25443
rect -10644 25423 -10642 25443
rect -9996 25423 -9994 25443
rect -9900 25423 -9898 25443
rect -9732 25423 -9730 25443
rect -9516 25423 -9514 25443
rect -9348 25423 -9346 25443
rect -9180 25423 -9178 25443
rect -8436 25423 -8434 25443
rect -8364 25423 -8362 25443
rect -8340 25423 -8338 25443
rect -8268 25423 -8266 25443
rect -8145 25440 -8131 25443
rect -8121 25443 -4291 25447
rect -8121 25440 -8107 25443
rect -8100 25440 -8097 25443
rect -8004 25423 -8002 25443
rect -7932 25423 -7930 25443
rect -7620 25423 -7618 25443
rect -7524 25423 -7522 25443
rect -7356 25423 -7354 25443
rect -7308 25423 -7306 25443
rect -7212 25423 -7210 25443
rect -7044 25423 -7042 25443
rect -6948 25423 -6946 25443
rect -6852 25423 -6850 25443
rect -6780 25423 -6778 25443
rect -6756 25423 -6754 25443
rect -6660 25423 -6658 25443
rect -6612 25423 -6610 25443
rect -6516 25423 -6514 25443
rect -6372 25423 -6370 25443
rect -6167 25438 -6164 25443
rect -6156 25438 -6154 25443
rect -6157 25424 -6154 25438
rect -6060 25440 -6058 25443
rect -6191 25423 -6157 25424
rect -6060 25423 -6057 25440
rect -6036 25423 -6034 25443
rect -5892 25423 -5890 25443
rect -5196 25423 -5194 25443
rect -5193 25440 -5179 25443
rect -5172 25440 -5169 25443
rect -5100 25423 -5098 25443
rect -5001 25440 -4987 25443
rect -4980 25440 -4977 25443
rect -4881 25440 -4867 25443
rect -4785 25440 -4771 25443
rect -4569 25440 -4555 25443
rect -4500 25423 -4498 25443
rect -4449 25440 -4435 25443
rect -4404 25423 -4402 25443
rect -4308 25423 -4306 25443
rect -4305 25440 -4291 25443
rect -4281 25443 18917 25447
rect -4281 25440 -4267 25443
rect -4260 25440 -4257 25443
rect -4164 25423 -4162 25443
rect -4020 25423 -4018 25443
rect -3876 25423 -3874 25443
rect -3732 25423 -3730 25443
rect -3564 25423 -3562 25443
rect -3516 25423 -3514 25443
rect -3468 25423 -3466 25443
rect -3420 25423 -3418 25443
rect -3324 25423 -3322 25443
rect -3228 25423 -3226 25443
rect -3132 25423 -3130 25443
rect -3108 25423 -3105 25440
rect -3012 25423 -3010 25443
rect -2964 25423 -2962 25443
rect -2916 25423 -2914 25443
rect -2892 25423 -2890 25443
rect -2868 25423 -2866 25443
rect -2820 25423 -2818 25443
rect -2796 25423 -2794 25443
rect -2772 25423 -2770 25443
rect -2676 25423 -2674 25443
rect -2580 25423 -2578 25443
rect -2364 25423 -2362 25443
rect -2316 25423 -2314 25443
rect -2268 25423 -2266 25443
rect -2244 25423 -2242 25443
rect -2172 25423 -2170 25443
rect -2148 25423 -2146 25443
rect -2076 25423 -2074 25443
rect -2052 25423 -2050 25443
rect -1980 25423 -1978 25443
rect -1884 25423 -1882 25443
rect -1572 25423 -1570 25443
rect -1476 25423 -1474 25443
rect -1380 25423 -1378 25443
rect -1356 25423 -1354 25443
rect -1308 25424 -1306 25443
rect -1343 25423 -1285 25424
rect -1260 25423 -1258 25443
rect -1140 25423 -1138 25443
rect -708 25423 -706 25443
rect -612 25423 -610 25443
rect -588 25423 -586 25443
rect -540 25423 -538 25443
rect -492 25423 -490 25443
rect -444 25423 -442 25443
rect -396 25423 -394 25443
rect -359 25438 -356 25443
rect -349 25424 -346 25438
rect -348 25423 -346 25424
rect -300 25423 -298 25443
rect -276 25423 -274 25443
rect -228 25440 -226 25443
rect -228 25423 -225 25440
rect -12 25423 -10 25443
rect 156 25423 158 25443
rect 204 25423 206 25443
rect 252 25423 254 25443
rect 348 25423 350 25443
rect 468 25423 470 25443
rect 492 25423 494 25443
rect 564 25423 566 25443
rect 588 25423 590 25443
rect 636 25423 638 25443
rect 660 25423 662 25443
rect 732 25423 734 25443
rect 1092 25423 1094 25443
rect 1140 25423 1142 25443
rect 1236 25423 1238 25443
rect 1308 25423 1310 25443
rect 1332 25423 1334 25443
rect 1380 25423 1382 25443
rect 1428 25423 1430 25443
rect 1476 25423 1478 25443
rect 1644 25424 1646 25443
rect 1633 25423 1667 25424
rect 1692 25423 1694 25443
rect 1740 25424 1742 25443
rect 1729 25423 1763 25424
rect 1788 25423 1790 25443
rect 2028 25423 2030 25443
rect 2076 25423 2078 25443
rect 2100 25423 2102 25443
rect 2124 25423 2126 25443
rect 2172 25423 2174 25443
rect 2220 25424 2222 25443
rect 2209 25423 2243 25424
rect 2316 25423 2318 25443
rect 2412 25423 2414 25443
rect 2460 25423 2462 25443
rect 2508 25423 2510 25443
rect 2580 25423 2582 25443
rect 2604 25423 2606 25443
rect 2676 25423 2678 25443
rect 2700 25424 2702 25443
rect 2689 25423 2723 25424
rect 2748 25423 2750 25443
rect 2772 25423 2774 25443
rect 2796 25424 2798 25443
rect 2785 25423 2819 25424
rect 2844 25423 2846 25443
rect 2868 25423 2870 25443
rect 2892 25423 2894 25443
rect 2940 25423 2942 25443
rect 3012 25423 3014 25443
rect 3108 25423 3110 25443
rect 3145 25423 3179 25424
rect 3252 25423 3254 25443
rect 3348 25423 3350 25443
rect 3396 25423 3398 25443
rect 3564 25423 3566 25443
rect 3636 25423 3638 25443
rect 3660 25423 3662 25443
rect 3732 25423 3734 25443
rect 3780 25423 3783 25440
rect 3828 25423 3830 25443
rect 3924 25423 3926 25443
rect 4020 25423 4022 25443
rect 4044 25423 4046 25443
rect 4092 25423 4094 25443
rect 4140 25423 4142 25443
rect 4188 25423 4190 25443
rect 4236 25423 4238 25443
rect 4308 25423 4310 25443
rect 4332 25423 4334 25443
rect 4404 25423 4406 25443
rect 4500 25423 4502 25443
rect 4596 25423 4598 25443
rect 4692 25423 4694 25443
rect 4860 25423 4862 25443
rect 4956 25423 4958 25443
rect 4980 25423 4982 25443
rect 5052 25423 5054 25443
rect 5124 25423 5126 25443
rect 5220 25423 5222 25443
rect 5268 25423 5270 25443
rect 5388 25423 5390 25443
rect 5484 25423 5486 25443
rect 5508 25423 5510 25443
rect 5532 25423 5534 25443
rect 5628 25423 5630 25443
rect 5652 25423 5654 25443
rect 5748 25423 5750 25443
rect 5796 25423 5798 25443
rect 5844 25423 5846 25443
rect 5892 25423 5894 25443
rect 6132 25423 6134 25443
rect 6180 25423 6182 25443
rect 6228 25423 6230 25443
rect 6252 25423 6254 25443
rect 6276 25423 6278 25443
rect 6324 25423 6326 25443
rect 6372 25423 6374 25443
rect 6409 25423 6467 25424
rect 6492 25423 6494 25443
rect 6588 25423 6590 25443
rect 6612 25423 6614 25443
rect 6660 25423 6662 25443
rect 6684 25423 6686 25443
rect 6708 25423 6710 25443
rect 6780 25423 6782 25443
rect 6804 25423 6806 25443
rect 6900 25423 6902 25443
rect 6924 25423 6926 25443
rect 7020 25423 7022 25443
rect 7068 25423 7070 25443
rect 7164 25423 7166 25443
rect 7236 25423 7238 25443
rect 7332 25423 7334 25443
rect 7380 25423 7382 25443
rect 7428 25423 7430 25443
rect 7452 25423 7454 25443
rect 7476 25423 7478 25443
rect 7524 25423 7526 25443
rect 7548 25423 7550 25443
rect 7572 25423 7574 25443
rect 7620 25423 7622 25443
rect 7644 25423 7646 25443
rect 7668 25423 7670 25443
rect 7956 25423 7958 25443
rect 8028 25423 8030 25443
rect 8124 25423 8126 25443
rect 8268 25423 8270 25443
rect 8340 25423 8342 25443
rect 8364 25423 8366 25443
rect 8436 25423 8438 25443
rect 8652 25423 8654 25443
rect 8700 25423 8702 25443
rect 8748 25423 8750 25443
rect 8820 25423 8822 25443
rect 8844 25423 8846 25443
rect 8868 25423 8870 25443
rect 9516 25423 9518 25443
rect 9660 25423 9662 25443
rect 9684 25423 9686 25443
rect 9756 25423 9758 25443
rect 9780 25423 9782 25443
rect 9804 25423 9806 25443
rect 9852 25423 9854 25443
rect 9900 25423 9902 25443
rect 9948 25423 9950 25443
rect 10068 25423 10070 25443
rect 10116 25423 10118 25443
rect 10164 25423 10166 25443
rect 10188 25423 10190 25443
rect 10212 25423 10214 25443
rect 10284 25423 10286 25443
rect 10332 25423 10334 25443
rect 10380 25423 10382 25443
rect 10428 25423 10430 25443
rect 10476 25423 10478 25443
rect 10500 25423 10502 25443
rect 10524 25423 10526 25443
rect 10572 25423 10574 25443
rect 10596 25423 10598 25443
rect 10620 25423 10622 25443
rect 10692 25423 10694 25443
rect 10716 25423 10718 25443
rect 10788 25423 10790 25443
rect 10956 25423 10958 25443
rect 11004 25423 11006 25443
rect 11052 25423 11054 25443
rect 11100 25423 11102 25443
rect 11172 25423 11174 25443
rect 11220 25423 11222 25443
rect 11340 25423 11342 25443
rect 11436 25423 11438 25443
rect 11532 25423 11534 25443
rect 11580 25423 11582 25443
rect 11628 25423 11630 25443
rect 11676 25423 11678 25443
rect 11724 25423 11726 25443
rect 11772 25423 11774 25443
rect 11796 25423 11798 25443
rect 11892 25423 11894 25443
rect 11988 25423 11990 25443
rect 12060 25423 12062 25443
rect 12132 25423 12134 25443
rect 12228 25423 12230 25443
rect 12276 25423 12278 25443
rect 12324 25423 12326 25443
rect 12420 25423 12422 25443
rect 12444 25423 12446 25443
rect 12492 25423 12494 25443
rect 12516 25423 12518 25443
rect 12540 25423 12542 25443
rect 12588 25423 12590 25443
rect 12636 25423 12638 25443
rect 12732 25423 12734 25443
rect 12756 25423 12758 25443
rect 12804 25423 12806 25443
rect 12828 25423 12830 25443
rect 12852 25423 12854 25443
rect 12948 25423 12950 25443
rect 12972 25423 12974 25443
rect 13044 25423 13046 25443
rect 13068 25423 13070 25443
rect 13116 25423 13118 25443
rect 13284 25423 13286 25443
rect 13332 25423 13334 25443
rect 13572 25423 13574 25443
rect 13620 25423 13622 25443
rect 13668 25423 13670 25443
rect 13716 25423 13718 25443
rect 13764 25423 13766 25443
rect 13860 25423 13862 25443
rect 13956 25423 13958 25443
rect 14004 25423 14006 25443
rect 14100 25423 14102 25443
rect 15180 25423 15182 25443
rect 15276 25423 15278 25443
rect 15420 25423 15422 25443
rect 15492 25423 15494 25443
rect 15660 25423 15662 25443
rect 15708 25423 15710 25443
rect 15732 25423 15734 25443
rect 15756 25423 15758 25443
rect 15804 25423 15806 25443
rect 15828 25423 15830 25443
rect 15852 25423 15854 25443
rect 15900 25423 15902 25443
rect 15948 25423 15950 25443
rect 16044 25423 16046 25443
rect 16068 25423 16070 25443
rect 16164 25423 16166 25443
rect 16260 25423 16262 25443
rect 16308 25423 16310 25443
rect 16332 25423 16334 25443
rect 16356 25423 16358 25443
rect 16404 25423 16406 25443
rect 16452 25423 16454 25443
rect 16548 25423 16550 25443
rect 16572 25423 16574 25443
rect 16620 25423 16622 25443
rect 16668 25423 16670 25443
rect 16716 25423 16718 25443
rect 16764 25423 16766 25443
rect 16812 25423 16814 25443
rect 16884 25423 16886 25443
rect 16908 25423 16910 25443
rect 16921 25423 16979 25424
rect 16980 25423 16982 25443
rect 17052 25423 17054 25443
rect 17196 25423 17198 25443
rect 17220 25423 17222 25443
rect 17292 25423 17294 25443
rect 17316 25423 17318 25443
rect 18084 25423 18086 25443
rect 18132 25423 18134 25443
rect 18228 25423 18230 25443
rect 18396 25423 18398 25443
rect 18492 25423 18494 25443
rect 18516 25423 18518 25443
rect 18564 25423 18566 25443
rect 18612 25423 18614 25443
rect 18660 25423 18662 25443
rect 18756 25423 18758 25443
rect 18900 25423 18902 25443
rect 18903 25440 18917 25443
rect 18924 25443 20885 25447
rect 18924 25440 18941 25443
rect 18924 25423 18926 25440
rect 18996 25423 18998 25443
rect 19020 25423 19022 25443
rect 19092 25423 19094 25443
rect 19116 25423 19118 25443
rect 19140 25423 19142 25443
rect 19188 25423 19190 25443
rect 19236 25423 19238 25443
rect 19332 25423 19334 25443
rect 19476 25423 19478 25443
rect 19788 25423 19790 25443
rect 19836 25423 19838 25443
rect 19860 25423 19862 25443
rect 19884 25423 19886 25443
rect 19932 25423 19934 25443
rect 19956 25423 19958 25443
rect 19980 25423 19982 25443
rect 20028 25423 20030 25443
rect 20052 25423 20054 25443
rect 20076 25423 20078 25443
rect 20148 25423 20150 25443
rect 20172 25423 20174 25443
rect 20196 25423 20198 25443
rect 20268 25423 20270 25443
rect 20292 25423 20294 25443
rect 20388 25423 20390 25443
rect 20412 25423 20414 25443
rect 20508 25423 20510 25443
rect 20556 25423 20558 25443
rect 20604 25423 20606 25443
rect 20871 25440 20885 25443
rect 20895 25443 25595 25447
rect 20895 25440 20909 25443
rect 20916 25440 20919 25443
rect 20964 25423 20966 25443
rect 21012 25423 21014 25443
rect 21060 25424 21062 25443
rect 21025 25423 21083 25424
rect 21108 25423 21110 25443
rect 21204 25423 21206 25443
rect 21300 25423 21302 25443
rect 21324 25423 21326 25443
rect 21444 25423 21446 25443
rect 21468 25423 21470 25443
rect 21564 25423 21566 25443
rect 21588 25423 21590 25443
rect 21684 25423 21686 25443
rect 21708 25423 21710 25443
rect 21828 25423 21830 25443
rect 21924 25423 21926 25443
rect 22068 25423 22070 25443
rect 22188 25423 22190 25443
rect 22212 25423 22214 25443
rect 22884 25423 22886 25443
rect 22980 25423 22982 25443
rect 23076 25423 23078 25443
rect 23100 25423 23102 25443
rect 23124 25423 23126 25443
rect 23244 25423 23246 25443
rect 23340 25423 23342 25443
rect 23412 25423 23414 25443
rect 23460 25423 23462 25443
rect 23508 25423 23510 25443
rect 23556 25423 23558 25443
rect 23604 25423 23606 25443
rect 23652 25423 23654 25443
rect 23676 25423 23678 25443
rect 23772 25423 23774 25443
rect 23820 25423 23822 25443
rect 23916 25423 23918 25443
rect 24012 25423 24014 25443
rect 24060 25423 24062 25443
rect 24156 25423 24158 25443
rect 24492 25423 24494 25443
rect 24516 25423 24518 25443
rect 24588 25423 24590 25443
rect 24612 25423 24614 25443
rect 24684 25423 24686 25443
rect 24732 25423 24734 25443
rect 24756 25423 24758 25443
rect 24780 25423 24782 25443
rect 24852 25423 24854 25443
rect 24876 25423 24878 25443
rect 24972 25423 24974 25443
rect 25068 25423 25070 25443
rect 25164 25423 25166 25443
rect 25260 25423 25262 25443
rect 25284 25423 25286 25443
rect 25356 25423 25358 25443
rect 25380 25423 25382 25443
rect 25404 25424 25406 25443
rect 25500 25424 25502 25443
rect 25393 25423 25451 25424
rect 25489 25423 25523 25424
rect -14903 25419 -11779 25423
rect -14903 25416 -14899 25419
rect -14892 25416 -14889 25419
rect -14783 25399 -14749 25400
rect -14676 25399 -14674 25419
rect -14460 25399 -14458 25419
rect -14100 25399 -14098 25419
rect -14004 25399 -14002 25419
rect -13788 25399 -13786 25419
rect -13428 25399 -13426 25419
rect -12756 25399 -12754 25419
rect -12660 25399 -12658 25419
rect -12348 25399 -12346 25419
rect -12252 25399 -12250 25419
rect -12156 25399 -12154 25419
rect -12060 25399 -12058 25419
rect -11793 25416 -11779 25419
rect -11772 25419 -3115 25423
rect -11772 25416 -11755 25419
rect -11772 25399 -11770 25416
rect -11676 25399 -11674 25419
rect -11508 25399 -11506 25419
rect -11436 25399 -11434 25419
rect -11412 25399 -11410 25419
rect -11340 25399 -11338 25419
rect -11196 25399 -11194 25419
rect -11100 25399 -11098 25419
rect -10764 25399 -10762 25419
rect -10644 25399 -10642 25419
rect -9996 25399 -9994 25419
rect -9900 25399 -9898 25419
rect -9732 25399 -9730 25419
rect -9516 25399 -9514 25419
rect -9348 25399 -9346 25419
rect -9335 25399 -9277 25400
rect -9180 25399 -9178 25419
rect -8577 25416 -8563 25419
rect -8436 25399 -8434 25419
rect -8364 25399 -8362 25419
rect -8340 25399 -8338 25419
rect -8268 25399 -8266 25419
rect -8004 25399 -8002 25419
rect -7932 25399 -7930 25419
rect -7620 25399 -7618 25419
rect -7524 25399 -7522 25419
rect -7356 25399 -7354 25419
rect -7308 25399 -7306 25419
rect -7212 25399 -7210 25419
rect -7044 25399 -7042 25419
rect -6948 25399 -6946 25419
rect -6852 25399 -6850 25419
rect -6780 25399 -6778 25419
rect -6756 25399 -6754 25419
rect -6660 25399 -6658 25419
rect -6612 25399 -6610 25419
rect -6516 25399 -6514 25419
rect -6372 25399 -6370 25419
rect -6081 25416 -6067 25419
rect -6060 25416 -6057 25419
rect -6036 25399 -6034 25419
rect -5892 25399 -5890 25419
rect -5196 25399 -5194 25419
rect -5100 25399 -5098 25419
rect -4500 25399 -4498 25419
rect -4404 25399 -4402 25419
rect -4308 25399 -4306 25419
rect -4164 25399 -4162 25419
rect -4020 25399 -4018 25419
rect -3876 25399 -3874 25419
rect -3732 25399 -3730 25419
rect -3671 25399 -3589 25400
rect -3564 25399 -3562 25419
rect -3516 25399 -3514 25419
rect -3468 25399 -3466 25419
rect -3420 25399 -3418 25419
rect -3324 25399 -3322 25419
rect -3228 25399 -3226 25419
rect -3132 25399 -3130 25419
rect -3129 25416 -3115 25419
rect -3108 25419 -259 25423
rect -3108 25416 -3091 25419
rect -3108 25399 -3106 25416
rect -3012 25399 -3010 25419
rect -2964 25399 -2962 25419
rect -2916 25399 -2914 25419
rect -2892 25399 -2890 25419
rect -2868 25399 -2866 25419
rect -2820 25399 -2818 25419
rect -2796 25399 -2794 25419
rect -2772 25399 -2770 25419
rect -2676 25399 -2674 25419
rect -2580 25399 -2578 25419
rect -2364 25399 -2362 25419
rect -2316 25399 -2314 25419
rect -2268 25399 -2266 25419
rect -2244 25399 -2242 25419
rect -2172 25399 -2170 25419
rect -2148 25399 -2146 25419
rect -2076 25399 -2074 25419
rect -2052 25399 -2050 25419
rect -1980 25399 -1978 25419
rect -1884 25399 -1882 25419
rect -1857 25416 -1843 25419
rect -1572 25399 -1570 25419
rect -1476 25399 -1474 25419
rect -1380 25399 -1378 25419
rect -1356 25399 -1354 25419
rect -1319 25414 -1316 25419
rect -1308 25414 -1306 25419
rect -1309 25400 -1306 25414
rect -1260 25399 -1258 25419
rect -1236 25399 -1233 25416
rect -1140 25399 -1138 25419
rect -708 25399 -706 25419
rect -612 25399 -610 25419
rect -588 25399 -586 25419
rect -540 25399 -538 25419
rect -492 25399 -490 25419
rect -444 25399 -442 25419
rect -396 25399 -394 25419
rect -348 25399 -346 25419
rect -300 25399 -298 25419
rect -276 25399 -274 25419
rect -273 25416 -259 25419
rect -249 25419 3773 25423
rect -249 25416 -235 25419
rect -228 25416 -225 25419
rect -12 25399 -10 25419
rect 156 25399 158 25419
rect 204 25399 206 25419
rect 252 25399 254 25419
rect 348 25399 350 25419
rect 468 25399 470 25419
rect 492 25399 494 25419
rect 564 25399 566 25419
rect 588 25399 590 25419
rect 636 25399 638 25419
rect 660 25399 662 25419
rect 732 25399 734 25419
rect 1092 25399 1094 25419
rect 1140 25399 1142 25419
rect 1236 25399 1238 25419
rect 1308 25399 1310 25419
rect 1332 25399 1334 25419
rect 1380 25399 1382 25419
rect 1428 25399 1430 25419
rect 1476 25399 1478 25419
rect 1633 25414 1636 25419
rect 1644 25414 1646 25419
rect 1643 25400 1646 25414
rect 1692 25399 1694 25419
rect 1729 25414 1732 25419
rect 1740 25416 1742 25419
rect 1740 25414 1743 25416
rect 1739 25400 1743 25414
rect 1788 25399 1790 25419
rect 2028 25399 2030 25419
rect 2076 25399 2078 25419
rect 2100 25399 2102 25419
rect 2124 25399 2126 25419
rect 2172 25399 2174 25419
rect 2209 25414 2212 25419
rect 2220 25414 2222 25419
rect 2219 25400 2222 25414
rect 2316 25416 2318 25419
rect 2316 25399 2319 25416
rect 2412 25399 2414 25419
rect 2460 25399 2462 25419
rect 2508 25399 2510 25419
rect 2580 25399 2582 25419
rect 2604 25399 2606 25419
rect 2676 25399 2678 25419
rect 2689 25414 2692 25419
rect 2700 25414 2702 25419
rect 2699 25400 2702 25414
rect 2748 25400 2750 25419
rect 2713 25399 2771 25400
rect 2772 25399 2774 25419
rect 2785 25414 2788 25419
rect 2796 25416 2798 25419
rect 2796 25414 2799 25416
rect 2795 25400 2799 25414
rect 2844 25399 2846 25419
rect 2868 25399 2870 25419
rect 2892 25416 2894 25419
rect 2892 25399 2895 25416
rect 2940 25399 2942 25419
rect 3012 25399 3014 25419
rect 3108 25399 3110 25419
rect 3252 25416 3254 25419
rect 3252 25399 3255 25416
rect 3348 25399 3350 25419
rect 3396 25399 3398 25419
rect 3564 25399 3566 25419
rect 3636 25399 3638 25419
rect 3660 25399 3662 25419
rect 3732 25399 3734 25419
rect 3759 25416 3773 25419
rect 3780 25419 25523 25423
rect 3780 25416 3797 25419
rect 3780 25399 3782 25416
rect 3828 25399 3830 25419
rect 3924 25399 3926 25419
rect 4020 25399 4022 25419
rect 4044 25399 4046 25419
rect 4092 25399 4094 25419
rect 4140 25399 4142 25419
rect 4188 25399 4190 25419
rect 4236 25399 4238 25419
rect 4308 25399 4310 25419
rect 4332 25399 4334 25419
rect 4404 25399 4406 25419
rect 4500 25399 4502 25419
rect 4596 25399 4598 25419
rect 4692 25399 4694 25419
rect 4860 25399 4862 25419
rect 4956 25399 4958 25419
rect 4980 25399 4982 25419
rect 5052 25399 5054 25419
rect 5124 25399 5126 25419
rect 5220 25399 5222 25419
rect 5268 25399 5270 25419
rect 5388 25399 5390 25419
rect 5484 25399 5486 25419
rect 5508 25399 5510 25419
rect 5532 25399 5534 25419
rect 5628 25399 5630 25419
rect 5652 25399 5654 25419
rect 5748 25399 5750 25419
rect 5796 25399 5798 25419
rect 5844 25399 5846 25419
rect 5892 25399 5894 25419
rect 6073 25399 6107 25400
rect 6132 25399 6134 25419
rect 6180 25399 6182 25419
rect 6228 25399 6230 25419
rect 6252 25399 6254 25419
rect 6276 25399 6278 25419
rect 6324 25399 6326 25419
rect 6372 25399 6374 25419
rect 6409 25414 6412 25419
rect 6419 25400 6422 25414
rect 6420 25399 6422 25400
rect 6492 25399 6494 25419
rect 6516 25399 6519 25416
rect 6588 25399 6590 25419
rect 6612 25399 6614 25419
rect 6660 25399 6662 25419
rect 6684 25399 6686 25419
rect 6708 25399 6710 25419
rect 6780 25399 6782 25419
rect 6804 25399 6806 25419
rect 6900 25399 6902 25419
rect 6924 25399 6926 25419
rect 7020 25399 7022 25419
rect 7068 25399 7070 25419
rect 7164 25399 7166 25419
rect 7236 25399 7238 25419
rect 7332 25399 7334 25419
rect 7380 25399 7382 25419
rect 7428 25399 7430 25419
rect 7452 25399 7454 25419
rect 7476 25399 7478 25419
rect 7524 25399 7526 25419
rect 7548 25399 7550 25419
rect 7572 25399 7574 25419
rect 7620 25399 7622 25419
rect 7644 25399 7646 25419
rect 7668 25399 7670 25419
rect 7956 25399 7958 25419
rect 8028 25399 8030 25419
rect 8124 25399 8126 25419
rect 8268 25399 8270 25419
rect 8340 25399 8342 25419
rect 8364 25399 8366 25419
rect 8436 25399 8438 25419
rect 8652 25399 8654 25419
rect 8700 25399 8702 25419
rect 8748 25399 8750 25419
rect 8820 25399 8822 25419
rect 8844 25399 8846 25419
rect 8868 25399 8870 25419
rect 9516 25399 9518 25419
rect 9660 25399 9662 25419
rect 9684 25399 9686 25419
rect 9756 25399 9758 25419
rect 9780 25399 9782 25419
rect 9804 25399 9806 25419
rect 9852 25399 9854 25419
rect 9900 25399 9902 25419
rect 9948 25399 9950 25419
rect 10068 25400 10070 25419
rect 10033 25399 10091 25400
rect 10116 25399 10118 25419
rect 10164 25399 10166 25419
rect 10188 25399 10190 25419
rect 10212 25399 10214 25419
rect 10284 25399 10286 25419
rect 10332 25399 10334 25419
rect 10380 25399 10382 25419
rect 10428 25399 10430 25419
rect 10476 25399 10478 25419
rect 10500 25399 10502 25419
rect 10524 25399 10526 25419
rect 10572 25399 10574 25419
rect 10596 25399 10598 25419
rect 10620 25399 10622 25419
rect 10692 25399 10694 25419
rect 10716 25399 10718 25419
rect 10788 25399 10790 25419
rect 10956 25399 10958 25419
rect 11004 25399 11006 25419
rect 11052 25399 11054 25419
rect 11100 25399 11102 25419
rect 11172 25399 11174 25419
rect 11220 25399 11222 25419
rect 11340 25399 11342 25419
rect 11436 25399 11438 25419
rect 11532 25399 11534 25419
rect 11580 25399 11582 25419
rect 11628 25399 11630 25419
rect 11676 25399 11678 25419
rect 11724 25399 11726 25419
rect 11772 25399 11774 25419
rect 11796 25399 11798 25419
rect 11892 25399 11894 25419
rect 11988 25399 11990 25419
rect 12060 25399 12062 25419
rect 12132 25399 12134 25419
rect 12228 25399 12230 25419
rect 12276 25399 12278 25419
rect 12324 25399 12326 25419
rect 12420 25399 12422 25419
rect 12444 25399 12446 25419
rect 12492 25399 12494 25419
rect 12516 25399 12518 25419
rect 12540 25399 12542 25419
rect 12588 25399 12590 25419
rect 12636 25399 12638 25419
rect 12732 25399 12734 25419
rect 12756 25399 12758 25419
rect 12804 25399 12806 25419
rect 12828 25399 12830 25419
rect 12852 25399 12854 25419
rect 12948 25399 12950 25419
rect 12972 25399 12974 25419
rect 13044 25399 13046 25419
rect 13068 25399 13070 25419
rect 13116 25399 13118 25419
rect 13284 25399 13286 25419
rect 13332 25399 13334 25419
rect 13572 25399 13574 25419
rect 13620 25399 13622 25419
rect 13668 25399 13670 25419
rect 13716 25399 13718 25419
rect 13764 25399 13766 25419
rect 13860 25399 13862 25419
rect 13956 25399 13958 25419
rect 14004 25399 14006 25419
rect 14100 25399 14102 25419
rect 15180 25399 15182 25419
rect 15276 25399 15278 25419
rect 15420 25399 15422 25419
rect 15492 25399 15494 25419
rect 15660 25399 15662 25419
rect 15708 25399 15710 25419
rect 15732 25399 15734 25419
rect 15756 25399 15758 25419
rect 15804 25399 15806 25419
rect 15828 25399 15830 25419
rect 15852 25399 15854 25419
rect 15900 25399 15902 25419
rect 15948 25399 15950 25419
rect 16044 25399 16046 25419
rect 16068 25399 16070 25419
rect 16164 25399 16166 25419
rect 16260 25399 16262 25419
rect 16308 25399 16310 25419
rect 16332 25399 16334 25419
rect 16356 25399 16358 25419
rect 16404 25399 16406 25419
rect 16452 25399 16454 25419
rect 16548 25399 16550 25419
rect 16572 25399 16574 25419
rect 16620 25399 16622 25419
rect 16668 25399 16670 25419
rect 16716 25399 16718 25419
rect 16764 25399 16766 25419
rect 16812 25399 16814 25419
rect 16884 25399 16886 25419
rect 16908 25399 16910 25419
rect 16980 25399 16982 25419
rect 17052 25416 17054 25419
rect 17052 25399 17055 25416
rect 17137 25399 17195 25400
rect 17196 25399 17198 25419
rect 17220 25399 17222 25419
rect 17292 25399 17294 25419
rect 17316 25399 17318 25419
rect 18084 25399 18086 25419
rect 18132 25399 18134 25419
rect 18228 25399 18230 25419
rect 18396 25399 18398 25419
rect 18492 25399 18494 25419
rect 18516 25399 18518 25419
rect 18564 25399 18566 25419
rect 18612 25399 18614 25419
rect 18660 25399 18662 25419
rect 18756 25399 18758 25419
rect 18900 25399 18902 25419
rect 18924 25399 18926 25419
rect 18996 25399 18998 25419
rect 19020 25399 19022 25419
rect 19092 25399 19094 25419
rect 19116 25399 19118 25419
rect 19140 25399 19142 25419
rect 19188 25399 19190 25419
rect 19236 25399 19238 25419
rect 19332 25399 19334 25419
rect 19369 25399 19403 25400
rect 19476 25399 19478 25419
rect 19788 25399 19790 25419
rect 19836 25399 19838 25419
rect 19860 25399 19862 25419
rect 19884 25399 19886 25419
rect 19932 25399 19934 25419
rect 19956 25399 19958 25419
rect 19980 25399 19982 25419
rect 20028 25399 20030 25419
rect 20052 25399 20054 25419
rect 20076 25399 20078 25419
rect 20148 25399 20150 25419
rect 20172 25399 20174 25419
rect 20196 25399 20198 25419
rect 20268 25399 20270 25419
rect 20292 25399 20294 25419
rect 20388 25399 20390 25419
rect 20412 25399 20414 25419
rect 20425 25399 20483 25400
rect 20508 25399 20510 25419
rect 20556 25399 20558 25419
rect 20604 25399 20606 25419
rect 20964 25399 20966 25419
rect 21012 25399 21014 25419
rect 21049 25414 21052 25419
rect 21060 25414 21062 25419
rect 21059 25400 21062 25414
rect 21108 25399 21110 25419
rect 21204 25399 21206 25419
rect 21300 25399 21302 25419
rect 21324 25399 21326 25419
rect 21444 25399 21446 25419
rect 21468 25399 21470 25419
rect 21564 25399 21566 25419
rect 21588 25399 21590 25419
rect 21684 25399 21686 25419
rect 21708 25399 21710 25419
rect 21828 25399 21830 25419
rect 21924 25399 21926 25419
rect 22068 25399 22070 25419
rect 22188 25399 22190 25419
rect 22212 25399 22214 25419
rect 22884 25399 22886 25419
rect 22980 25399 22982 25419
rect 23076 25399 23078 25419
rect 23100 25399 23102 25419
rect 23124 25399 23126 25419
rect 23244 25399 23246 25419
rect 23340 25399 23342 25419
rect 23412 25399 23414 25419
rect 23460 25399 23462 25419
rect 23508 25399 23510 25419
rect 23556 25399 23558 25419
rect 23604 25399 23606 25419
rect 23652 25399 23654 25419
rect 23676 25399 23678 25419
rect 23772 25399 23774 25419
rect 23820 25399 23822 25419
rect 23916 25399 23918 25419
rect 24012 25399 24014 25419
rect 24060 25399 24062 25419
rect 24156 25399 24158 25419
rect 24492 25399 24494 25419
rect 24516 25399 24518 25419
rect 24588 25399 24590 25419
rect 24612 25399 24614 25419
rect 24684 25399 24686 25419
rect 24732 25399 24734 25419
rect 24756 25399 24758 25419
rect 24780 25399 24782 25419
rect 24852 25399 24854 25419
rect 24876 25399 24878 25419
rect 24972 25399 24974 25419
rect 25068 25399 25070 25419
rect 25164 25399 25166 25419
rect 25260 25399 25262 25419
rect 25284 25399 25286 25419
rect 25356 25399 25358 25419
rect 25380 25400 25382 25419
rect 25393 25414 25396 25419
rect 25404 25414 25406 25419
rect 25489 25414 25492 25419
rect 25500 25416 25502 25419
rect 25500 25414 25503 25416
rect 25403 25400 25406 25414
rect 25499 25406 25503 25414
rect 25513 25406 25517 25414
rect 25499 25400 25513 25406
rect 25369 25399 25403 25400
rect -14783 25395 -1243 25399
rect -14676 25392 -14674 25395
rect -14676 25376 -14673 25392
rect -14687 25375 -14653 25376
rect -14460 25375 -14458 25395
rect -14100 25375 -14098 25395
rect -14004 25375 -14002 25395
rect -13788 25375 -13786 25395
rect -13665 25392 -13651 25395
rect -13428 25375 -13426 25395
rect -13391 25375 -13357 25376
rect -12756 25375 -12754 25395
rect -12660 25376 -12658 25395
rect -12671 25375 -12637 25376
rect -12348 25375 -12346 25395
rect -12252 25375 -12250 25395
rect -12156 25375 -12154 25395
rect -12060 25375 -12058 25395
rect -11772 25375 -11770 25395
rect -11676 25375 -11674 25395
rect -11508 25375 -11506 25395
rect -11436 25375 -11434 25395
rect -11412 25375 -11410 25395
rect -11340 25375 -11338 25395
rect -11196 25375 -11194 25395
rect -11100 25375 -11098 25395
rect -10764 25375 -10762 25395
rect -10644 25375 -10642 25395
rect -9996 25375 -9994 25395
rect -9900 25375 -9898 25395
rect -9732 25375 -9730 25395
rect -9516 25375 -9514 25395
rect -9348 25375 -9346 25395
rect -9228 25375 -9225 25392
rect -9180 25375 -9178 25395
rect -8436 25375 -8434 25395
rect -8364 25375 -8362 25395
rect -8340 25375 -8338 25395
rect -8268 25375 -8266 25395
rect -8004 25375 -8002 25395
rect -7932 25375 -7930 25395
rect -7620 25375 -7618 25395
rect -7524 25375 -7522 25395
rect -7356 25375 -7354 25395
rect -7308 25375 -7306 25395
rect -7212 25375 -7210 25395
rect -7044 25375 -7042 25395
rect -6948 25375 -6946 25395
rect -6887 25375 -6853 25376
rect -6852 25375 -6850 25395
rect -6780 25375 -6778 25395
rect -6756 25375 -6754 25395
rect -6660 25375 -6658 25395
rect -6612 25375 -6610 25395
rect -6516 25375 -6514 25395
rect -6372 25375 -6370 25395
rect -6105 25392 -6091 25395
rect -6036 25375 -6034 25395
rect -5892 25375 -5890 25395
rect -5196 25375 -5194 25395
rect -5100 25375 -5098 25395
rect -4823 25375 -4765 25376
rect -4500 25375 -4498 25395
rect -4404 25375 -4402 25395
rect -4308 25375 -4306 25395
rect -4164 25375 -4162 25395
rect -4020 25375 -4018 25395
rect -3876 25375 -3874 25395
rect -3732 25375 -3730 25395
rect -3647 25390 -3644 25395
rect -3564 25392 -3562 25395
rect -3516 25392 -3514 25395
rect -3637 25376 -3634 25390
rect -3636 25375 -3634 25376
rect -3564 25375 -3561 25392
rect -3516 25375 -3513 25392
rect -3468 25375 -3466 25395
rect -3420 25375 -3418 25395
rect -3324 25375 -3322 25395
rect -3228 25375 -3226 25395
rect -3132 25375 -3130 25395
rect -3108 25375 -3106 25395
rect -3012 25375 -3010 25395
rect -2964 25375 -2962 25395
rect -2916 25375 -2914 25395
rect -2892 25375 -2890 25395
rect -2868 25375 -2866 25395
rect -2820 25375 -2818 25395
rect -2796 25375 -2794 25395
rect -2772 25375 -2770 25395
rect -2676 25375 -2674 25395
rect -2580 25375 -2578 25395
rect -2364 25375 -2362 25395
rect -2316 25375 -2314 25395
rect -2268 25375 -2266 25395
rect -2244 25375 -2242 25395
rect -2172 25375 -2170 25395
rect -2148 25375 -2146 25395
rect -2076 25375 -2074 25395
rect -2052 25375 -2050 25395
rect -1980 25375 -1978 25395
rect -1884 25375 -1882 25395
rect -1572 25375 -1570 25395
rect -1476 25375 -1474 25395
rect -1380 25375 -1378 25395
rect -1356 25375 -1354 25395
rect -1260 25375 -1258 25395
rect -1257 25392 -1243 25395
rect -1236 25395 6509 25399
rect -1236 25392 -1219 25395
rect -1236 25375 -1234 25392
rect -1140 25375 -1138 25395
rect -708 25375 -706 25395
rect -695 25375 -613 25376
rect -612 25375 -610 25395
rect -588 25375 -586 25395
rect -540 25375 -538 25395
rect -492 25375 -490 25395
rect -444 25375 -442 25395
rect -396 25375 -394 25395
rect -348 25375 -346 25395
rect -300 25375 -298 25395
rect -276 25375 -274 25395
rect -12 25375 -10 25395
rect 156 25375 158 25395
rect 204 25375 206 25395
rect 252 25375 254 25395
rect 348 25375 350 25395
rect 468 25375 470 25395
rect 492 25375 494 25395
rect 564 25375 566 25395
rect 588 25375 590 25395
rect 636 25375 638 25395
rect 660 25375 662 25395
rect 732 25375 734 25395
rect 1092 25375 1094 25395
rect 1140 25375 1142 25395
rect 1236 25375 1238 25395
rect 1308 25375 1310 25395
rect 1332 25375 1334 25395
rect 1380 25375 1382 25395
rect 1428 25375 1430 25395
rect 1476 25375 1478 25395
rect 1692 25375 1694 25395
rect 1719 25392 1733 25395
rect 1788 25375 1790 25395
rect 1815 25392 1829 25395
rect 2028 25375 2030 25395
rect 2076 25375 2078 25395
rect 2100 25375 2102 25395
rect 2124 25375 2126 25395
rect 2172 25376 2174 25395
rect 2295 25392 2309 25395
rect 2316 25392 2319 25395
rect 2137 25375 2195 25376
rect 2412 25375 2414 25395
rect 2460 25375 2462 25395
rect 2508 25375 2510 25395
rect 2580 25375 2582 25395
rect 2604 25375 2606 25395
rect 2676 25375 2678 25395
rect 2737 25390 2740 25395
rect 2748 25390 2750 25395
rect 2747 25376 2750 25390
rect 2772 25375 2774 25395
rect 2775 25392 2789 25395
rect 2844 25392 2846 25395
rect 2844 25375 2847 25392
rect 2868 25375 2870 25395
rect 2871 25392 2885 25395
rect 2892 25392 2895 25395
rect 2940 25375 2942 25395
rect 3012 25375 3014 25395
rect 3108 25375 3110 25395
rect 3231 25392 3245 25395
rect 3252 25392 3255 25395
rect 3348 25375 3350 25395
rect 3396 25375 3398 25395
rect 3564 25375 3566 25395
rect 3636 25375 3638 25395
rect 3660 25375 3662 25395
rect 3732 25375 3734 25395
rect 3780 25375 3782 25395
rect 3828 25375 3830 25395
rect 3924 25375 3926 25395
rect 4020 25375 4022 25395
rect 4044 25375 4046 25395
rect 4092 25375 4094 25395
rect 4140 25375 4142 25395
rect 4188 25375 4190 25395
rect 4236 25375 4238 25395
rect 4308 25375 4310 25395
rect 4332 25375 4334 25395
rect 4404 25375 4406 25395
rect 4500 25375 4502 25395
rect 4596 25375 4598 25395
rect 4692 25375 4694 25395
rect 4860 25375 4862 25395
rect 4956 25375 4958 25395
rect 4980 25375 4982 25395
rect 5052 25375 5054 25395
rect 5124 25375 5126 25395
rect 5220 25375 5222 25395
rect 5268 25375 5270 25395
rect 5388 25375 5390 25395
rect 5484 25375 5486 25395
rect 5508 25375 5510 25395
rect 5532 25375 5534 25395
rect 5628 25375 5630 25395
rect 5652 25375 5654 25395
rect 5748 25375 5750 25395
rect 5796 25375 5798 25395
rect 5844 25375 5846 25395
rect 5892 25375 5894 25395
rect 6132 25375 6134 25395
rect 6180 25392 6182 25395
rect 6180 25375 6183 25392
rect 6228 25375 6230 25395
rect 6252 25375 6254 25395
rect 6276 25375 6278 25395
rect 6324 25375 6326 25395
rect 6372 25375 6374 25395
rect 6420 25375 6422 25395
rect 6492 25375 6494 25395
rect 6495 25392 6509 25395
rect 6516 25395 17021 25399
rect 6516 25392 6533 25395
rect 6516 25375 6518 25392
rect 6588 25375 6590 25395
rect 6612 25375 6614 25395
rect 6660 25375 6662 25395
rect 6684 25375 6686 25395
rect 6708 25375 6710 25395
rect 6780 25375 6782 25395
rect 6804 25375 6806 25395
rect 6900 25375 6902 25395
rect 6924 25375 6926 25395
rect 6937 25375 6995 25376
rect 7020 25375 7022 25395
rect 7068 25375 7070 25395
rect 7164 25375 7166 25395
rect 7236 25375 7238 25395
rect 7332 25375 7334 25395
rect 7380 25375 7382 25395
rect 7428 25375 7430 25395
rect 7452 25375 7454 25395
rect 7476 25375 7478 25395
rect 7524 25375 7526 25395
rect 7548 25375 7550 25395
rect 7572 25375 7574 25395
rect 7620 25375 7622 25395
rect 7644 25375 7646 25395
rect 7668 25375 7670 25395
rect 7956 25375 7958 25395
rect 8028 25375 8030 25395
rect 8124 25375 8126 25395
rect 8268 25375 8270 25395
rect 8340 25375 8342 25395
rect 8364 25375 8366 25395
rect 8436 25375 8438 25395
rect 8652 25375 8654 25395
rect 8700 25375 8702 25395
rect 8748 25375 8750 25395
rect 8820 25375 8822 25395
rect 8844 25375 8846 25395
rect 8868 25375 8870 25395
rect 9516 25375 9518 25395
rect 9660 25375 9662 25395
rect 9684 25375 9686 25395
rect 9756 25375 9758 25395
rect 9780 25375 9782 25395
rect 9804 25375 9806 25395
rect 9852 25375 9854 25395
rect 9900 25375 9902 25395
rect 9948 25375 9950 25395
rect 10033 25390 10036 25395
rect 10057 25390 10060 25395
rect 10068 25390 10070 25395
rect 10043 25376 10046 25390
rect 10067 25376 10070 25390
rect 10044 25375 10046 25376
rect 10116 25375 10118 25395
rect 10164 25392 10166 25395
rect 10164 25375 10167 25392
rect 10188 25375 10190 25395
rect 10212 25375 10214 25395
rect 10284 25375 10286 25395
rect 10332 25375 10334 25395
rect 10380 25375 10382 25395
rect 10428 25375 10430 25395
rect 10476 25375 10478 25395
rect 10500 25375 10502 25395
rect 10524 25375 10526 25395
rect 10572 25375 10574 25395
rect 10596 25375 10598 25395
rect 10620 25375 10622 25395
rect 10692 25375 10694 25395
rect 10716 25375 10718 25395
rect 10788 25375 10790 25395
rect 10956 25375 10958 25395
rect 11004 25375 11006 25395
rect 11052 25375 11054 25395
rect 11100 25375 11102 25395
rect 11172 25375 11174 25395
rect 11220 25375 11222 25395
rect 11340 25375 11342 25395
rect 11436 25375 11438 25395
rect 11532 25375 11534 25395
rect 11580 25375 11582 25395
rect 11628 25375 11630 25395
rect 11676 25375 11678 25395
rect 11724 25375 11726 25395
rect 11772 25375 11774 25395
rect 11796 25375 11798 25395
rect 11892 25375 11894 25395
rect 11988 25375 11990 25395
rect 12060 25375 12062 25395
rect 12132 25375 12134 25395
rect 12228 25375 12230 25395
rect 12276 25375 12278 25395
rect 12324 25375 12326 25395
rect 12420 25375 12422 25395
rect 12444 25375 12446 25395
rect 12492 25375 12494 25395
rect 12516 25375 12518 25395
rect 12540 25375 12542 25395
rect 12588 25375 12590 25395
rect 12636 25375 12638 25395
rect 12732 25375 12734 25395
rect 12756 25375 12758 25395
rect 12804 25375 12806 25395
rect 12828 25375 12830 25395
rect 12852 25376 12854 25395
rect 12841 25375 12875 25376
rect 12948 25375 12950 25395
rect 12972 25375 12974 25395
rect 13044 25375 13046 25395
rect 13068 25375 13070 25395
rect 13116 25375 13118 25395
rect 13284 25375 13286 25395
rect 13332 25375 13334 25395
rect 13572 25375 13574 25395
rect 13620 25375 13622 25395
rect 13668 25375 13670 25395
rect 13716 25375 13718 25395
rect 13764 25375 13766 25395
rect 13860 25375 13862 25395
rect 13956 25375 13958 25395
rect 14004 25375 14006 25395
rect 14100 25375 14102 25395
rect 15145 25375 15179 25376
rect 15180 25375 15182 25395
rect 15276 25375 15278 25395
rect 15420 25375 15422 25395
rect 15492 25375 15494 25395
rect 15660 25375 15662 25395
rect 15708 25375 15710 25395
rect 15732 25375 15734 25395
rect 15756 25375 15758 25395
rect 15804 25375 15806 25395
rect 15828 25375 15830 25395
rect 15852 25375 15854 25395
rect 15900 25375 15902 25395
rect 15948 25375 15950 25395
rect 16044 25375 16046 25395
rect 16068 25375 16070 25395
rect 16164 25375 16166 25395
rect 16260 25375 16262 25395
rect 16308 25375 16310 25395
rect 16332 25375 16334 25395
rect 16356 25376 16358 25395
rect 16345 25375 16379 25376
rect 16404 25375 16406 25395
rect 16452 25375 16454 25395
rect 16548 25375 16550 25395
rect 16572 25375 16574 25395
rect 16620 25375 16622 25395
rect 16668 25375 16670 25395
rect 16716 25375 16718 25395
rect 16764 25375 16766 25395
rect 16812 25375 16814 25395
rect 16884 25375 16886 25395
rect 16908 25375 16910 25395
rect 16980 25375 16982 25395
rect 17007 25392 17021 25395
rect 17031 25395 21125 25399
rect 17031 25392 17045 25395
rect 17052 25392 17055 25395
rect 17137 25390 17140 25395
rect 17147 25376 17150 25390
rect 17148 25375 17150 25376
rect 17196 25375 17198 25395
rect 17220 25375 17222 25395
rect 17292 25375 17294 25395
rect 17316 25375 17318 25395
rect 18084 25376 18086 25395
rect 18049 25375 18107 25376
rect 18132 25375 18134 25395
rect 18228 25375 18230 25395
rect 18396 25375 18398 25395
rect 18492 25375 18494 25395
rect 18516 25375 18518 25395
rect 18564 25375 18566 25395
rect 18612 25375 18614 25395
rect 18660 25375 18662 25395
rect 18756 25375 18758 25395
rect 18900 25375 18902 25395
rect 18924 25375 18926 25395
rect 18996 25375 18998 25395
rect 19020 25375 19022 25395
rect 19092 25375 19094 25395
rect 19116 25375 19118 25395
rect 19140 25375 19142 25395
rect 19188 25375 19190 25395
rect 19236 25375 19238 25395
rect 19332 25375 19334 25395
rect 19476 25392 19478 25395
rect 19476 25375 19479 25392
rect 19788 25375 19790 25395
rect 19836 25375 19838 25395
rect 19860 25375 19862 25395
rect 19884 25375 19886 25395
rect 19932 25375 19934 25395
rect 19956 25375 19958 25395
rect 19980 25375 19982 25395
rect 20028 25375 20030 25395
rect 20052 25375 20054 25395
rect 20076 25375 20078 25395
rect 20148 25375 20150 25395
rect 20172 25375 20174 25395
rect 20196 25375 20198 25395
rect 20268 25375 20270 25395
rect 20292 25375 20294 25395
rect 20388 25375 20390 25395
rect 20412 25375 20414 25395
rect 20508 25375 20510 25395
rect 20556 25392 20558 25395
rect 20556 25375 20559 25392
rect 20604 25375 20606 25395
rect 20964 25375 20966 25395
rect 21012 25375 21014 25395
rect 21108 25375 21110 25395
rect 21111 25392 21125 25395
rect 21135 25395 25403 25399
rect 21135 25392 21149 25395
rect 21204 25375 21206 25395
rect 21300 25375 21302 25395
rect 21324 25375 21326 25395
rect 21444 25375 21446 25395
rect 21468 25375 21470 25395
rect 21564 25375 21566 25395
rect 21588 25375 21590 25395
rect 21684 25375 21686 25395
rect 21708 25375 21710 25395
rect 21828 25375 21830 25395
rect 21924 25375 21926 25395
rect 22068 25375 22070 25395
rect 22188 25375 22190 25395
rect 22212 25375 22214 25395
rect 22884 25375 22886 25395
rect 22980 25375 22982 25395
rect 23076 25375 23078 25395
rect 23100 25375 23102 25395
rect 23124 25375 23126 25395
rect 23244 25375 23246 25395
rect 23340 25375 23342 25395
rect 23412 25375 23414 25395
rect 23460 25375 23462 25395
rect 23508 25375 23510 25395
rect 23556 25375 23558 25395
rect 23604 25375 23606 25395
rect 23652 25375 23654 25395
rect 23676 25375 23678 25395
rect 23689 25375 23747 25376
rect 23772 25375 23774 25395
rect 23820 25375 23822 25395
rect 23916 25375 23918 25395
rect 24012 25375 24014 25395
rect 24060 25375 24062 25395
rect 24156 25375 24158 25395
rect 24492 25375 24494 25395
rect 24516 25375 24518 25395
rect 24588 25375 24590 25395
rect 24612 25375 24614 25395
rect 24684 25375 24686 25395
rect 24732 25375 24734 25395
rect 24756 25375 24758 25395
rect 24780 25375 24782 25395
rect 24852 25375 24854 25395
rect 24876 25375 24878 25395
rect 24972 25375 24974 25395
rect 25068 25375 25070 25395
rect 25164 25375 25166 25395
rect 25260 25375 25262 25395
rect 25284 25376 25286 25395
rect 25356 25376 25358 25395
rect 25369 25390 25372 25395
rect 25380 25390 25382 25395
rect 25379 25376 25382 25390
rect 25273 25375 25331 25376
rect 25345 25375 25379 25376
rect -14687 25371 -9235 25375
rect -14687 25368 -14683 25371
rect -14676 25368 -14673 25371
rect -14567 25351 -14533 25352
rect -14460 25351 -14458 25371
rect -14100 25351 -14098 25371
rect -14004 25351 -14002 25371
rect -13788 25351 -13786 25371
rect -13428 25351 -13426 25371
rect -12756 25351 -12754 25371
rect -12671 25366 -12668 25371
rect -12660 25366 -12658 25371
rect -12661 25352 -12658 25366
rect -12743 25351 -12685 25352
rect -12348 25351 -12346 25371
rect -12252 25351 -12250 25371
rect -12156 25351 -12154 25371
rect -12060 25351 -12058 25371
rect -11772 25351 -11770 25371
rect -11676 25351 -11674 25371
rect -11508 25351 -11506 25371
rect -11436 25351 -11434 25371
rect -11412 25351 -11410 25371
rect -11340 25351 -11338 25371
rect -11196 25351 -11194 25371
rect -11100 25351 -11098 25371
rect -10764 25351 -10762 25371
rect -10644 25351 -10642 25371
rect -9996 25351 -9994 25371
rect -9900 25351 -9898 25371
rect -9732 25351 -9730 25371
rect -9516 25352 -9514 25371
rect -9551 25351 -9493 25352
rect -9348 25351 -9346 25371
rect -9249 25368 -9235 25371
rect -9228 25371 -3547 25375
rect -9228 25368 -9211 25371
rect -9228 25351 -9226 25368
rect -9180 25352 -9178 25371
rect -9215 25351 -9157 25352
rect -8436 25351 -8434 25371
rect -8364 25351 -8362 25371
rect -8340 25351 -8338 25371
rect -8268 25351 -8266 25371
rect -8004 25351 -8002 25371
rect -7932 25351 -7930 25371
rect -7620 25351 -7618 25371
rect -7524 25351 -7522 25371
rect -7356 25351 -7354 25371
rect -7308 25351 -7306 25371
rect -7212 25351 -7210 25371
rect -7044 25351 -7042 25371
rect -6948 25351 -6946 25371
rect -6852 25351 -6850 25371
rect -6780 25368 -6778 25371
rect -6780 25351 -6777 25368
rect -6756 25351 -6754 25371
rect -6660 25351 -6658 25371
rect -6612 25351 -6610 25371
rect -6516 25351 -6514 25371
rect -6372 25351 -6370 25371
rect -6036 25351 -6034 25371
rect -5892 25351 -5890 25371
rect -5196 25351 -5194 25371
rect -5100 25351 -5098 25371
rect -4716 25351 -4713 25368
rect -4500 25351 -4498 25371
rect -4404 25351 -4402 25371
rect -4308 25351 -4306 25371
rect -4164 25351 -4162 25371
rect -4020 25351 -4018 25371
rect -3876 25351 -3874 25371
rect -3732 25351 -3730 25371
rect -3636 25351 -3634 25371
rect -3585 25368 -3571 25371
rect -3564 25368 -3547 25371
rect -3537 25371 2813 25375
rect -3537 25368 -3523 25371
rect -3516 25368 -3513 25371
rect -3551 25351 -3493 25352
rect -3468 25351 -3466 25371
rect -3420 25351 -3418 25371
rect -3324 25351 -3322 25371
rect -3228 25351 -3226 25371
rect -3132 25351 -3130 25371
rect -3108 25351 -3106 25371
rect -3012 25351 -3010 25371
rect -2964 25351 -2962 25371
rect -2916 25351 -2914 25371
rect -2892 25351 -2890 25371
rect -2868 25351 -2866 25371
rect -2820 25351 -2818 25371
rect -2796 25351 -2794 25371
rect -2772 25351 -2770 25371
rect -2676 25351 -2674 25371
rect -2580 25351 -2578 25371
rect -2364 25351 -2362 25371
rect -2316 25351 -2314 25371
rect -2268 25351 -2266 25371
rect -2244 25351 -2242 25371
rect -2172 25351 -2170 25371
rect -2148 25351 -2146 25371
rect -2076 25351 -2074 25371
rect -2052 25351 -2050 25371
rect -1980 25351 -1978 25371
rect -1884 25351 -1882 25371
rect -1572 25351 -1570 25371
rect -1476 25351 -1474 25371
rect -1380 25351 -1378 25371
rect -1356 25351 -1354 25371
rect -1260 25351 -1258 25371
rect -1236 25351 -1234 25371
rect -1140 25351 -1138 25371
rect -708 25351 -706 25371
rect -671 25366 -668 25371
rect -661 25352 -658 25366
rect -660 25351 -658 25352
rect -612 25351 -610 25371
rect -588 25368 -586 25371
rect -540 25368 -538 25371
rect -588 25351 -585 25368
rect -540 25351 -537 25368
rect -492 25351 -490 25371
rect -444 25351 -442 25371
rect -396 25351 -394 25371
rect -348 25351 -346 25371
rect -300 25351 -298 25371
rect -276 25351 -274 25371
rect -12 25351 -10 25371
rect 156 25351 158 25371
rect 204 25351 206 25371
rect 252 25351 254 25371
rect 348 25351 350 25371
rect 468 25351 470 25371
rect 492 25351 494 25371
rect 564 25351 566 25371
rect 588 25351 590 25371
rect 636 25351 638 25371
rect 660 25351 662 25371
rect 732 25351 734 25371
rect 1092 25351 1094 25371
rect 1140 25351 1142 25371
rect 1236 25351 1238 25371
rect 1308 25351 1310 25371
rect 1332 25351 1334 25371
rect 1380 25351 1382 25371
rect 1428 25351 1430 25371
rect 1476 25351 1478 25371
rect 1692 25351 1694 25371
rect 1788 25351 1790 25371
rect 2028 25351 2030 25371
rect 2076 25351 2078 25371
rect 2100 25351 2102 25371
rect 2124 25351 2126 25371
rect 2161 25366 2164 25371
rect 2172 25366 2174 25371
rect 2171 25352 2174 25366
rect 2244 25351 2247 25368
rect 2412 25351 2414 25371
rect 2460 25351 2462 25371
rect 2508 25351 2510 25371
rect 2580 25351 2582 25371
rect 2604 25351 2606 25371
rect 2676 25351 2678 25371
rect 2772 25351 2774 25371
rect 2799 25368 2813 25371
rect 2823 25371 10133 25375
rect 2823 25368 2837 25371
rect 2844 25368 2847 25371
rect 2868 25351 2870 25371
rect 2940 25351 2942 25371
rect 3012 25351 3014 25371
rect 3108 25351 3110 25371
rect 3348 25351 3350 25371
rect 3396 25351 3398 25371
rect 3564 25351 3566 25371
rect 3636 25351 3638 25371
rect 3660 25351 3662 25371
rect 3732 25351 3734 25371
rect 3780 25351 3782 25371
rect 3828 25351 3830 25371
rect 3924 25351 3926 25371
rect 4020 25351 4022 25371
rect 4044 25351 4046 25371
rect 4092 25351 4094 25371
rect 4140 25351 4142 25371
rect 4188 25351 4190 25371
rect 4236 25351 4238 25371
rect 4308 25351 4310 25371
rect 4332 25351 4334 25371
rect 4404 25351 4406 25371
rect 4500 25351 4502 25371
rect 4596 25351 4598 25371
rect 4692 25351 4694 25371
rect 4860 25351 4862 25371
rect 4956 25351 4958 25371
rect 4980 25351 4982 25371
rect 5052 25351 5054 25371
rect 5124 25351 5126 25371
rect 5220 25351 5222 25371
rect 5268 25351 5270 25371
rect 5388 25351 5390 25371
rect 5484 25351 5486 25371
rect 5508 25351 5510 25371
rect 5532 25351 5534 25371
rect 5628 25351 5630 25371
rect 5652 25351 5654 25371
rect 5748 25351 5750 25371
rect 5796 25351 5798 25371
rect 5844 25351 5846 25371
rect 5892 25351 5894 25371
rect 6132 25351 6134 25371
rect 6159 25368 6173 25371
rect 6180 25368 6183 25371
rect 6228 25351 6230 25371
rect 6252 25351 6254 25371
rect 6276 25351 6278 25371
rect 6324 25351 6326 25371
rect 6372 25351 6374 25371
rect 6420 25351 6422 25371
rect 6492 25351 6494 25371
rect 6516 25351 6518 25371
rect 6588 25351 6590 25371
rect 6612 25351 6614 25371
rect 6660 25351 6662 25371
rect 6684 25351 6686 25371
rect 6708 25351 6710 25371
rect 6780 25351 6782 25371
rect 6804 25351 6806 25371
rect 6900 25351 6902 25371
rect 6924 25351 6926 25371
rect 7020 25351 7022 25371
rect 7068 25368 7070 25371
rect 7068 25351 7071 25368
rect 7164 25351 7166 25371
rect 7236 25351 7238 25371
rect 7332 25351 7334 25371
rect 7380 25351 7382 25371
rect 7428 25351 7430 25371
rect 7452 25351 7454 25371
rect 7476 25351 7478 25371
rect 7524 25351 7526 25371
rect 7548 25351 7550 25371
rect 7572 25351 7574 25371
rect 7620 25351 7622 25371
rect 7644 25351 7646 25371
rect 7668 25351 7670 25371
rect 7897 25351 7955 25352
rect 7956 25351 7958 25371
rect 8028 25351 8030 25371
rect 8124 25351 8126 25371
rect 8268 25351 8270 25371
rect 8340 25351 8342 25371
rect 8364 25351 8366 25371
rect 8436 25351 8438 25371
rect 8652 25351 8654 25371
rect 8700 25351 8702 25371
rect 8748 25351 8750 25371
rect 8820 25351 8822 25371
rect 8844 25351 8846 25371
rect 8868 25351 8870 25371
rect 9516 25351 9518 25371
rect 9660 25351 9662 25371
rect 9684 25351 9686 25371
rect 9756 25351 9758 25371
rect 9780 25351 9782 25371
rect 9804 25351 9806 25371
rect 9852 25351 9854 25371
rect 9900 25351 9902 25371
rect 9948 25351 9950 25371
rect 10044 25351 10046 25371
rect 10116 25351 10118 25371
rect 10119 25368 10133 25371
rect 10143 25371 17237 25375
rect 10143 25368 10157 25371
rect 10164 25368 10167 25371
rect 10188 25351 10190 25371
rect 10212 25351 10214 25371
rect 10284 25351 10286 25371
rect 10332 25351 10334 25371
rect 10380 25351 10382 25371
rect 10428 25351 10430 25371
rect 10476 25351 10478 25371
rect 10500 25351 10502 25371
rect 10524 25351 10526 25371
rect 10572 25351 10574 25371
rect 10596 25351 10598 25371
rect 10620 25351 10622 25371
rect 10692 25351 10694 25371
rect 10716 25351 10718 25371
rect 10788 25351 10790 25371
rect 10956 25351 10958 25371
rect 11004 25351 11006 25371
rect 11052 25351 11054 25371
rect 11100 25351 11102 25371
rect 11172 25351 11174 25371
rect 11220 25351 11222 25371
rect 11340 25351 11342 25371
rect 11436 25351 11438 25371
rect 11532 25351 11534 25371
rect 11580 25351 11582 25371
rect 11628 25351 11630 25371
rect 11676 25351 11678 25371
rect 11724 25351 11726 25371
rect 11772 25351 11774 25371
rect 11796 25351 11798 25371
rect 11892 25351 11894 25371
rect 11988 25351 11990 25371
rect 12060 25351 12062 25371
rect 12132 25351 12134 25371
rect 12228 25351 12230 25371
rect 12276 25351 12278 25371
rect 12324 25351 12326 25371
rect 12420 25351 12422 25371
rect 12444 25351 12446 25371
rect 12492 25351 12494 25371
rect 12516 25351 12518 25371
rect 12540 25351 12542 25371
rect 12588 25351 12590 25371
rect 12636 25351 12638 25371
rect 12732 25351 12734 25371
rect 12756 25351 12758 25371
rect 12804 25351 12806 25371
rect 12828 25351 12830 25371
rect 12841 25366 12844 25371
rect 12852 25366 12854 25371
rect 12851 25352 12854 25366
rect 12948 25368 12950 25371
rect 12948 25351 12951 25368
rect 12972 25351 12974 25371
rect 13044 25351 13046 25371
rect 13068 25351 13070 25371
rect 13116 25351 13118 25371
rect 13284 25351 13286 25371
rect 13332 25351 13334 25371
rect 13572 25351 13574 25371
rect 13620 25351 13622 25371
rect 13668 25351 13670 25371
rect 13716 25351 13718 25371
rect 13764 25351 13766 25371
rect 13860 25351 13862 25371
rect 13956 25351 13958 25371
rect 14004 25351 14006 25371
rect 14100 25351 14102 25371
rect 15180 25351 15182 25371
rect 15276 25351 15278 25371
rect 15420 25351 15422 25371
rect 15492 25351 15494 25371
rect 15660 25351 15662 25371
rect 15708 25351 15710 25371
rect 15732 25351 15734 25371
rect 15756 25351 15758 25371
rect 15804 25351 15806 25371
rect 15828 25351 15830 25371
rect 15852 25351 15854 25371
rect 15900 25351 15902 25371
rect 15948 25351 15950 25371
rect 16044 25351 16046 25371
rect 16068 25351 16070 25371
rect 16164 25351 16166 25371
rect 16260 25351 16262 25371
rect 16308 25351 16310 25371
rect 16332 25351 16334 25371
rect 16345 25366 16348 25371
rect 16356 25366 16358 25371
rect 16355 25352 16358 25366
rect 16404 25351 16406 25371
rect 16452 25368 16454 25371
rect 16452 25351 16455 25368
rect 16548 25351 16550 25371
rect 16572 25351 16574 25371
rect 16620 25351 16622 25371
rect 16668 25351 16670 25371
rect 16716 25351 16718 25371
rect 16764 25351 16766 25371
rect 16812 25351 16814 25371
rect 16884 25351 16886 25371
rect 16908 25351 16910 25371
rect 16980 25351 16982 25371
rect 17148 25351 17150 25371
rect 17196 25351 17198 25371
rect 17220 25351 17222 25371
rect 17223 25368 17237 25371
rect 17247 25371 20525 25375
rect 17247 25368 17261 25371
rect 17292 25351 17294 25371
rect 17316 25351 17318 25371
rect 18073 25366 18076 25371
rect 18084 25366 18086 25371
rect 18083 25352 18086 25366
rect 18132 25351 18134 25371
rect 18228 25351 18230 25371
rect 18396 25351 18398 25371
rect 18492 25351 18494 25371
rect 18516 25351 18518 25371
rect 18564 25351 18566 25371
rect 18612 25351 18614 25371
rect 18660 25351 18662 25371
rect 18756 25351 18758 25371
rect 18900 25351 18902 25371
rect 18924 25351 18926 25371
rect 18996 25351 18998 25371
rect 19020 25351 19022 25371
rect 19092 25351 19094 25371
rect 19116 25351 19118 25371
rect 19140 25351 19142 25371
rect 19188 25351 19190 25371
rect 19236 25351 19238 25371
rect 19332 25351 19334 25371
rect 19455 25368 19469 25371
rect 19476 25368 19479 25371
rect 19788 25351 19790 25371
rect 19836 25351 19838 25371
rect 19860 25351 19862 25371
rect 19884 25351 19886 25371
rect 19932 25351 19934 25371
rect 19956 25351 19958 25371
rect 19980 25351 19982 25371
rect 20028 25351 20030 25371
rect 20052 25351 20054 25371
rect 20076 25351 20078 25371
rect 20148 25351 20150 25371
rect 20172 25351 20174 25371
rect 20196 25351 20198 25371
rect 20268 25351 20270 25371
rect 20292 25351 20294 25371
rect 20388 25351 20390 25371
rect 20412 25351 20414 25371
rect 20508 25351 20510 25371
rect 20511 25368 20525 25371
rect 20535 25371 25379 25375
rect 20535 25368 20549 25371
rect 20556 25368 20559 25371
rect 20604 25351 20606 25371
rect 20964 25351 20966 25371
rect 21012 25351 21014 25371
rect 21108 25351 21110 25371
rect 21204 25351 21206 25371
rect 21300 25351 21302 25371
rect 21324 25351 21326 25371
rect 21444 25351 21446 25371
rect 21468 25351 21470 25371
rect 21564 25351 21566 25371
rect 21588 25351 21590 25371
rect 21684 25351 21686 25371
rect 21708 25351 21710 25371
rect 21828 25351 21830 25371
rect 21924 25351 21926 25371
rect 22068 25351 22070 25371
rect 22188 25351 22190 25371
rect 22212 25351 22214 25371
rect 22884 25351 22886 25371
rect 22980 25351 22982 25371
rect 23076 25351 23078 25371
rect 23100 25351 23102 25371
rect 23124 25351 23126 25371
rect 23244 25351 23246 25371
rect 23340 25351 23342 25371
rect 23412 25351 23414 25371
rect 23460 25351 23462 25371
rect 23508 25351 23510 25371
rect 23556 25351 23558 25371
rect 23604 25351 23606 25371
rect 23652 25351 23654 25371
rect 23676 25351 23678 25371
rect 23689 25366 23692 25371
rect 23699 25352 23702 25366
rect 23700 25351 23702 25352
rect 23772 25351 23774 25371
rect 23820 25368 23822 25371
rect 23796 25351 23799 25368
rect 23820 25351 23823 25368
rect 23916 25351 23918 25371
rect 24012 25351 24014 25371
rect 24060 25351 24062 25371
rect 24156 25351 24158 25371
rect 24492 25351 24494 25371
rect 24516 25351 24518 25371
rect 24588 25351 24590 25371
rect 24612 25351 24614 25371
rect 24684 25351 24686 25371
rect 24732 25351 24734 25371
rect 24756 25351 24758 25371
rect 24780 25351 24782 25371
rect 24852 25351 24854 25371
rect 24876 25351 24878 25371
rect 24972 25352 24974 25371
rect 25068 25352 25070 25371
rect 25164 25352 25166 25371
rect 25260 25352 25262 25371
rect 25273 25366 25276 25371
rect 25284 25366 25286 25371
rect 25345 25366 25348 25371
rect 25356 25366 25358 25371
rect 25283 25352 25286 25366
rect 25355 25352 25358 25366
rect 25369 25358 25373 25366
rect 25359 25352 25369 25358
rect 24961 25351 24995 25352
rect -14567 25347 -4723 25351
rect -14460 25344 -14458 25347
rect -14460 25328 -14457 25344
rect -14471 25327 -14437 25328
rect -14100 25327 -14098 25347
rect -14004 25327 -14002 25347
rect -13788 25327 -13786 25347
rect -13727 25327 -13693 25328
rect -13428 25327 -13426 25347
rect -13305 25344 -13291 25347
rect -12756 25327 -12754 25347
rect -12585 25344 -12571 25347
rect -12636 25327 -12633 25344
rect -12348 25327 -12346 25347
rect -12252 25327 -12250 25347
rect -12156 25327 -12154 25347
rect -12060 25327 -12058 25347
rect -11772 25327 -11770 25347
rect -11676 25327 -11674 25347
rect -11508 25327 -11506 25347
rect -11436 25327 -11434 25347
rect -11412 25327 -11410 25347
rect -11340 25327 -11338 25347
rect -11196 25327 -11194 25347
rect -11100 25327 -11098 25347
rect -10764 25327 -10762 25347
rect -10644 25327 -10642 25347
rect -9996 25327 -9994 25347
rect -9900 25327 -9898 25347
rect -9732 25327 -9730 25347
rect -9527 25342 -9524 25347
rect -9516 25342 -9514 25347
rect -9517 25328 -9514 25342
rect -9444 25327 -9441 25344
rect -9348 25327 -9346 25347
rect -9228 25327 -9226 25347
rect -9191 25342 -9188 25347
rect -9180 25342 -9178 25347
rect -9181 25328 -9178 25342
rect -9108 25327 -9105 25344
rect -8436 25327 -8434 25347
rect -8364 25327 -8362 25347
rect -8340 25327 -8338 25347
rect -8268 25327 -8266 25347
rect -8004 25327 -8002 25347
rect -7932 25327 -7930 25347
rect -7620 25327 -7618 25347
rect -7524 25327 -7522 25347
rect -7356 25327 -7354 25347
rect -7308 25327 -7306 25347
rect -7212 25327 -7210 25347
rect -7044 25327 -7042 25347
rect -6948 25327 -6946 25347
rect -6852 25327 -6850 25347
rect -6801 25344 -6787 25347
rect -6780 25344 -6777 25347
rect -6756 25327 -6754 25347
rect -6660 25327 -6658 25347
rect -6612 25327 -6610 25347
rect -6516 25327 -6514 25347
rect -6372 25327 -6370 25347
rect -6036 25327 -6034 25347
rect -5892 25327 -5890 25347
rect -5196 25327 -5194 25347
rect -5100 25327 -5098 25347
rect -4737 25344 -4723 25347
rect -4716 25347 -571 25351
rect -4716 25344 -4699 25347
rect -4716 25327 -4714 25344
rect -4500 25327 -4498 25347
rect -4404 25327 -4402 25347
rect -4308 25327 -4306 25347
rect -4164 25327 -4162 25347
rect -4020 25327 -4018 25347
rect -3876 25327 -3874 25347
rect -3732 25327 -3730 25347
rect -3636 25327 -3634 25347
rect -3551 25342 -3548 25347
rect -3541 25328 -3538 25342
rect -3540 25327 -3538 25328
rect -3468 25327 -3466 25347
rect -3420 25344 -3418 25347
rect -3420 25327 -3417 25344
rect -3324 25327 -3322 25347
rect -3228 25327 -3226 25347
rect -3132 25327 -3130 25347
rect -3108 25327 -3106 25347
rect -3012 25327 -3010 25347
rect -2964 25327 -2962 25347
rect -2916 25327 -2914 25347
rect -2892 25327 -2890 25347
rect -2868 25327 -2866 25347
rect -2820 25327 -2818 25347
rect -2796 25327 -2794 25347
rect -2772 25327 -2770 25347
rect -2676 25327 -2674 25347
rect -2580 25327 -2578 25347
rect -2364 25327 -2362 25347
rect -2316 25327 -2314 25347
rect -2268 25327 -2266 25347
rect -2244 25327 -2242 25347
rect -2172 25327 -2170 25347
rect -2148 25327 -2146 25347
rect -2076 25327 -2074 25347
rect -2052 25327 -2050 25347
rect -1980 25327 -1978 25347
rect -1884 25327 -1882 25347
rect -1572 25327 -1570 25347
rect -1476 25327 -1474 25347
rect -1380 25328 -1378 25347
rect -1391 25327 -1357 25328
rect -1356 25327 -1354 25347
rect -1260 25327 -1258 25347
rect -1236 25327 -1234 25347
rect -1140 25327 -1138 25347
rect -708 25327 -706 25347
rect -660 25327 -658 25347
rect -612 25327 -610 25347
rect -609 25344 -595 25347
rect -588 25344 -571 25347
rect -561 25347 2237 25351
rect -561 25344 -547 25347
rect -540 25344 -537 25347
rect -492 25327 -490 25347
rect -444 25327 -442 25347
rect -396 25327 -394 25347
rect -348 25327 -346 25347
rect -300 25327 -298 25347
rect -276 25327 -274 25347
rect -12 25327 -10 25347
rect 156 25327 158 25347
rect 204 25327 206 25347
rect 252 25327 254 25347
rect 348 25327 350 25347
rect 468 25327 470 25347
rect 492 25327 494 25347
rect 564 25327 566 25347
rect 588 25327 590 25347
rect 636 25327 638 25347
rect 660 25327 662 25347
rect 732 25327 734 25347
rect 1092 25327 1094 25347
rect 1140 25327 1142 25347
rect 1236 25327 1238 25347
rect 1308 25327 1310 25347
rect 1332 25327 1334 25347
rect 1380 25327 1382 25347
rect 1428 25327 1430 25347
rect 1476 25327 1478 25347
rect 1692 25327 1694 25347
rect 1788 25327 1790 25347
rect 2028 25327 2030 25347
rect 2076 25327 2078 25347
rect 2100 25327 2102 25347
rect 2124 25327 2126 25347
rect 2223 25344 2237 25347
rect 2244 25347 7037 25351
rect 2244 25344 2261 25347
rect 2244 25327 2246 25344
rect 2412 25327 2414 25347
rect 2460 25327 2462 25347
rect 2508 25327 2510 25347
rect 2580 25328 2582 25347
rect 2569 25327 2603 25328
rect 2604 25327 2606 25347
rect 2676 25327 2678 25347
rect 2772 25327 2774 25347
rect 2868 25327 2870 25347
rect 2940 25327 2942 25347
rect 3012 25327 3014 25347
rect 3108 25327 3110 25347
rect 3348 25327 3350 25347
rect 3396 25327 3398 25347
rect 3564 25327 3566 25347
rect 3636 25327 3638 25347
rect 3660 25327 3662 25347
rect 3732 25327 3734 25347
rect 3780 25327 3782 25347
rect 3828 25327 3830 25347
rect 3924 25327 3926 25347
rect 4020 25327 4022 25347
rect 4044 25327 4046 25347
rect 4092 25327 4094 25347
rect 4140 25327 4142 25347
rect 4188 25327 4190 25347
rect 4236 25327 4238 25347
rect 4308 25327 4310 25347
rect 4332 25327 4334 25347
rect 4404 25327 4406 25347
rect 4500 25327 4502 25347
rect 4596 25327 4598 25347
rect 4692 25327 4694 25347
rect 4860 25327 4862 25347
rect 4956 25327 4958 25347
rect 4980 25327 4982 25347
rect 5052 25327 5054 25347
rect 5124 25327 5126 25347
rect 5220 25327 5222 25347
rect 5268 25327 5270 25347
rect 5388 25327 5390 25347
rect 5484 25327 5486 25347
rect 5508 25327 5510 25347
rect 5532 25327 5534 25347
rect 5628 25327 5630 25347
rect 5652 25327 5654 25347
rect 5748 25327 5750 25347
rect 5796 25327 5798 25347
rect 5809 25327 5843 25328
rect 5844 25327 5846 25347
rect 5892 25327 5894 25347
rect 6132 25327 6134 25347
rect 6228 25327 6230 25347
rect 6252 25327 6254 25347
rect 6276 25327 6278 25347
rect 6324 25327 6326 25347
rect 6372 25327 6374 25347
rect 6420 25327 6422 25347
rect 6492 25327 6494 25347
rect 6516 25327 6518 25347
rect 6588 25327 6590 25347
rect 6612 25327 6614 25347
rect 6660 25327 6662 25347
rect 6684 25327 6686 25347
rect 6708 25327 6710 25347
rect 6780 25327 6782 25347
rect 6804 25327 6806 25347
rect 6900 25327 6902 25347
rect 6924 25327 6926 25347
rect 7020 25327 7022 25347
rect 7023 25344 7037 25347
rect 7047 25347 18149 25351
rect 7047 25344 7061 25347
rect 7068 25344 7071 25347
rect 7164 25327 7166 25347
rect 7236 25327 7238 25347
rect 7332 25327 7334 25347
rect 7380 25327 7382 25347
rect 7428 25327 7430 25347
rect 7452 25327 7454 25347
rect 7476 25327 7478 25347
rect 7524 25327 7526 25347
rect 7548 25327 7550 25347
rect 7572 25327 7574 25347
rect 7620 25327 7622 25347
rect 7644 25327 7646 25347
rect 7668 25327 7670 25347
rect 7897 25342 7900 25347
rect 7907 25328 7910 25342
rect 7908 25327 7910 25328
rect 7956 25327 7958 25347
rect 8028 25344 8030 25347
rect 8028 25327 8031 25344
rect 8124 25327 8126 25347
rect 8268 25327 8270 25347
rect 8340 25327 8342 25347
rect 8364 25327 8366 25347
rect 8436 25327 8438 25347
rect 8652 25327 8654 25347
rect 8700 25327 8702 25347
rect 8748 25327 8750 25347
rect 8820 25327 8822 25347
rect 8844 25327 8846 25347
rect 8868 25327 8870 25347
rect 9516 25327 9518 25347
rect 9660 25327 9662 25347
rect 9684 25327 9686 25347
rect 9756 25327 9758 25347
rect 9780 25327 9782 25347
rect 9804 25327 9806 25347
rect 9852 25327 9854 25347
rect 9900 25327 9902 25347
rect 9948 25327 9950 25347
rect 10044 25327 10046 25347
rect 10116 25327 10118 25347
rect 10188 25327 10190 25347
rect 10212 25327 10214 25347
rect 10284 25327 10286 25347
rect 10332 25327 10334 25347
rect 10380 25327 10382 25347
rect 10428 25327 10430 25347
rect 10476 25327 10478 25347
rect 10500 25327 10502 25347
rect 10524 25327 10526 25347
rect 10572 25327 10574 25347
rect 10596 25327 10598 25347
rect 10620 25327 10622 25347
rect 10692 25327 10694 25347
rect 10716 25327 10718 25347
rect 10788 25327 10790 25347
rect 10956 25327 10958 25347
rect 11004 25327 11006 25347
rect 11052 25327 11054 25347
rect 11100 25327 11102 25347
rect 11172 25327 11174 25347
rect 11220 25327 11222 25347
rect 11340 25327 11342 25347
rect 11436 25327 11438 25347
rect 11532 25327 11534 25347
rect 11580 25327 11582 25347
rect 11628 25327 11630 25347
rect 11676 25327 11678 25347
rect 11724 25327 11726 25347
rect 11772 25327 11774 25347
rect 11796 25327 11798 25347
rect 11892 25327 11894 25347
rect 11988 25327 11990 25347
rect 12060 25327 12062 25347
rect 12132 25327 12134 25347
rect 12228 25327 12230 25347
rect 12276 25327 12278 25347
rect 12324 25327 12326 25347
rect 12420 25327 12422 25347
rect 12444 25327 12446 25347
rect 12492 25327 12494 25347
rect 12516 25327 12518 25347
rect 12540 25327 12542 25347
rect 12588 25327 12590 25347
rect 12636 25327 12638 25347
rect 12732 25327 12734 25347
rect 12756 25327 12758 25347
rect 12804 25327 12806 25347
rect 12828 25327 12830 25347
rect 12927 25344 12941 25347
rect 12948 25344 12951 25347
rect 12972 25327 12974 25347
rect 13044 25327 13046 25347
rect 13068 25327 13070 25347
rect 13116 25327 13118 25347
rect 13284 25327 13286 25347
rect 13332 25327 13334 25347
rect 13572 25327 13574 25347
rect 13620 25327 13622 25347
rect 13668 25327 13670 25347
rect 13716 25327 13718 25347
rect 13764 25327 13766 25347
rect 13860 25327 13862 25347
rect 13956 25327 13958 25347
rect 14004 25327 14006 25347
rect 14100 25327 14102 25347
rect 15180 25327 15182 25347
rect 15231 25344 15245 25347
rect 15276 25327 15278 25347
rect 15420 25327 15422 25347
rect 15492 25327 15494 25347
rect 15660 25327 15662 25347
rect 15708 25327 15710 25347
rect 15732 25327 15734 25347
rect 15756 25327 15758 25347
rect 15804 25327 15806 25347
rect 15828 25327 15830 25347
rect 15852 25327 15854 25347
rect 15900 25327 15902 25347
rect 15948 25327 15950 25347
rect 16009 25327 16043 25328
rect 16044 25327 16046 25347
rect 16068 25327 16070 25347
rect 16164 25327 16166 25347
rect 16260 25327 16262 25347
rect 16308 25328 16310 25347
rect 16273 25327 16331 25328
rect 16332 25327 16334 25347
rect 16404 25327 16406 25347
rect 16431 25344 16445 25347
rect 16452 25344 16455 25347
rect 16548 25327 16550 25347
rect 16572 25327 16574 25347
rect 16620 25327 16622 25347
rect 16668 25327 16670 25347
rect 16716 25327 16718 25347
rect 16764 25327 16766 25347
rect 16812 25327 16814 25347
rect 16884 25327 16886 25347
rect 16908 25327 16910 25347
rect 16980 25327 16982 25347
rect 17148 25327 17150 25347
rect 17196 25327 17198 25347
rect 17220 25327 17222 25347
rect 17292 25327 17294 25347
rect 17316 25327 17318 25347
rect 18132 25327 18134 25347
rect 18135 25344 18149 25347
rect 18159 25347 23789 25351
rect 18159 25344 18173 25347
rect 18228 25327 18230 25347
rect 18289 25327 18323 25328
rect 18396 25327 18398 25347
rect 18492 25327 18494 25347
rect 18516 25327 18518 25347
rect 18564 25327 18566 25347
rect 18612 25327 18614 25347
rect 18660 25327 18662 25347
rect 18756 25327 18758 25347
rect 18900 25327 18902 25347
rect 18924 25327 18926 25347
rect 18996 25327 18998 25347
rect 19020 25327 19022 25347
rect 19092 25327 19094 25347
rect 19116 25327 19118 25347
rect 19140 25327 19142 25347
rect 19188 25327 19190 25347
rect 19236 25327 19238 25347
rect 19332 25327 19334 25347
rect 19788 25327 19790 25347
rect 19836 25327 19838 25347
rect 19860 25327 19862 25347
rect 19884 25327 19886 25347
rect 19932 25327 19934 25347
rect 19956 25327 19958 25347
rect 19980 25327 19982 25347
rect 20028 25327 20030 25347
rect 20052 25327 20054 25347
rect 20076 25327 20078 25347
rect 20148 25327 20150 25347
rect 20172 25327 20174 25347
rect 20196 25327 20198 25347
rect 20268 25327 20270 25347
rect 20292 25327 20294 25347
rect 20388 25327 20390 25347
rect 20412 25327 20414 25347
rect 20508 25327 20510 25347
rect 20604 25327 20606 25347
rect 20964 25327 20966 25347
rect 21012 25327 21014 25347
rect 21108 25327 21110 25347
rect 21204 25327 21206 25347
rect 21300 25327 21302 25347
rect 21324 25327 21326 25347
rect 21444 25327 21446 25347
rect 21468 25327 21470 25347
rect 21564 25327 21566 25347
rect 21588 25327 21590 25347
rect 21684 25327 21686 25347
rect 21708 25327 21710 25347
rect 21828 25327 21830 25347
rect 21924 25327 21926 25347
rect 22068 25327 22070 25347
rect 22188 25327 22190 25347
rect 22212 25327 22214 25347
rect 22884 25327 22886 25347
rect 22980 25327 22982 25347
rect 23076 25327 23078 25347
rect 23100 25327 23102 25347
rect 23124 25327 23126 25347
rect 23244 25327 23246 25347
rect 23340 25327 23342 25347
rect 23412 25327 23414 25347
rect 23460 25327 23462 25347
rect 23508 25327 23510 25347
rect 23556 25327 23558 25347
rect 23604 25327 23606 25347
rect 23652 25327 23654 25347
rect 23676 25327 23678 25347
rect 23700 25327 23702 25347
rect 23772 25327 23774 25347
rect 23775 25344 23789 25347
rect 23796 25347 24995 25351
rect 25057 25351 25091 25352
rect 25153 25351 25211 25352
rect 25249 25351 25283 25352
rect 25057 25347 25283 25351
rect 23796 25344 23813 25347
rect 23820 25344 23823 25347
rect 23796 25327 23798 25344
rect 23916 25327 23918 25347
rect 24012 25327 24014 25347
rect 24060 25327 24062 25347
rect 24156 25327 24158 25347
rect 24492 25327 24494 25347
rect 24516 25327 24518 25347
rect 24588 25327 24590 25347
rect 24612 25327 24614 25347
rect 24625 25327 24659 25328
rect 24684 25327 24686 25347
rect 24732 25327 24734 25347
rect 24756 25327 24758 25347
rect 24780 25327 24782 25347
rect 24852 25327 24854 25347
rect 24876 25327 24878 25347
rect 24961 25342 24964 25347
rect 24972 25342 24974 25347
rect 25057 25342 25060 25347
rect 25068 25344 25070 25347
rect 25068 25342 25071 25344
rect 25153 25342 25156 25347
rect 25164 25344 25166 25347
rect 25164 25342 25167 25344
rect 25249 25342 25252 25347
rect 25260 25344 25262 25347
rect 25260 25342 25263 25344
rect 24971 25328 24974 25342
rect 25067 25328 25071 25342
rect 25163 25328 25167 25342
rect 25259 25334 25263 25342
rect 25273 25334 25277 25342
rect 25259 25328 25273 25334
rect 24889 25327 24923 25328
rect -14471 25323 -12643 25327
rect -14471 25320 -14467 25323
rect -14460 25320 -14457 25323
rect -14351 25303 -14317 25304
rect -14100 25303 -14098 25323
rect -14004 25303 -14002 25323
rect -13788 25303 -13786 25323
rect -13428 25303 -13426 25323
rect -12756 25303 -12754 25323
rect -12657 25320 -12643 25323
rect -12636 25323 -9451 25327
rect -12636 25320 -12619 25323
rect -12636 25303 -12634 25320
rect -12348 25303 -12346 25323
rect -12252 25303 -12250 25323
rect -12156 25303 -12154 25323
rect -12060 25303 -12058 25323
rect -11772 25303 -11770 25323
rect -11676 25303 -11674 25323
rect -11508 25303 -11506 25323
rect -11436 25303 -11434 25323
rect -11412 25303 -11410 25323
rect -11340 25303 -11338 25323
rect -11196 25303 -11194 25323
rect -11100 25303 -11098 25323
rect -10764 25303 -10762 25323
rect -10644 25303 -10642 25323
rect -9996 25303 -9994 25323
rect -9900 25303 -9898 25323
rect -9732 25303 -9730 25323
rect -9465 25320 -9451 25323
rect -9444 25323 -9115 25327
rect -9444 25320 -9427 25323
rect -9444 25303 -9442 25320
rect -9348 25303 -9346 25323
rect -9228 25303 -9226 25323
rect -9129 25320 -9115 25323
rect -9108 25323 -3451 25327
rect -9108 25320 -9091 25323
rect -9108 25303 -9106 25320
rect -8436 25303 -8434 25323
rect -8364 25303 -8362 25323
rect -8340 25303 -8338 25323
rect -8268 25303 -8266 25323
rect -8004 25303 -8002 25323
rect -7932 25303 -7930 25323
rect -7727 25303 -7693 25304
rect -7620 25303 -7618 25323
rect -7524 25303 -7522 25323
rect -7356 25303 -7354 25323
rect -7308 25303 -7306 25323
rect -7212 25303 -7210 25323
rect -7044 25303 -7042 25323
rect -6948 25303 -6946 25323
rect -6852 25303 -6850 25323
rect -6756 25303 -6754 25323
rect -6660 25303 -6658 25323
rect -6612 25303 -6610 25323
rect -6516 25303 -6514 25323
rect -6372 25303 -6370 25323
rect -6036 25303 -6034 25323
rect -5892 25303 -5890 25323
rect -5196 25303 -5194 25323
rect -5100 25303 -5098 25323
rect -4716 25303 -4714 25323
rect -4500 25303 -4498 25323
rect -4404 25303 -4402 25323
rect -4308 25303 -4306 25323
rect -4164 25303 -4162 25323
rect -4020 25303 -4018 25323
rect -3876 25303 -3874 25323
rect -3732 25303 -3730 25323
rect -3636 25303 -3634 25323
rect -3540 25303 -3538 25323
rect -3468 25303 -3466 25323
rect -3465 25320 -3451 25323
rect -3441 25323 7997 25327
rect -3441 25320 -3427 25323
rect -3420 25320 -3417 25323
rect -3324 25303 -3322 25323
rect -3228 25304 -3226 25323
rect -3239 25303 -3205 25304
rect -3132 25303 -3130 25323
rect -3108 25303 -3106 25323
rect -3012 25303 -3010 25323
rect -2964 25303 -2962 25323
rect -2916 25303 -2914 25323
rect -2892 25303 -2890 25323
rect -2868 25303 -2866 25323
rect -2820 25303 -2818 25323
rect -2796 25303 -2794 25323
rect -2772 25303 -2770 25323
rect -2676 25303 -2674 25323
rect -2580 25303 -2578 25323
rect -2364 25303 -2362 25323
rect -2316 25303 -2314 25323
rect -2268 25303 -2266 25323
rect -2244 25303 -2242 25323
rect -2172 25303 -2170 25323
rect -2148 25303 -2146 25323
rect -2076 25303 -2074 25323
rect -2052 25303 -2050 25323
rect -1980 25303 -1978 25323
rect -1884 25303 -1882 25323
rect -1572 25303 -1570 25323
rect -1476 25303 -1474 25323
rect -1391 25318 -1388 25323
rect -1380 25318 -1378 25323
rect -1381 25304 -1378 25318
rect -1356 25303 -1354 25323
rect -1260 25303 -1258 25323
rect -1236 25303 -1234 25323
rect -1140 25303 -1138 25323
rect -983 25303 -925 25304
rect -708 25303 -706 25323
rect -660 25303 -658 25323
rect -612 25303 -610 25323
rect -492 25303 -490 25323
rect -444 25303 -442 25323
rect -396 25303 -394 25323
rect -348 25303 -346 25323
rect -300 25303 -298 25323
rect -276 25303 -274 25323
rect -12 25303 -10 25323
rect 156 25303 158 25323
rect 204 25303 206 25323
rect 252 25303 254 25323
rect 348 25303 350 25323
rect 468 25303 470 25323
rect 492 25303 494 25323
rect 564 25303 566 25323
rect 588 25303 590 25323
rect 636 25303 638 25323
rect 660 25303 662 25323
rect 732 25303 734 25323
rect 1092 25303 1094 25323
rect 1140 25303 1142 25323
rect 1236 25303 1238 25323
rect 1308 25303 1310 25323
rect 1332 25303 1334 25323
rect 1380 25303 1382 25323
rect 1428 25303 1430 25323
rect 1476 25303 1478 25323
rect 1692 25303 1694 25323
rect 1788 25303 1790 25323
rect 2028 25303 2030 25323
rect 2076 25303 2078 25323
rect 2100 25303 2102 25323
rect 2124 25303 2126 25323
rect 2244 25303 2246 25323
rect 2412 25303 2414 25323
rect 2460 25303 2462 25323
rect 2508 25303 2510 25323
rect 2569 25318 2572 25323
rect 2580 25318 2582 25323
rect 2579 25304 2582 25318
rect 2604 25303 2606 25323
rect 2676 25320 2678 25323
rect 2676 25303 2679 25320
rect 2772 25303 2774 25323
rect 2868 25303 2870 25323
rect 2940 25303 2942 25323
rect 3012 25303 3014 25323
rect 3108 25303 3110 25323
rect 3348 25303 3350 25323
rect 3396 25303 3398 25323
rect 3564 25303 3566 25323
rect 3636 25303 3638 25323
rect 3660 25303 3662 25323
rect 3732 25303 3734 25323
rect 3780 25303 3782 25323
rect 3828 25303 3830 25323
rect 3924 25303 3926 25323
rect 3937 25303 3971 25304
rect 4020 25303 4022 25323
rect 4044 25304 4046 25323
rect 4033 25303 4067 25304
rect 4092 25303 4094 25323
rect 4140 25304 4142 25323
rect 4129 25303 4163 25304
rect 4188 25303 4190 25323
rect 4236 25304 4238 25323
rect 4225 25303 4259 25304
rect 4308 25303 4310 25323
rect 4332 25304 4334 25323
rect 4321 25303 4355 25304
rect 4404 25303 4406 25323
rect 4500 25303 4502 25323
rect 4596 25303 4598 25323
rect 4692 25303 4694 25323
rect 4860 25303 4862 25323
rect 4956 25303 4958 25323
rect 4980 25303 4982 25323
rect 5052 25303 5054 25323
rect 5124 25303 5126 25323
rect 5220 25303 5222 25323
rect 5268 25303 5270 25323
rect 5388 25303 5390 25323
rect 5484 25303 5486 25323
rect 5508 25303 5510 25323
rect 5532 25303 5534 25323
rect 5628 25303 5630 25323
rect 5652 25303 5654 25323
rect 5748 25303 5750 25323
rect 5796 25303 5798 25323
rect 5844 25303 5846 25323
rect 5892 25303 5894 25323
rect 6132 25303 6134 25323
rect 6228 25303 6230 25323
rect 6252 25303 6254 25323
rect 6276 25303 6278 25323
rect 6324 25303 6326 25323
rect 6372 25303 6374 25323
rect 6420 25303 6422 25323
rect 6492 25303 6494 25323
rect 6516 25303 6518 25323
rect 6588 25303 6590 25323
rect 6612 25303 6614 25323
rect 6660 25303 6662 25323
rect 6684 25303 6686 25323
rect 6708 25303 6710 25323
rect 6780 25303 6782 25323
rect 6804 25303 6806 25323
rect 6900 25303 6902 25323
rect 6924 25303 6926 25323
rect 7020 25303 7022 25323
rect 7164 25303 7166 25323
rect 7236 25303 7238 25323
rect 7332 25303 7334 25323
rect 7380 25303 7382 25323
rect 7428 25303 7430 25323
rect 7452 25303 7454 25323
rect 7476 25303 7478 25323
rect 7524 25303 7526 25323
rect 7548 25303 7550 25323
rect 7572 25303 7574 25323
rect 7620 25303 7622 25323
rect 7644 25303 7646 25323
rect 7668 25303 7670 25323
rect 7908 25303 7910 25323
rect 7956 25303 7958 25323
rect 7983 25320 7997 25323
rect 8007 25323 24923 25327
rect 8007 25320 8021 25323
rect 8028 25320 8031 25323
rect 8124 25303 8126 25323
rect 8268 25303 8270 25323
rect 8340 25303 8342 25323
rect 8364 25303 8366 25323
rect 8436 25304 8438 25323
rect 8401 25303 8459 25304
rect 8652 25303 8654 25323
rect 8700 25303 8702 25323
rect 8748 25303 8750 25323
rect 8820 25303 8822 25323
rect 8844 25303 8846 25323
rect 8868 25303 8870 25323
rect 9516 25303 9518 25323
rect 9660 25303 9662 25323
rect 9684 25303 9686 25323
rect 9756 25303 9758 25323
rect 9780 25303 9782 25323
rect 9804 25303 9806 25323
rect 9852 25303 9854 25323
rect 9900 25303 9902 25323
rect 9948 25303 9950 25323
rect 10044 25303 10046 25323
rect 10116 25303 10118 25323
rect 10188 25303 10190 25323
rect 10212 25303 10214 25323
rect 10284 25303 10286 25323
rect 10332 25303 10334 25323
rect 10380 25303 10382 25323
rect 10428 25303 10430 25323
rect 10476 25303 10478 25323
rect 10500 25303 10502 25323
rect 10524 25303 10526 25323
rect 10572 25303 10574 25323
rect 10596 25303 10598 25323
rect 10620 25303 10622 25323
rect 10692 25303 10694 25323
rect 10716 25303 10718 25323
rect 10788 25303 10790 25323
rect 10956 25303 10958 25323
rect 11004 25303 11006 25323
rect 11052 25303 11054 25323
rect 11100 25303 11102 25323
rect 11172 25303 11174 25323
rect 11220 25303 11222 25323
rect 11340 25303 11342 25323
rect 11436 25303 11438 25323
rect 11532 25303 11534 25323
rect 11580 25303 11582 25323
rect 11628 25303 11630 25323
rect 11676 25303 11678 25323
rect 11724 25303 11726 25323
rect 11772 25303 11774 25323
rect 11796 25303 11798 25323
rect 11892 25303 11894 25323
rect 11988 25303 11990 25323
rect 12060 25303 12062 25323
rect 12132 25303 12134 25323
rect 12228 25303 12230 25323
rect 12276 25303 12278 25323
rect 12324 25303 12326 25323
rect 12420 25303 12422 25323
rect 12444 25303 12446 25323
rect 12492 25303 12494 25323
rect 12516 25303 12518 25323
rect 12540 25303 12542 25323
rect 12588 25303 12590 25323
rect 12636 25303 12638 25323
rect 12732 25303 12734 25323
rect 12756 25303 12758 25323
rect 12804 25303 12806 25323
rect 12828 25303 12830 25323
rect 12972 25303 12974 25323
rect 13044 25303 13046 25323
rect 13068 25303 13070 25323
rect 13116 25303 13118 25323
rect 13284 25303 13286 25323
rect 13332 25303 13334 25323
rect 13572 25303 13574 25323
rect 13620 25303 13622 25323
rect 13668 25303 13670 25323
rect 13716 25303 13718 25323
rect 13764 25303 13766 25323
rect 13860 25303 13862 25323
rect 13956 25303 13958 25323
rect 14004 25303 14006 25323
rect 14100 25303 14102 25323
rect 15180 25303 15182 25323
rect 15276 25303 15278 25323
rect 15420 25303 15422 25323
rect 15492 25303 15494 25323
rect 15660 25303 15662 25323
rect 15708 25303 15710 25323
rect 15732 25303 15734 25323
rect 15756 25303 15758 25323
rect 15804 25303 15806 25323
rect 15828 25303 15830 25323
rect 15852 25303 15854 25323
rect 15900 25303 15902 25323
rect 15948 25303 15950 25323
rect 16044 25303 16046 25323
rect 16068 25303 16070 25323
rect 16164 25303 16166 25323
rect 16260 25303 16262 25323
rect 16297 25318 16300 25323
rect 16308 25318 16310 25323
rect 16307 25304 16310 25318
rect 16332 25303 16334 25323
rect 16404 25320 16406 25323
rect 16404 25303 16407 25320
rect 16548 25303 16550 25323
rect 16572 25303 16574 25323
rect 16620 25303 16622 25323
rect 16668 25303 16670 25323
rect 16716 25303 16718 25323
rect 16764 25303 16766 25323
rect 16812 25303 16814 25323
rect 16884 25303 16886 25323
rect 16908 25303 16910 25323
rect 16980 25303 16982 25323
rect 17148 25303 17150 25323
rect 17196 25303 17198 25323
rect 17220 25303 17222 25323
rect 17292 25303 17294 25323
rect 17316 25303 17318 25323
rect 18132 25303 18134 25323
rect 18228 25303 18230 25323
rect 18396 25320 18398 25323
rect 18396 25303 18399 25320
rect 18492 25303 18494 25323
rect 18516 25303 18518 25323
rect 18564 25303 18566 25323
rect 18612 25303 18614 25323
rect 18660 25303 18662 25323
rect 18756 25303 18758 25323
rect 18900 25303 18902 25323
rect 18924 25303 18926 25323
rect 18996 25303 18998 25323
rect 19020 25303 19022 25323
rect 19092 25303 19094 25323
rect 19116 25303 19118 25323
rect 19140 25303 19142 25323
rect 19188 25303 19190 25323
rect 19236 25303 19238 25323
rect 19332 25304 19334 25323
rect 19297 25303 19355 25304
rect 19788 25303 19790 25323
rect 19836 25303 19838 25323
rect 19860 25303 19862 25323
rect 19884 25303 19886 25323
rect 19932 25303 19934 25323
rect 19956 25303 19958 25323
rect 19980 25303 19982 25323
rect 20028 25303 20030 25323
rect 20052 25303 20054 25323
rect 20076 25303 20078 25323
rect 20148 25303 20150 25323
rect 20172 25303 20174 25323
rect 20196 25303 20198 25323
rect 20268 25303 20270 25323
rect 20292 25303 20294 25323
rect 20388 25303 20390 25323
rect 20412 25303 20414 25323
rect 20508 25303 20510 25323
rect 20604 25303 20606 25323
rect 20964 25303 20966 25323
rect 21012 25303 21014 25323
rect 21108 25303 21110 25323
rect 21204 25303 21206 25323
rect 21300 25303 21302 25323
rect 21324 25303 21326 25323
rect 21444 25303 21446 25323
rect 21468 25303 21470 25323
rect 21564 25303 21566 25323
rect 21588 25303 21590 25323
rect 21684 25303 21686 25323
rect 21708 25303 21710 25323
rect 21828 25303 21830 25323
rect 21924 25303 21926 25323
rect 22068 25303 22070 25323
rect 22188 25303 22190 25323
rect 22212 25303 22214 25323
rect 22884 25303 22886 25323
rect 22980 25303 22982 25323
rect 23076 25303 23078 25323
rect 23100 25303 23102 25323
rect 23124 25303 23126 25323
rect 23244 25303 23246 25323
rect 23340 25303 23342 25323
rect 23412 25303 23414 25323
rect 23460 25303 23462 25323
rect 23508 25303 23510 25323
rect 23556 25303 23558 25323
rect 23604 25303 23606 25323
rect 23652 25303 23654 25323
rect 23676 25303 23678 25323
rect 23700 25303 23702 25323
rect 23772 25303 23774 25323
rect 23796 25303 23798 25323
rect 23916 25303 23918 25323
rect 24012 25303 24014 25323
rect 24060 25303 24062 25323
rect 24156 25303 24158 25323
rect 24492 25303 24494 25323
rect 24516 25303 24518 25323
rect 24588 25303 24590 25323
rect 24612 25303 24614 25323
rect 24684 25303 24686 25323
rect 24732 25320 24734 25323
rect 24732 25303 24735 25320
rect 24756 25303 24758 25323
rect 24780 25303 24782 25323
rect 24852 25303 24854 25323
rect 24876 25304 24878 25323
rect 24865 25303 24899 25304
rect -14351 25299 16373 25303
rect -14207 25279 -14173 25280
rect -14100 25279 -14098 25299
rect -14004 25279 -14002 25299
rect -13788 25279 -13786 25299
rect -13641 25296 -13627 25299
rect -13428 25279 -13426 25299
rect -12959 25279 -12901 25280
rect -12756 25279 -12754 25299
rect -12636 25279 -12634 25299
rect -12348 25279 -12346 25299
rect -12252 25279 -12250 25299
rect -12156 25279 -12154 25299
rect -12060 25279 -12058 25299
rect -11772 25279 -11770 25299
rect -11676 25279 -11674 25299
rect -11508 25279 -11506 25299
rect -11436 25279 -11434 25299
rect -11412 25279 -11410 25299
rect -11340 25279 -11338 25299
rect -11196 25279 -11194 25299
rect -11100 25279 -11098 25299
rect -10764 25279 -10762 25299
rect -10644 25279 -10642 25299
rect -9996 25279 -9994 25299
rect -9900 25279 -9898 25299
rect -9732 25279 -9730 25299
rect -9695 25279 -9661 25280
rect -9444 25279 -9442 25299
rect -9348 25279 -9346 25299
rect -9228 25279 -9226 25299
rect -9108 25279 -9106 25299
rect -8591 25279 -8557 25280
rect -8436 25279 -8434 25299
rect -8399 25279 -8365 25280
rect -8364 25279 -8362 25299
rect -8340 25279 -8338 25299
rect -8268 25279 -8266 25299
rect -8004 25279 -8002 25299
rect -7932 25279 -7930 25299
rect -7620 25296 -7618 25299
rect -7620 25279 -7617 25296
rect -7524 25279 -7522 25299
rect -7356 25279 -7354 25299
rect -7308 25279 -7306 25299
rect -7212 25279 -7210 25299
rect -7044 25279 -7042 25299
rect -6948 25279 -6946 25299
rect -6852 25279 -6850 25299
rect -6756 25279 -6754 25299
rect -6660 25279 -6658 25299
rect -6612 25279 -6610 25299
rect -6516 25279 -6514 25299
rect -6372 25279 -6370 25299
rect -6036 25279 -6034 25299
rect -5892 25279 -5890 25299
rect -5196 25279 -5194 25299
rect -5100 25279 -5098 25299
rect -4716 25279 -4714 25299
rect -4500 25279 -4498 25299
rect -4404 25279 -4402 25299
rect -4308 25279 -4306 25299
rect -4164 25279 -4162 25299
rect -4020 25279 -4018 25299
rect -3876 25279 -3874 25299
rect -3732 25279 -3730 25299
rect -3636 25279 -3634 25299
rect -3540 25279 -3538 25299
rect -3468 25279 -3466 25299
rect -3324 25279 -3322 25299
rect -3239 25294 -3236 25299
rect -3228 25294 -3226 25299
rect -3229 25280 -3226 25294
rect -3132 25296 -3130 25299
rect -3132 25279 -3129 25296
rect -3108 25279 -3106 25299
rect -3012 25279 -3010 25299
rect -2964 25279 -2962 25299
rect -2916 25279 -2914 25299
rect -2892 25279 -2890 25299
rect -2868 25279 -2866 25299
rect -2820 25279 -2818 25299
rect -2796 25279 -2794 25299
rect -2772 25279 -2770 25299
rect -2676 25279 -2674 25299
rect -2580 25279 -2578 25299
rect -2364 25279 -2362 25299
rect -2316 25279 -2314 25299
rect -2268 25279 -2266 25299
rect -2244 25279 -2242 25299
rect -2172 25279 -2170 25299
rect -2148 25279 -2146 25299
rect -2076 25279 -2074 25299
rect -2052 25279 -2050 25299
rect -1980 25279 -1978 25299
rect -1884 25279 -1882 25299
rect -1572 25279 -1570 25299
rect -1476 25279 -1474 25299
rect -1356 25279 -1354 25299
rect -1305 25296 -1291 25299
rect -1260 25279 -1258 25299
rect -1236 25279 -1234 25299
rect -1140 25279 -1138 25299
rect -876 25279 -873 25296
rect -708 25279 -706 25299
rect -660 25279 -658 25299
rect -612 25279 -610 25299
rect -492 25279 -490 25299
rect -444 25279 -442 25299
rect -396 25279 -394 25299
rect -348 25279 -346 25299
rect -300 25279 -298 25299
rect -276 25279 -274 25299
rect -12 25279 -10 25299
rect 156 25279 158 25299
rect 204 25279 206 25299
rect 252 25279 254 25299
rect 348 25279 350 25299
rect 468 25279 470 25299
rect 492 25279 494 25299
rect 564 25279 566 25299
rect 588 25279 590 25299
rect 636 25279 638 25299
rect 660 25279 662 25299
rect 732 25279 734 25299
rect 1092 25279 1094 25299
rect 1140 25279 1142 25299
rect 1236 25279 1238 25299
rect 1308 25279 1310 25299
rect 1332 25279 1334 25299
rect 1380 25279 1382 25299
rect 1428 25279 1430 25299
rect 1476 25279 1478 25299
rect 1692 25279 1694 25299
rect 1788 25279 1790 25299
rect 2028 25279 2030 25299
rect 2076 25279 2078 25299
rect 2100 25279 2102 25299
rect 2124 25279 2126 25299
rect 2244 25279 2246 25299
rect 2412 25279 2414 25299
rect 2460 25279 2462 25299
rect 2508 25279 2510 25299
rect 2604 25279 2606 25299
rect 2655 25296 2669 25299
rect 2676 25296 2679 25299
rect 2772 25279 2774 25299
rect 2868 25279 2870 25299
rect 2940 25279 2942 25299
rect 3012 25279 3014 25299
rect 3108 25279 3110 25299
rect 3348 25280 3350 25299
rect 3313 25279 3371 25280
rect 3396 25279 3398 25299
rect 3564 25279 3566 25299
rect 3636 25279 3638 25299
rect 3660 25279 3662 25299
rect 3732 25279 3734 25299
rect 3780 25279 3782 25299
rect 3828 25279 3830 25299
rect 3924 25279 3926 25299
rect 4020 25279 4022 25299
rect 4033 25294 4036 25299
rect 4044 25296 4046 25299
rect 4044 25294 4047 25296
rect 4043 25280 4047 25294
rect 4092 25279 4094 25299
rect 4129 25294 4132 25299
rect 4140 25296 4142 25299
rect 4140 25294 4143 25296
rect 4139 25280 4143 25294
rect 4188 25279 4190 25299
rect 4225 25294 4228 25299
rect 4236 25296 4238 25299
rect 4236 25294 4239 25296
rect 4235 25280 4239 25294
rect 4308 25279 4310 25299
rect 4321 25294 4324 25299
rect 4332 25296 4334 25299
rect 4332 25294 4335 25296
rect 4331 25280 4335 25294
rect 4404 25279 4406 25299
rect 4500 25279 4502 25299
rect 4596 25279 4598 25299
rect 4692 25279 4694 25299
rect 4860 25279 4862 25299
rect 4956 25279 4958 25299
rect 4980 25279 4982 25299
rect 5052 25279 5054 25299
rect 5124 25279 5126 25299
rect 5220 25279 5222 25299
rect 5268 25279 5270 25299
rect 5388 25279 5390 25299
rect 5484 25279 5486 25299
rect 5508 25279 5510 25299
rect 5532 25279 5534 25299
rect 5628 25279 5630 25299
rect 5652 25279 5654 25299
rect 5748 25279 5750 25299
rect 5796 25279 5798 25299
rect 5844 25279 5846 25299
rect 5892 25279 5894 25299
rect 5895 25296 5909 25299
rect 6132 25279 6134 25299
rect 6228 25279 6230 25299
rect 6252 25279 6254 25299
rect 6276 25279 6278 25299
rect 6324 25279 6326 25299
rect 6372 25279 6374 25299
rect 6420 25279 6422 25299
rect 6492 25279 6494 25299
rect 6516 25279 6518 25299
rect 6588 25279 6590 25299
rect 6612 25279 6614 25299
rect 6660 25279 6662 25299
rect 6684 25279 6686 25299
rect 6708 25279 6710 25299
rect 6780 25279 6782 25299
rect 6804 25279 6806 25299
rect 6900 25279 6902 25299
rect 6924 25279 6926 25299
rect 7020 25279 7022 25299
rect 7164 25279 7166 25299
rect 7236 25279 7238 25299
rect 7332 25279 7334 25299
rect 7380 25279 7382 25299
rect 7428 25279 7430 25299
rect 7452 25279 7454 25299
rect 7476 25279 7478 25299
rect 7524 25279 7526 25299
rect 7548 25279 7550 25299
rect 7572 25279 7574 25299
rect 7620 25279 7622 25299
rect 7644 25279 7646 25299
rect 7668 25279 7670 25299
rect 7908 25279 7910 25299
rect 7956 25279 7958 25299
rect 8124 25279 8126 25299
rect 8268 25279 8270 25299
rect 8340 25279 8342 25299
rect 8364 25279 8366 25299
rect 8425 25294 8428 25299
rect 8436 25294 8438 25299
rect 8435 25280 8438 25294
rect 8652 25279 8654 25299
rect 8700 25279 8702 25299
rect 8748 25279 8750 25299
rect 8820 25279 8822 25299
rect 8844 25279 8846 25299
rect 8868 25279 8870 25299
rect 9516 25279 9518 25299
rect 9660 25279 9662 25299
rect 9684 25279 9686 25299
rect 9756 25279 9758 25299
rect 9780 25279 9782 25299
rect 9804 25279 9806 25299
rect 9852 25279 9854 25299
rect 9900 25279 9902 25299
rect 9948 25279 9950 25299
rect 10044 25279 10046 25299
rect 10116 25279 10118 25299
rect 10188 25279 10190 25299
rect 10212 25279 10214 25299
rect 10284 25279 10286 25299
rect 10332 25279 10334 25299
rect 10380 25279 10382 25299
rect 10428 25279 10430 25299
rect 10476 25279 10478 25299
rect 10500 25279 10502 25299
rect 10524 25279 10526 25299
rect 10572 25279 10574 25299
rect 10596 25279 10598 25299
rect 10620 25279 10622 25299
rect 10692 25279 10694 25299
rect 10716 25279 10718 25299
rect 10788 25279 10790 25299
rect 10956 25279 10958 25299
rect 11004 25279 11006 25299
rect 11052 25279 11054 25299
rect 11100 25279 11102 25299
rect 11172 25279 11174 25299
rect 11220 25279 11222 25299
rect 11340 25279 11342 25299
rect 11436 25279 11438 25299
rect 11532 25279 11534 25299
rect 11580 25279 11582 25299
rect 11628 25279 11630 25299
rect 11676 25279 11678 25299
rect 11724 25279 11726 25299
rect 11772 25279 11774 25299
rect 11796 25279 11798 25299
rect 11892 25279 11894 25299
rect 11988 25279 11990 25299
rect 12060 25279 12062 25299
rect 12132 25279 12134 25299
rect 12228 25279 12230 25299
rect 12276 25279 12278 25299
rect 12324 25279 12326 25299
rect 12420 25279 12422 25299
rect 12444 25279 12446 25299
rect 12492 25279 12494 25299
rect 12516 25279 12518 25299
rect 12540 25279 12542 25299
rect 12588 25279 12590 25299
rect 12636 25279 12638 25299
rect 12732 25279 12734 25299
rect 12756 25279 12758 25299
rect 12804 25279 12806 25299
rect 12828 25279 12830 25299
rect 12972 25279 12974 25299
rect 13044 25279 13046 25299
rect 13068 25279 13070 25299
rect 13116 25279 13118 25299
rect 13284 25279 13286 25299
rect 13332 25279 13334 25299
rect 13572 25279 13574 25299
rect 13620 25279 13622 25299
rect 13668 25279 13670 25299
rect 13716 25279 13718 25299
rect 13764 25279 13766 25299
rect 13860 25279 13862 25299
rect 13956 25279 13958 25299
rect 14004 25279 14006 25299
rect 14100 25279 14102 25299
rect 15180 25279 15182 25299
rect 15276 25279 15278 25299
rect 15420 25279 15422 25299
rect 15492 25279 15494 25299
rect 15660 25279 15662 25299
rect 15708 25279 15710 25299
rect 15732 25279 15734 25299
rect 15756 25279 15758 25299
rect 15804 25279 15806 25299
rect 15828 25279 15830 25299
rect 15852 25279 15854 25299
rect 15900 25279 15902 25299
rect 15948 25279 15950 25299
rect 16044 25279 16046 25299
rect 16068 25279 16070 25299
rect 16095 25296 16109 25299
rect 16164 25279 16166 25299
rect 16260 25279 16262 25299
rect 16332 25279 16334 25299
rect 16359 25296 16373 25299
rect 16383 25299 24899 25303
rect 16383 25296 16397 25299
rect 16404 25296 16407 25299
rect 16548 25279 16550 25299
rect 16572 25279 16574 25299
rect 16620 25279 16622 25299
rect 16668 25279 16670 25299
rect 16716 25279 16718 25299
rect 16764 25279 16766 25299
rect 16812 25279 16814 25299
rect 16884 25279 16886 25299
rect 16908 25279 16910 25299
rect 16980 25279 16982 25299
rect 17148 25279 17150 25299
rect 17196 25279 17198 25299
rect 17220 25279 17222 25299
rect 17292 25279 17294 25299
rect 17316 25279 17318 25299
rect 18132 25279 18134 25299
rect 18228 25279 18230 25299
rect 18375 25296 18389 25299
rect 18396 25296 18399 25299
rect 18492 25279 18494 25299
rect 18516 25279 18518 25299
rect 18564 25279 18566 25299
rect 18612 25279 18614 25299
rect 18660 25279 18662 25299
rect 18756 25279 18758 25299
rect 18900 25279 18902 25299
rect 18924 25279 18926 25299
rect 18996 25279 18998 25299
rect 19020 25279 19022 25299
rect 19092 25279 19094 25299
rect 19116 25279 19118 25299
rect 19140 25279 19142 25299
rect 19188 25279 19190 25299
rect 19236 25279 19238 25299
rect 19321 25294 19324 25299
rect 19332 25294 19334 25299
rect 19331 25280 19334 25294
rect 19788 25279 19790 25299
rect 19836 25279 19838 25299
rect 19860 25279 19862 25299
rect 19884 25279 19886 25299
rect 19932 25279 19934 25299
rect 19956 25279 19958 25299
rect 19980 25279 19982 25299
rect 20028 25279 20030 25299
rect 20052 25279 20054 25299
rect 20076 25279 20078 25299
rect 20148 25279 20150 25299
rect 20172 25279 20174 25299
rect 20196 25279 20198 25299
rect 20268 25279 20270 25299
rect 20292 25279 20294 25299
rect 20388 25279 20390 25299
rect 20412 25279 20414 25299
rect 20508 25279 20510 25299
rect 20604 25279 20606 25299
rect 20964 25279 20966 25299
rect 21012 25279 21014 25299
rect 21108 25279 21110 25299
rect 21204 25279 21206 25299
rect 21300 25279 21302 25299
rect 21324 25279 21326 25299
rect 21444 25279 21446 25299
rect 21468 25279 21470 25299
rect 21564 25279 21566 25299
rect 21588 25279 21590 25299
rect 21684 25279 21686 25299
rect 21708 25279 21710 25299
rect 21828 25279 21830 25299
rect 21924 25279 21926 25299
rect 22068 25279 22070 25299
rect 22188 25279 22190 25299
rect 22212 25279 22214 25299
rect 22884 25279 22886 25299
rect 22980 25279 22982 25299
rect 23076 25279 23078 25299
rect 23100 25279 23102 25299
rect 23124 25279 23126 25299
rect 23244 25279 23246 25299
rect 23340 25279 23342 25299
rect 23412 25279 23414 25299
rect 23460 25279 23462 25299
rect 23508 25279 23510 25299
rect 23556 25279 23558 25299
rect 23604 25279 23606 25299
rect 23652 25279 23654 25299
rect 23676 25279 23678 25299
rect 23700 25279 23702 25299
rect 23772 25279 23774 25299
rect 23796 25279 23798 25299
rect 23916 25279 23918 25299
rect 24012 25279 24014 25299
rect 24060 25279 24062 25299
rect 24156 25279 24158 25299
rect 24492 25279 24494 25299
rect 24516 25279 24518 25299
rect 24588 25279 24590 25299
rect 24612 25279 24614 25299
rect 24684 25279 24686 25299
rect 24711 25296 24725 25299
rect 24732 25296 24735 25299
rect 24756 25279 24758 25299
rect 24780 25279 24782 25299
rect 24852 25280 24854 25299
rect 24865 25294 24868 25299
rect 24876 25294 24878 25299
rect 24875 25280 24878 25294
rect 24841 25279 24875 25280
rect -14207 25275 -883 25279
rect -14100 25272 -14098 25275
rect -14100 25256 -14097 25272
rect -14111 25255 -14077 25256
rect -14004 25255 -14002 25275
rect -13788 25255 -13786 25275
rect -13428 25255 -13426 25275
rect -12852 25255 -12849 25272
rect -12756 25255 -12754 25275
rect -12636 25255 -12634 25275
rect -12348 25256 -12346 25275
rect -12359 25255 -12325 25256
rect -12252 25255 -12250 25275
rect -12156 25255 -12154 25275
rect -12060 25255 -12058 25275
rect -11772 25255 -11770 25275
rect -11759 25255 -11701 25256
rect -11676 25255 -11674 25275
rect -11508 25255 -11506 25275
rect -11436 25255 -11434 25275
rect -11412 25255 -11410 25275
rect -11340 25255 -11338 25275
rect -11196 25255 -11194 25275
rect -11100 25255 -11098 25275
rect -10764 25255 -10762 25275
rect -10644 25255 -10642 25275
rect -9996 25255 -9994 25275
rect -9900 25255 -9898 25275
rect -9732 25255 -9730 25275
rect -9444 25255 -9442 25275
rect -9348 25255 -9346 25275
rect -9228 25255 -9226 25275
rect -9108 25255 -9106 25275
rect -8436 25255 -8434 25275
rect -8364 25255 -8362 25275
rect -8340 25255 -8338 25275
rect -8268 25255 -8266 25275
rect -8004 25255 -8002 25275
rect -7932 25255 -7930 25275
rect -7641 25272 -7627 25275
rect -7620 25272 -7617 25275
rect -7799 25255 -7765 25256
rect -7524 25255 -7522 25275
rect -7356 25255 -7354 25275
rect -7308 25255 -7306 25275
rect -7212 25255 -7210 25275
rect -7044 25255 -7042 25275
rect -6948 25255 -6946 25275
rect -6852 25255 -6850 25275
rect -6756 25255 -6754 25275
rect -6660 25255 -6658 25275
rect -6612 25255 -6610 25275
rect -6516 25255 -6514 25275
rect -6372 25255 -6370 25275
rect -6036 25256 -6034 25275
rect -6047 25255 -6013 25256
rect -5892 25255 -5890 25275
rect -5196 25255 -5194 25275
rect -5100 25255 -5098 25275
rect -4716 25255 -4714 25275
rect -4500 25255 -4498 25275
rect -4404 25255 -4402 25275
rect -4308 25255 -4306 25275
rect -4164 25255 -4162 25275
rect -4020 25255 -4018 25275
rect -3876 25255 -3874 25275
rect -3732 25255 -3730 25275
rect -3636 25255 -3634 25275
rect -3540 25255 -3538 25275
rect -3468 25255 -3466 25275
rect -3324 25255 -3322 25275
rect -3153 25272 -3139 25275
rect -3132 25272 -3129 25275
rect -3108 25255 -3106 25275
rect -3012 25255 -3010 25275
rect -2964 25255 -2962 25275
rect -2916 25255 -2914 25275
rect -2892 25255 -2890 25275
rect -2868 25255 -2866 25275
rect -2820 25255 -2818 25275
rect -2796 25255 -2794 25275
rect -2772 25255 -2770 25275
rect -2676 25255 -2674 25275
rect -2580 25255 -2578 25275
rect -2364 25255 -2362 25275
rect -2316 25255 -2314 25275
rect -2268 25255 -2266 25275
rect -2244 25255 -2242 25275
rect -2172 25255 -2170 25275
rect -2148 25255 -2146 25275
rect -2076 25255 -2074 25275
rect -2052 25255 -2050 25275
rect -1980 25255 -1978 25275
rect -1884 25255 -1882 25275
rect -1572 25255 -1570 25275
rect -1476 25255 -1474 25275
rect -1356 25255 -1354 25275
rect -1260 25255 -1258 25275
rect -1236 25255 -1234 25275
rect -1140 25255 -1138 25275
rect -897 25272 -883 25275
rect -876 25275 8501 25279
rect -876 25272 -859 25275
rect -876 25255 -874 25272
rect -708 25256 -706 25275
rect -719 25255 -685 25256
rect -660 25255 -658 25275
rect -612 25255 -610 25275
rect -492 25255 -490 25275
rect -444 25255 -442 25275
rect -396 25255 -394 25275
rect -348 25255 -346 25275
rect -300 25255 -298 25275
rect -276 25255 -274 25275
rect -12 25255 -10 25275
rect 156 25255 158 25275
rect 204 25255 206 25275
rect 252 25255 254 25275
rect 348 25255 350 25275
rect 468 25255 470 25275
rect 492 25255 494 25275
rect 564 25255 566 25275
rect 588 25255 590 25275
rect 636 25255 638 25275
rect 660 25255 662 25275
rect 732 25255 734 25275
rect 1092 25255 1094 25275
rect 1140 25255 1142 25275
rect 1236 25255 1238 25275
rect 1308 25255 1310 25275
rect 1332 25255 1334 25275
rect 1380 25255 1382 25275
rect 1428 25255 1430 25275
rect 1476 25255 1478 25275
rect 1692 25255 1694 25275
rect 1788 25255 1790 25275
rect 2028 25255 2030 25275
rect 2076 25255 2078 25275
rect 2100 25255 2102 25275
rect 2124 25255 2126 25275
rect 2244 25255 2246 25275
rect 2412 25255 2414 25275
rect 2460 25255 2462 25275
rect 2508 25255 2510 25275
rect 2604 25255 2606 25275
rect 2772 25255 2774 25275
rect 2868 25255 2870 25275
rect 2940 25255 2942 25275
rect 3012 25255 3014 25275
rect 3108 25255 3110 25275
rect 3337 25270 3340 25275
rect 3348 25270 3350 25275
rect 3347 25256 3350 25270
rect 3396 25255 3398 25275
rect 3564 25255 3566 25275
rect 3636 25255 3638 25275
rect 3660 25255 3662 25275
rect 3732 25255 3734 25275
rect 3780 25255 3782 25275
rect 3828 25255 3830 25275
rect 3924 25255 3926 25275
rect 4020 25255 4022 25275
rect 4023 25272 4037 25275
rect 4092 25255 4094 25275
rect 4119 25272 4133 25275
rect 4188 25255 4190 25275
rect 4215 25272 4229 25275
rect 4308 25255 4310 25275
rect 4311 25272 4325 25275
rect 4404 25255 4406 25275
rect 4407 25272 4421 25275
rect 4500 25255 4502 25275
rect 4596 25255 4598 25275
rect 4692 25255 4694 25275
rect 4860 25255 4862 25275
rect 4956 25255 4958 25275
rect 4980 25255 4982 25275
rect 5052 25255 5054 25275
rect 5124 25255 5126 25275
rect 5220 25255 5222 25275
rect 5268 25255 5270 25275
rect 5388 25255 5390 25275
rect 5484 25255 5486 25275
rect 5508 25255 5510 25275
rect 5532 25255 5534 25275
rect 5628 25255 5630 25275
rect 5652 25255 5654 25275
rect 5748 25255 5750 25275
rect 5796 25255 5798 25275
rect 5844 25255 5846 25275
rect 5892 25255 5894 25275
rect 6132 25255 6134 25275
rect 6228 25255 6230 25275
rect 6252 25255 6254 25275
rect 6276 25255 6278 25275
rect 6324 25255 6326 25275
rect 6372 25255 6374 25275
rect 6420 25255 6422 25275
rect 6492 25255 6494 25275
rect 6516 25255 6518 25275
rect 6588 25255 6590 25275
rect 6612 25255 6614 25275
rect 6660 25255 6662 25275
rect 6684 25255 6686 25275
rect 6708 25255 6710 25275
rect 6780 25255 6782 25275
rect 6804 25255 6806 25275
rect 6900 25255 6902 25275
rect 6924 25255 6926 25275
rect 7020 25255 7022 25275
rect 7164 25255 7166 25275
rect 7236 25255 7238 25275
rect 7332 25255 7334 25275
rect 7380 25255 7382 25275
rect 7428 25255 7430 25275
rect 7452 25255 7454 25275
rect 7476 25255 7478 25275
rect 7524 25255 7526 25275
rect 7548 25255 7550 25275
rect 7572 25255 7574 25275
rect 7620 25255 7622 25275
rect 7644 25255 7646 25275
rect 7668 25255 7670 25275
rect 7908 25255 7910 25275
rect 7956 25255 7958 25275
rect 8124 25255 8126 25275
rect 8268 25256 8270 25275
rect 8257 25255 8291 25256
rect 8340 25255 8342 25275
rect 8364 25255 8366 25275
rect 8487 25272 8501 25275
rect 8511 25275 19397 25279
rect 8511 25272 8525 25275
rect 8652 25255 8654 25275
rect 8700 25255 8702 25275
rect 8748 25255 8750 25275
rect 8820 25255 8822 25275
rect 8844 25255 8846 25275
rect 8868 25255 8870 25275
rect 9516 25255 9518 25275
rect 9660 25255 9662 25275
rect 9684 25255 9686 25275
rect 9756 25255 9758 25275
rect 9780 25255 9782 25275
rect 9804 25255 9806 25275
rect 9852 25255 9854 25275
rect 9900 25255 9902 25275
rect 9948 25255 9950 25275
rect 9961 25255 9995 25256
rect 10044 25255 10046 25275
rect 10116 25255 10118 25275
rect 10188 25255 10190 25275
rect 10212 25255 10214 25275
rect 10284 25255 10286 25275
rect 10332 25255 10334 25275
rect 10380 25255 10382 25275
rect 10428 25255 10430 25275
rect 10476 25255 10478 25275
rect 10500 25255 10502 25275
rect 10524 25255 10526 25275
rect 10572 25255 10574 25275
rect 10596 25255 10598 25275
rect 10620 25255 10622 25275
rect 10692 25256 10694 25275
rect 10681 25255 10715 25256
rect 10716 25255 10718 25275
rect 10788 25255 10790 25275
rect 10956 25255 10958 25275
rect 11004 25255 11006 25275
rect 11052 25255 11054 25275
rect 11100 25255 11102 25275
rect 11172 25255 11174 25275
rect 11220 25255 11222 25275
rect 11340 25255 11342 25275
rect 11436 25255 11438 25275
rect 11532 25255 11534 25275
rect 11580 25255 11582 25275
rect 11628 25255 11630 25275
rect 11676 25255 11678 25275
rect 11724 25255 11726 25275
rect 11772 25255 11774 25275
rect 11796 25255 11798 25275
rect 11892 25255 11894 25275
rect 11988 25255 11990 25275
rect 12025 25255 12059 25256
rect 12060 25255 12062 25275
rect 12132 25255 12134 25275
rect 12228 25255 12230 25275
rect 12276 25255 12278 25275
rect 12324 25255 12326 25275
rect 12420 25255 12422 25275
rect 12444 25255 12446 25275
rect 12492 25255 12494 25275
rect 12516 25255 12518 25275
rect 12540 25255 12542 25275
rect 12588 25255 12590 25275
rect 12636 25255 12638 25275
rect 12732 25255 12734 25275
rect 12756 25255 12758 25275
rect 12804 25255 12806 25275
rect 12828 25255 12830 25275
rect 12972 25255 12974 25275
rect 13044 25255 13046 25275
rect 13068 25255 13070 25275
rect 13116 25255 13118 25275
rect 13284 25255 13286 25275
rect 13332 25255 13334 25275
rect 13572 25255 13574 25275
rect 13620 25255 13622 25275
rect 13668 25255 13670 25275
rect 13716 25255 13718 25275
rect 13764 25255 13766 25275
rect 13860 25255 13862 25275
rect 13956 25255 13958 25275
rect 14004 25255 14006 25275
rect 14100 25255 14102 25275
rect 15180 25255 15182 25275
rect 15276 25255 15278 25275
rect 15420 25255 15422 25275
rect 15492 25255 15494 25275
rect 15660 25255 15662 25275
rect 15708 25255 15710 25275
rect 15732 25255 15734 25275
rect 15756 25255 15758 25275
rect 15804 25255 15806 25275
rect 15828 25255 15830 25275
rect 15852 25255 15854 25275
rect 15900 25255 15902 25275
rect 15948 25255 15950 25275
rect 16044 25255 16046 25275
rect 16068 25255 16070 25275
rect 16164 25255 16166 25275
rect 16260 25255 16262 25275
rect 16332 25255 16334 25275
rect 16548 25255 16550 25275
rect 16572 25255 16574 25275
rect 16620 25255 16622 25275
rect 16668 25255 16670 25275
rect 16716 25255 16718 25275
rect 16764 25255 16766 25275
rect 16812 25255 16814 25275
rect 16884 25255 16886 25275
rect 16908 25255 16910 25275
rect 16980 25255 16982 25275
rect 17148 25255 17150 25275
rect 17196 25255 17198 25275
rect 17220 25255 17222 25275
rect 17292 25255 17294 25275
rect 17316 25255 17318 25275
rect 18132 25255 18134 25275
rect 18228 25255 18230 25275
rect 18492 25255 18494 25275
rect 18516 25255 18518 25275
rect 18564 25255 18566 25275
rect 18612 25255 18614 25275
rect 18660 25255 18662 25275
rect 18756 25255 18758 25275
rect 18900 25255 18902 25275
rect 18924 25255 18926 25275
rect 18996 25255 18998 25275
rect 19020 25255 19022 25275
rect 19092 25255 19094 25275
rect 19116 25256 19118 25275
rect 19105 25255 19139 25256
rect 19140 25255 19142 25275
rect 19188 25255 19190 25275
rect 19236 25255 19238 25275
rect 19383 25272 19397 25275
rect 19407 25275 24875 25279
rect 19407 25272 19421 25275
rect 19788 25255 19790 25275
rect 19836 25255 19838 25275
rect 19860 25255 19862 25275
rect 19884 25255 19886 25275
rect 19932 25255 19934 25275
rect 19956 25255 19958 25275
rect 19980 25255 19982 25275
rect 20028 25255 20030 25275
rect 20052 25255 20054 25275
rect 20076 25255 20078 25275
rect 20148 25256 20150 25275
rect 20113 25255 20171 25256
rect 20172 25255 20174 25275
rect 20196 25255 20198 25275
rect 20268 25255 20270 25275
rect 20292 25255 20294 25275
rect 20388 25255 20390 25275
rect 20412 25255 20414 25275
rect 20508 25255 20510 25275
rect 20604 25255 20606 25275
rect 20964 25255 20966 25275
rect 21012 25255 21014 25275
rect 21108 25255 21110 25275
rect 21204 25255 21206 25275
rect 21300 25255 21302 25275
rect 21324 25255 21326 25275
rect 21444 25255 21446 25275
rect 21468 25255 21470 25275
rect 21564 25255 21566 25275
rect 21588 25255 21590 25275
rect 21684 25255 21686 25275
rect 21708 25255 21710 25275
rect 21828 25255 21830 25275
rect 21924 25255 21926 25275
rect 22068 25255 22070 25275
rect 22188 25255 22190 25275
rect 22212 25255 22214 25275
rect 22884 25255 22886 25275
rect 22980 25255 22982 25275
rect 23076 25255 23078 25275
rect 23100 25255 23102 25275
rect 23124 25255 23126 25275
rect 23244 25255 23246 25275
rect 23340 25255 23342 25275
rect 23412 25255 23414 25275
rect 23460 25255 23462 25275
rect 23508 25255 23510 25275
rect 23556 25255 23558 25275
rect 23604 25255 23606 25275
rect 23652 25255 23654 25275
rect 23676 25255 23678 25275
rect 23700 25255 23702 25275
rect 23772 25255 23774 25275
rect 23796 25255 23798 25275
rect 23916 25255 23918 25275
rect 24012 25255 24014 25275
rect 24060 25255 24062 25275
rect 24156 25255 24158 25275
rect 24492 25255 24494 25275
rect 24516 25255 24518 25275
rect 24588 25255 24590 25275
rect 24612 25255 24614 25275
rect 24684 25255 24686 25275
rect 24756 25255 24758 25275
rect 24780 25256 24782 25275
rect 24841 25270 24844 25275
rect 24852 25270 24854 25275
rect 24851 25256 24854 25270
rect 24769 25255 24803 25256
rect -14111 25251 -12859 25255
rect -14111 25248 -14107 25251
rect -14100 25248 -14097 25251
rect -14004 25248 -14002 25251
rect -14004 25232 -14001 25248
rect -14015 25231 -13981 25232
rect -13788 25231 -13786 25251
rect -13428 25231 -13426 25251
rect -12873 25248 -12859 25251
rect -12852 25251 3413 25255
rect -12852 25248 -12835 25251
rect -12852 25231 -12850 25248
rect -12756 25231 -12754 25251
rect -12636 25231 -12634 25251
rect -12359 25246 -12356 25251
rect -12348 25246 -12346 25251
rect -12349 25232 -12346 25246
rect -12252 25248 -12250 25251
rect -12252 25231 -12249 25248
rect -12156 25231 -12154 25251
rect -12060 25231 -12058 25251
rect -11772 25231 -11770 25251
rect -11676 25231 -11674 25251
rect -11652 25231 -11649 25248
rect -11508 25231 -11506 25251
rect -11436 25231 -11434 25251
rect -11412 25231 -11410 25251
rect -11340 25231 -11338 25251
rect -11196 25231 -11194 25251
rect -11100 25231 -11098 25251
rect -10764 25231 -10762 25251
rect -10644 25231 -10642 25251
rect -10103 25231 -10069 25232
rect -9996 25231 -9994 25251
rect -9900 25231 -9898 25251
rect -9732 25231 -9730 25251
rect -9609 25248 -9595 25251
rect -9444 25231 -9442 25251
rect -9348 25231 -9346 25251
rect -9228 25231 -9226 25251
rect -9108 25231 -9106 25251
rect -8505 25248 -8491 25251
rect -8436 25231 -8434 25251
rect -8364 25231 -8362 25251
rect -8340 25231 -8338 25251
rect -8313 25248 -8299 25251
rect -8268 25231 -8266 25251
rect -8004 25231 -8002 25251
rect -7932 25231 -7930 25251
rect -7524 25231 -7522 25251
rect -7356 25231 -7354 25251
rect -7308 25231 -7306 25251
rect -7212 25231 -7210 25251
rect -7044 25231 -7042 25251
rect -6948 25231 -6946 25251
rect -6852 25231 -6850 25251
rect -6756 25231 -6754 25251
rect -6660 25231 -6658 25251
rect -6612 25231 -6610 25251
rect -6516 25231 -6514 25251
rect -6372 25231 -6370 25251
rect -6047 25246 -6044 25251
rect -6036 25246 -6034 25251
rect -6037 25232 -6034 25246
rect -5892 25231 -5890 25251
rect -5447 25231 -5389 25232
rect -5196 25231 -5194 25251
rect -5100 25231 -5098 25251
rect -4716 25231 -4714 25251
rect -4500 25231 -4498 25251
rect -4404 25231 -4402 25251
rect -4308 25231 -4306 25251
rect -4164 25231 -4162 25251
rect -4020 25231 -4018 25251
rect -3876 25231 -3874 25251
rect -3732 25231 -3730 25251
rect -3636 25231 -3634 25251
rect -3540 25231 -3538 25251
rect -3468 25231 -3466 25251
rect -3324 25231 -3322 25251
rect -3108 25231 -3106 25251
rect -3012 25231 -3010 25251
rect -2964 25231 -2962 25251
rect -2916 25231 -2914 25251
rect -2892 25231 -2890 25251
rect -2868 25231 -2866 25251
rect -2820 25231 -2818 25251
rect -2796 25231 -2794 25251
rect -2772 25231 -2770 25251
rect -2676 25231 -2674 25251
rect -2580 25232 -2578 25251
rect -2591 25231 -2557 25232
rect -2364 25231 -2362 25251
rect -2316 25231 -2314 25251
rect -2268 25232 -2266 25251
rect -2279 25231 -2245 25232
rect -2244 25231 -2242 25251
rect -2172 25231 -2170 25251
rect -2148 25231 -2146 25251
rect -2076 25231 -2074 25251
rect -2052 25231 -2050 25251
rect -1980 25231 -1978 25251
rect -1884 25231 -1882 25251
rect -1572 25231 -1570 25251
rect -1476 25231 -1474 25251
rect -1356 25231 -1354 25251
rect -1260 25231 -1258 25251
rect -1236 25231 -1234 25251
rect -1140 25231 -1138 25251
rect -876 25231 -874 25251
rect -719 25246 -716 25251
rect -708 25246 -706 25251
rect -709 25232 -706 25246
rect -660 25231 -658 25251
rect -612 25248 -610 25251
rect -612 25232 -609 25248
rect -623 25231 -589 25232
rect -492 25231 -490 25251
rect -444 25231 -442 25251
rect -396 25231 -394 25251
rect -348 25231 -346 25251
rect -300 25232 -298 25251
rect -311 25231 -277 25232
rect -276 25231 -274 25251
rect -12 25231 -10 25251
rect 156 25231 158 25251
rect 204 25231 206 25251
rect 252 25231 254 25251
rect 348 25231 350 25251
rect 468 25231 470 25251
rect 492 25231 494 25251
rect 564 25231 566 25251
rect 588 25231 590 25251
rect 636 25231 638 25251
rect 660 25231 662 25251
rect 732 25231 734 25251
rect 1092 25231 1094 25251
rect 1140 25231 1142 25251
rect 1236 25231 1238 25251
rect 1308 25231 1310 25251
rect 1332 25231 1334 25251
rect 1380 25231 1382 25251
rect 1428 25231 1430 25251
rect 1476 25231 1478 25251
rect 1692 25231 1694 25251
rect 1788 25231 1790 25251
rect 2028 25231 2030 25251
rect 2076 25231 2078 25251
rect 2100 25231 2102 25251
rect 2124 25231 2126 25251
rect 2244 25231 2246 25251
rect 2412 25231 2414 25251
rect 2460 25231 2462 25251
rect 2508 25231 2510 25251
rect 2604 25231 2606 25251
rect 2772 25231 2774 25251
rect 2868 25231 2870 25251
rect 2940 25231 2942 25251
rect 3012 25231 3014 25251
rect 3108 25231 3110 25251
rect 3396 25231 3398 25251
rect 3399 25248 3413 25251
rect 3423 25251 24803 25255
rect 3423 25248 3437 25251
rect 3564 25231 3566 25251
rect 3636 25231 3638 25251
rect 3660 25231 3662 25251
rect 3732 25231 3734 25251
rect 3780 25231 3782 25251
rect 3828 25231 3830 25251
rect 3924 25231 3926 25251
rect 4020 25231 4022 25251
rect 4092 25231 4094 25251
rect 4188 25231 4190 25251
rect 4308 25231 4310 25251
rect 4404 25231 4406 25251
rect 4500 25231 4502 25251
rect 4596 25231 4598 25251
rect 4692 25231 4694 25251
rect 4860 25231 4862 25251
rect 4956 25231 4958 25251
rect 4980 25231 4982 25251
rect 5052 25231 5054 25251
rect 5124 25231 5126 25251
rect 5220 25231 5222 25251
rect 5268 25231 5270 25251
rect 5388 25231 5390 25251
rect 5484 25231 5486 25251
rect 5508 25231 5510 25251
rect 5532 25231 5534 25251
rect 5628 25231 5630 25251
rect 5652 25231 5654 25251
rect 5748 25231 5750 25251
rect 5796 25231 5798 25251
rect 5844 25231 5846 25251
rect 5892 25231 5894 25251
rect 6132 25231 6134 25251
rect 6228 25231 6230 25251
rect 6252 25231 6254 25251
rect 6276 25231 6278 25251
rect 6324 25231 6326 25251
rect 6372 25231 6374 25251
rect 6420 25231 6422 25251
rect 6492 25231 6494 25251
rect 6516 25231 6518 25251
rect 6588 25231 6590 25251
rect 6612 25231 6614 25251
rect 6660 25231 6662 25251
rect 6684 25231 6686 25251
rect 6708 25231 6710 25251
rect 6780 25231 6782 25251
rect 6804 25231 6806 25251
rect 6900 25231 6902 25251
rect 6924 25231 6926 25251
rect 7020 25231 7022 25251
rect 7164 25231 7166 25251
rect 7236 25231 7238 25251
rect 7332 25232 7334 25251
rect 7297 25231 7355 25232
rect 7380 25231 7382 25251
rect 7428 25231 7430 25251
rect 7452 25231 7454 25251
rect 7476 25231 7478 25251
rect 7524 25231 7526 25251
rect 7548 25231 7550 25251
rect 7572 25231 7574 25251
rect 7620 25231 7622 25251
rect 7644 25231 7646 25251
rect 7668 25231 7670 25251
rect 7908 25231 7910 25251
rect 7956 25231 7958 25251
rect 8124 25231 8126 25251
rect 8257 25246 8260 25251
rect 8268 25246 8270 25251
rect 8267 25232 8270 25246
rect 8340 25231 8342 25251
rect 8364 25248 8366 25251
rect 8364 25231 8367 25248
rect 8652 25231 8654 25251
rect 8700 25231 8702 25251
rect 8748 25231 8750 25251
rect 8820 25231 8822 25251
rect 8844 25231 8846 25251
rect 8868 25231 8870 25251
rect 9516 25231 9518 25251
rect 9660 25231 9662 25251
rect 9684 25231 9686 25251
rect 9756 25231 9758 25251
rect 9780 25231 9782 25251
rect 9804 25231 9806 25251
rect 9852 25231 9854 25251
rect 9900 25231 9902 25251
rect 9948 25231 9950 25251
rect 10044 25231 10046 25251
rect 10116 25231 10118 25251
rect 10188 25231 10190 25251
rect 10212 25231 10214 25251
rect 10284 25231 10286 25251
rect 10332 25231 10334 25251
rect 10380 25231 10382 25251
rect 10428 25231 10430 25251
rect 10476 25231 10478 25251
rect 10500 25231 10502 25251
rect 10524 25231 10526 25251
rect 10572 25231 10574 25251
rect 10596 25231 10598 25251
rect 10620 25231 10622 25251
rect 10681 25246 10684 25251
rect 10692 25246 10694 25251
rect 10691 25232 10694 25246
rect 10716 25231 10718 25251
rect 10788 25248 10790 25251
rect 10788 25231 10791 25248
rect 10956 25231 10958 25251
rect 11004 25231 11006 25251
rect 11052 25231 11054 25251
rect 11100 25231 11102 25251
rect 11172 25231 11174 25251
rect 11220 25231 11222 25251
rect 11340 25231 11342 25251
rect 11436 25231 11438 25251
rect 11473 25231 11507 25232
rect 11532 25231 11534 25251
rect 11580 25231 11582 25251
rect 11628 25231 11630 25251
rect 11676 25231 11678 25251
rect 11724 25231 11726 25251
rect 11772 25231 11774 25251
rect 11796 25231 11798 25251
rect 11892 25231 11894 25251
rect 11988 25231 11990 25251
rect 12060 25231 12062 25251
rect 12132 25248 12134 25251
rect 12132 25231 12135 25248
rect 12228 25231 12230 25251
rect 12276 25231 12278 25251
rect 12324 25231 12326 25251
rect 12420 25231 12422 25251
rect 12444 25231 12446 25251
rect 12492 25231 12494 25251
rect 12516 25231 12518 25251
rect 12540 25231 12542 25251
rect 12588 25231 12590 25251
rect 12636 25231 12638 25251
rect 12732 25231 12734 25251
rect 12756 25231 12758 25251
rect 12804 25231 12806 25251
rect 12828 25231 12830 25251
rect 12972 25231 12974 25251
rect 13044 25231 13046 25251
rect 13068 25231 13070 25251
rect 13116 25231 13118 25251
rect 13284 25231 13286 25251
rect 13332 25231 13334 25251
rect 13572 25231 13574 25251
rect 13620 25231 13622 25251
rect 13668 25231 13670 25251
rect 13716 25231 13718 25251
rect 13764 25231 13766 25251
rect 13860 25231 13862 25251
rect 13956 25231 13958 25251
rect 14004 25231 14006 25251
rect 14100 25231 14102 25251
rect 15180 25231 15182 25251
rect 15276 25231 15278 25251
rect 15420 25231 15422 25251
rect 15492 25231 15494 25251
rect 15660 25231 15662 25251
rect 15708 25231 15710 25251
rect 15732 25231 15734 25251
rect 15756 25231 15758 25251
rect 15804 25231 15806 25251
rect 15828 25231 15830 25251
rect 15852 25231 15854 25251
rect 15900 25232 15902 25251
rect 15865 25231 15923 25232
rect 15948 25231 15950 25251
rect 16044 25231 16046 25251
rect 16068 25231 16070 25251
rect 16164 25231 16166 25251
rect 16260 25231 16262 25251
rect 16332 25231 16334 25251
rect 16548 25231 16550 25251
rect 16572 25231 16574 25251
rect 16620 25231 16622 25251
rect 16668 25231 16670 25251
rect 16716 25231 16718 25251
rect 16764 25231 16766 25251
rect 16812 25231 16814 25251
rect 16884 25231 16886 25251
rect 16908 25231 16910 25251
rect 16980 25231 16982 25251
rect 17148 25231 17150 25251
rect 17196 25231 17198 25251
rect 17220 25231 17222 25251
rect 17292 25231 17294 25251
rect 17316 25231 17318 25251
rect 18132 25231 18134 25251
rect 18228 25231 18230 25251
rect 18492 25231 18494 25251
rect 18516 25231 18518 25251
rect 18564 25231 18566 25251
rect 18612 25231 18614 25251
rect 18660 25231 18662 25251
rect 18756 25231 18758 25251
rect 18900 25231 18902 25251
rect 18924 25231 18926 25251
rect 18996 25231 18998 25251
rect 19020 25231 19022 25251
rect 19092 25231 19094 25251
rect 19105 25246 19108 25251
rect 19116 25246 19118 25251
rect 19115 25232 19118 25246
rect 19140 25231 19142 25251
rect 19188 25231 19190 25251
rect 19236 25231 19238 25251
rect 19788 25231 19790 25251
rect 19836 25231 19838 25251
rect 19860 25231 19862 25251
rect 19884 25231 19886 25251
rect 19932 25232 19934 25251
rect 19897 25231 19955 25232
rect 19956 25231 19958 25251
rect 19980 25231 19982 25251
rect 20028 25231 20030 25251
rect 20052 25231 20054 25251
rect 20076 25231 20078 25251
rect 20113 25246 20116 25251
rect 20137 25246 20140 25251
rect 20148 25246 20150 25251
rect 20123 25232 20126 25246
rect 20147 25232 20150 25246
rect 20124 25231 20126 25232
rect 20172 25231 20174 25251
rect 20196 25231 20198 25251
rect 20268 25231 20270 25251
rect 20292 25231 20294 25251
rect 20388 25231 20390 25251
rect 20412 25231 20414 25251
rect 20508 25231 20510 25251
rect 20604 25231 20606 25251
rect 20964 25231 20966 25251
rect 21012 25231 21014 25251
rect 21108 25231 21110 25251
rect 21204 25231 21206 25251
rect 21300 25231 21302 25251
rect 21324 25231 21326 25251
rect 21444 25231 21446 25251
rect 21468 25231 21470 25251
rect 21564 25231 21566 25251
rect 21588 25231 21590 25251
rect 21684 25231 21686 25251
rect 21708 25231 21710 25251
rect 21828 25231 21830 25251
rect 21924 25231 21926 25251
rect 22068 25231 22070 25251
rect 22188 25231 22190 25251
rect 22212 25231 22214 25251
rect 22884 25231 22886 25251
rect 22980 25231 22982 25251
rect 23076 25231 23078 25251
rect 23100 25231 23102 25251
rect 23124 25231 23126 25251
rect 23244 25231 23246 25251
rect 23340 25231 23342 25251
rect 23412 25231 23414 25251
rect 23460 25231 23462 25251
rect 23508 25231 23510 25251
rect 23556 25231 23558 25251
rect 23604 25231 23606 25251
rect 23652 25231 23654 25251
rect 23676 25231 23678 25251
rect 23700 25231 23702 25251
rect 23772 25231 23774 25251
rect 23796 25231 23798 25251
rect 23916 25231 23918 25251
rect 24012 25231 24014 25251
rect 24060 25231 24062 25251
rect 24156 25231 24158 25251
rect 24492 25231 24494 25251
rect 24516 25231 24518 25251
rect 24588 25231 24590 25251
rect 24612 25231 24614 25251
rect 24684 25231 24686 25251
rect 24756 25232 24758 25251
rect 24769 25246 24772 25251
rect 24780 25246 24782 25251
rect 24779 25232 24782 25246
rect 24745 25231 24779 25232
rect -14015 25227 -11659 25231
rect -14015 25224 -14011 25227
rect -14004 25224 -14001 25227
rect -13895 25207 -13861 25208
rect -13788 25207 -13786 25227
rect -13428 25207 -13426 25227
rect -12852 25207 -12850 25227
rect -12756 25208 -12754 25227
rect -12767 25207 -12733 25208
rect -12636 25207 -12634 25227
rect -12273 25224 -12259 25227
rect -12252 25224 -12249 25227
rect -12263 25207 -12229 25208
rect -12156 25207 -12154 25227
rect -12060 25207 -12058 25227
rect -11772 25207 -11770 25227
rect -11676 25207 -11674 25227
rect -11673 25224 -11659 25227
rect -11652 25227 20213 25231
rect -11652 25224 -11635 25227
rect -11652 25207 -11650 25224
rect -11508 25207 -11506 25227
rect -11436 25207 -11434 25227
rect -11412 25207 -11410 25227
rect -11340 25207 -11338 25227
rect -11196 25207 -11194 25227
rect -11100 25207 -11098 25227
rect -10764 25207 -10762 25227
rect -10644 25207 -10642 25227
rect -9996 25224 -9994 25227
rect -9996 25207 -9993 25224
rect -9900 25207 -9898 25227
rect -9732 25207 -9730 25227
rect -9444 25207 -9442 25227
rect -9348 25207 -9346 25227
rect -9228 25207 -9226 25227
rect -9108 25207 -9106 25227
rect -8436 25207 -8434 25227
rect -8364 25207 -8362 25227
rect -8340 25207 -8338 25227
rect -8268 25207 -8266 25227
rect -8004 25207 -8002 25227
rect -7932 25207 -7930 25227
rect -7713 25224 -7699 25227
rect -7524 25207 -7522 25227
rect -7356 25207 -7354 25227
rect -7308 25207 -7306 25227
rect -7212 25207 -7210 25227
rect -7044 25207 -7042 25227
rect -6948 25207 -6946 25227
rect -6852 25207 -6850 25227
rect -6756 25207 -6754 25227
rect -6660 25207 -6658 25227
rect -6612 25207 -6610 25227
rect -6516 25207 -6514 25227
rect -6372 25207 -6370 25227
rect -5961 25224 -5947 25227
rect -6071 25207 -6037 25208
rect -5892 25207 -5890 25227
rect -5447 25222 -5444 25227
rect -5437 25208 -5434 25222
rect -5436 25207 -5434 25208
rect -5340 25207 -5337 25224
rect -5196 25207 -5194 25227
rect -5100 25207 -5098 25227
rect -4716 25207 -4714 25227
rect -4500 25207 -4498 25227
rect -4404 25207 -4402 25227
rect -4308 25207 -4306 25227
rect -4164 25207 -4162 25227
rect -4020 25207 -4018 25227
rect -3876 25207 -3874 25227
rect -3732 25207 -3730 25227
rect -3636 25207 -3634 25227
rect -3540 25207 -3538 25227
rect -3468 25207 -3466 25227
rect -3324 25207 -3322 25227
rect -3108 25207 -3106 25227
rect -3012 25207 -3010 25227
rect -2964 25207 -2962 25227
rect -2916 25207 -2914 25227
rect -2892 25207 -2890 25227
rect -2868 25207 -2866 25227
rect -2820 25207 -2818 25227
rect -2796 25207 -2794 25227
rect -2772 25207 -2770 25227
rect -2676 25207 -2674 25227
rect -2591 25222 -2588 25227
rect -2580 25222 -2578 25227
rect -2581 25208 -2578 25222
rect -2364 25207 -2362 25227
rect -2316 25207 -2314 25227
rect -2279 25222 -2276 25227
rect -2268 25222 -2266 25227
rect -2269 25208 -2266 25222
rect -2244 25207 -2242 25227
rect -2172 25224 -2170 25227
rect -2172 25207 -2169 25224
rect -2148 25207 -2146 25227
rect -2076 25207 -2074 25227
rect -2052 25207 -2050 25227
rect -1980 25207 -1978 25227
rect -1884 25207 -1882 25227
rect -1572 25207 -1570 25227
rect -1476 25207 -1474 25227
rect -1356 25207 -1354 25227
rect -1260 25207 -1258 25227
rect -1236 25207 -1234 25227
rect -1140 25207 -1138 25227
rect -876 25207 -874 25227
rect -660 25207 -658 25227
rect -633 25224 -619 25227
rect -612 25224 -609 25227
rect -492 25207 -490 25227
rect -444 25207 -442 25227
rect -396 25207 -394 25227
rect -348 25207 -346 25227
rect -311 25222 -308 25227
rect -300 25222 -298 25227
rect -301 25208 -298 25222
rect -276 25207 -274 25227
rect -12 25207 -10 25227
rect 156 25207 158 25227
rect 204 25207 206 25227
rect 252 25207 254 25227
rect 348 25207 350 25227
rect 468 25207 470 25227
rect 492 25207 494 25227
rect 564 25207 566 25227
rect 588 25207 590 25227
rect 636 25207 638 25227
rect 660 25207 662 25227
rect 732 25207 734 25227
rect 1092 25207 1094 25227
rect 1140 25207 1142 25227
rect 1236 25207 1238 25227
rect 1249 25207 1307 25208
rect 1308 25207 1310 25227
rect 1332 25207 1334 25227
rect 1380 25207 1382 25227
rect 1428 25207 1430 25227
rect 1476 25207 1478 25227
rect 1692 25207 1694 25227
rect 1788 25207 1790 25227
rect 2028 25207 2030 25227
rect 2076 25207 2078 25227
rect 2100 25207 2102 25227
rect 2124 25207 2126 25227
rect 2244 25207 2246 25227
rect 2412 25207 2414 25227
rect 2460 25207 2462 25227
rect 2508 25207 2510 25227
rect 2604 25207 2606 25227
rect 2772 25207 2774 25227
rect 2868 25207 2870 25227
rect 2940 25207 2942 25227
rect 3012 25207 3014 25227
rect 3108 25207 3110 25227
rect 3396 25207 3398 25227
rect 3564 25207 3566 25227
rect 3636 25207 3638 25227
rect 3660 25207 3662 25227
rect 3732 25207 3734 25227
rect 3780 25207 3782 25227
rect 3828 25207 3830 25227
rect 3924 25207 3926 25227
rect 4020 25207 4022 25227
rect 4092 25207 4094 25227
rect 4188 25207 4190 25227
rect 4308 25207 4310 25227
rect 4404 25207 4406 25227
rect 4500 25207 4502 25227
rect 4596 25207 4598 25227
rect 4633 25207 4667 25208
rect 4692 25207 4694 25227
rect 4860 25207 4862 25227
rect 4956 25207 4958 25227
rect 4980 25207 4982 25227
rect 5052 25207 5054 25227
rect 5124 25207 5126 25227
rect 5220 25207 5222 25227
rect 5268 25207 5270 25227
rect 5388 25207 5390 25227
rect 5484 25207 5486 25227
rect 5508 25207 5510 25227
rect 5532 25207 5534 25227
rect 5628 25207 5630 25227
rect 5652 25207 5654 25227
rect 5748 25207 5750 25227
rect 5796 25207 5798 25227
rect 5844 25207 5846 25227
rect 5892 25207 5894 25227
rect 6132 25207 6134 25227
rect 6228 25207 6230 25227
rect 6252 25207 6254 25227
rect 6276 25207 6278 25227
rect 6324 25207 6326 25227
rect 6372 25207 6374 25227
rect 6420 25207 6422 25227
rect 6492 25207 6494 25227
rect 6516 25207 6518 25227
rect 6588 25207 6590 25227
rect 6612 25207 6614 25227
rect 6660 25207 6662 25227
rect 6684 25207 6686 25227
rect 6708 25207 6710 25227
rect 6780 25207 6782 25227
rect 6804 25207 6806 25227
rect 6900 25207 6902 25227
rect 6924 25207 6926 25227
rect 7020 25207 7022 25227
rect 7164 25207 7166 25227
rect 7236 25207 7238 25227
rect 7297 25222 7300 25227
rect 7321 25222 7324 25227
rect 7332 25222 7334 25227
rect 7307 25208 7310 25222
rect 7331 25208 7334 25222
rect 7308 25207 7310 25208
rect 7380 25207 7382 25227
rect 7428 25224 7430 25227
rect 7428 25207 7431 25224
rect 7452 25207 7454 25227
rect 7476 25207 7478 25227
rect 7524 25207 7526 25227
rect 7548 25207 7550 25227
rect 7572 25207 7574 25227
rect 7620 25207 7622 25227
rect 7644 25207 7646 25227
rect 7668 25207 7670 25227
rect 7908 25207 7910 25227
rect 7956 25207 7958 25227
rect 8124 25207 8126 25227
rect 8209 25207 8267 25208
rect 8340 25207 8342 25227
rect 8343 25224 8357 25227
rect 8364 25224 8367 25227
rect 8652 25207 8654 25227
rect 8700 25207 8702 25227
rect 8748 25207 8750 25227
rect 8820 25207 8822 25227
rect 8844 25207 8846 25227
rect 8868 25207 8870 25227
rect 9516 25207 9518 25227
rect 9660 25207 9662 25227
rect 9684 25207 9686 25227
rect 9756 25207 9758 25227
rect 9780 25207 9782 25227
rect 9804 25207 9806 25227
rect 9852 25207 9854 25227
rect 9900 25207 9902 25227
rect 9948 25207 9950 25227
rect 10044 25207 10046 25227
rect 10047 25224 10061 25227
rect 10116 25207 10118 25227
rect 10188 25207 10190 25227
rect 10212 25207 10214 25227
rect 10284 25207 10286 25227
rect 10332 25207 10334 25227
rect 10380 25207 10382 25227
rect 10428 25207 10430 25227
rect 10476 25207 10478 25227
rect 10500 25207 10502 25227
rect 10524 25207 10526 25227
rect 10572 25207 10574 25227
rect 10596 25207 10598 25227
rect 10620 25207 10622 25227
rect 10716 25207 10718 25227
rect 10767 25224 10781 25227
rect 10788 25224 10791 25227
rect 10956 25207 10958 25227
rect 11004 25207 11006 25227
rect 11052 25207 11054 25227
rect 11100 25207 11102 25227
rect 11172 25207 11174 25227
rect 11220 25207 11222 25227
rect 11340 25207 11342 25227
rect 11436 25207 11438 25227
rect 11532 25207 11534 25227
rect 11580 25224 11582 25227
rect 11580 25207 11583 25224
rect 11628 25207 11630 25227
rect 11676 25207 11678 25227
rect 11724 25207 11726 25227
rect 11772 25207 11774 25227
rect 11796 25207 11798 25227
rect 11892 25207 11894 25227
rect 11988 25207 11990 25227
rect 12060 25207 12062 25227
rect 12111 25224 12125 25227
rect 12132 25224 12135 25227
rect 12228 25207 12230 25227
rect 12276 25207 12278 25227
rect 12324 25207 12326 25227
rect 12420 25207 12422 25227
rect 12444 25207 12446 25227
rect 12492 25208 12494 25227
rect 12457 25207 12515 25208
rect 12516 25207 12518 25227
rect 12540 25207 12542 25227
rect 12588 25207 12590 25227
rect 12636 25207 12638 25227
rect 12732 25207 12734 25227
rect 12756 25207 12758 25227
rect 12804 25207 12806 25227
rect 12828 25207 12830 25227
rect 12972 25207 12974 25227
rect 13044 25207 13046 25227
rect 13068 25207 13070 25227
rect 13116 25207 13118 25227
rect 13284 25207 13286 25227
rect 13332 25207 13334 25227
rect 13572 25207 13574 25227
rect 13620 25207 13622 25227
rect 13668 25207 13670 25227
rect 13716 25207 13718 25227
rect 13764 25207 13766 25227
rect 13860 25207 13862 25227
rect 13956 25207 13958 25227
rect 14004 25207 14006 25227
rect 14100 25207 14102 25227
rect 15180 25207 15182 25227
rect 15276 25207 15278 25227
rect 15420 25207 15422 25227
rect 15492 25207 15494 25227
rect 15660 25207 15662 25227
rect 15708 25207 15710 25227
rect 15732 25207 15734 25227
rect 15756 25207 15758 25227
rect 15804 25207 15806 25227
rect 15828 25207 15830 25227
rect 15852 25207 15854 25227
rect 15889 25222 15892 25227
rect 15900 25222 15902 25227
rect 15899 25208 15902 25222
rect 15948 25207 15950 25227
rect 15972 25207 15975 25224
rect 16044 25207 16046 25227
rect 16068 25207 16070 25227
rect 16164 25207 16166 25227
rect 16260 25207 16262 25227
rect 16332 25207 16334 25227
rect 16548 25207 16550 25227
rect 16572 25207 16574 25227
rect 16620 25207 16622 25227
rect 16668 25207 16670 25227
rect 16716 25207 16718 25227
rect 16764 25207 16766 25227
rect 16812 25207 16814 25227
rect 16884 25207 16886 25227
rect 16908 25207 16910 25227
rect 16980 25207 16982 25227
rect 17148 25207 17150 25227
rect 17196 25207 17198 25227
rect 17220 25207 17222 25227
rect 17292 25207 17294 25227
rect 17316 25207 17318 25227
rect 18132 25207 18134 25227
rect 18228 25207 18230 25227
rect 18492 25207 18494 25227
rect 18516 25207 18518 25227
rect 18564 25207 18566 25227
rect 18612 25207 18614 25227
rect 18660 25207 18662 25227
rect 18756 25207 18758 25227
rect 18900 25207 18902 25227
rect 18924 25207 18926 25227
rect 18996 25207 18998 25227
rect 19020 25207 19022 25227
rect 19092 25207 19094 25227
rect 19140 25207 19142 25227
rect 19188 25207 19190 25227
rect 19191 25224 19205 25227
rect 19236 25207 19238 25227
rect 19788 25207 19790 25227
rect 19836 25207 19838 25227
rect 19860 25207 19862 25227
rect 19884 25207 19886 25227
rect 19921 25222 19924 25227
rect 19932 25222 19934 25227
rect 19931 25208 19934 25222
rect 19956 25207 19958 25227
rect 19980 25207 19982 25227
rect 20028 25224 20030 25227
rect 20028 25207 20031 25224
rect 20052 25207 20054 25227
rect 20076 25207 20078 25227
rect 20124 25207 20126 25227
rect 20172 25207 20174 25227
rect 20196 25207 20198 25227
rect 20199 25224 20213 25227
rect 20223 25227 24779 25231
rect 20223 25224 20237 25227
rect 20268 25207 20270 25227
rect 20292 25207 20294 25227
rect 20388 25207 20390 25227
rect 20412 25207 20414 25227
rect 20508 25207 20510 25227
rect 20604 25207 20606 25227
rect 20964 25207 20966 25227
rect 21012 25207 21014 25227
rect 21108 25207 21110 25227
rect 21204 25207 21206 25227
rect 21300 25207 21302 25227
rect 21324 25207 21326 25227
rect 21444 25207 21446 25227
rect 21468 25207 21470 25227
rect 21564 25207 21566 25227
rect 21588 25207 21590 25227
rect 21684 25207 21686 25227
rect 21708 25207 21710 25227
rect 21828 25207 21830 25227
rect 21924 25207 21926 25227
rect 22068 25207 22070 25227
rect 22188 25207 22190 25227
rect 22212 25207 22214 25227
rect 22884 25207 22886 25227
rect 22980 25207 22982 25227
rect 23076 25207 23078 25227
rect 23100 25207 23102 25227
rect 23124 25207 23126 25227
rect 23244 25207 23246 25227
rect 23340 25207 23342 25227
rect 23412 25207 23414 25227
rect 23460 25207 23462 25227
rect 23508 25207 23510 25227
rect 23556 25207 23558 25227
rect 23604 25207 23606 25227
rect 23652 25207 23654 25227
rect 23676 25207 23678 25227
rect 23700 25207 23702 25227
rect 23772 25207 23774 25227
rect 23796 25207 23798 25227
rect 23916 25207 23918 25227
rect 24012 25207 24014 25227
rect 24060 25207 24062 25227
rect 24156 25207 24158 25227
rect 24492 25207 24494 25227
rect 24516 25207 24518 25227
rect 24588 25207 24590 25227
rect 24612 25207 24614 25227
rect 24684 25208 24686 25227
rect 24745 25222 24748 25227
rect 24756 25222 24758 25227
rect 24755 25208 24758 25222
rect 24649 25207 24707 25208
rect 24721 25207 24755 25208
rect -13895 25203 -5347 25207
rect -13788 25200 -13786 25203
rect -13788 25184 -13785 25200
rect -13799 25183 -13765 25184
rect -13428 25183 -13426 25203
rect -12852 25183 -12850 25203
rect -12767 25198 -12764 25203
rect -12756 25198 -12754 25203
rect -12757 25184 -12754 25198
rect -12636 25183 -12634 25203
rect -12156 25200 -12154 25203
rect -12156 25184 -12153 25200
rect -12311 25183 -12253 25184
rect -12191 25183 -12133 25184
rect -12060 25183 -12058 25203
rect -11772 25183 -11770 25203
rect -11676 25183 -11674 25203
rect -11652 25183 -11650 25203
rect -11508 25183 -11506 25203
rect -11436 25183 -11434 25203
rect -11412 25183 -11410 25203
rect -11340 25183 -11338 25203
rect -11196 25183 -11194 25203
rect -11100 25183 -11098 25203
rect -10764 25183 -10762 25203
rect -10644 25183 -10642 25203
rect -10017 25200 -10003 25203
rect -9996 25200 -9993 25203
rect -9900 25183 -9898 25203
rect -9732 25183 -9730 25203
rect -9444 25183 -9442 25203
rect -9348 25183 -9346 25203
rect -9228 25183 -9226 25203
rect -9108 25183 -9106 25203
rect -8436 25183 -8434 25203
rect -8364 25183 -8362 25203
rect -8340 25183 -8338 25203
rect -8268 25183 -8266 25203
rect -8004 25183 -8002 25203
rect -7932 25183 -7930 25203
rect -7524 25183 -7522 25203
rect -7356 25183 -7354 25203
rect -7308 25183 -7306 25203
rect -7212 25183 -7210 25203
rect -7044 25183 -7042 25203
rect -6948 25183 -6946 25203
rect -6852 25183 -6850 25203
rect -6756 25183 -6754 25203
rect -6660 25183 -6658 25203
rect -6612 25183 -6610 25203
rect -6516 25183 -6514 25203
rect -6372 25184 -6370 25203
rect -6479 25183 -6445 25184
rect -6383 25183 -6349 25184
rect -5892 25183 -5890 25203
rect -5436 25183 -5434 25203
rect -5361 25200 -5347 25203
rect -5340 25203 7397 25207
rect -5340 25200 -5323 25203
rect -5340 25183 -5338 25200
rect -5196 25183 -5194 25203
rect -5100 25183 -5098 25203
rect -4716 25183 -4714 25203
rect -4500 25183 -4498 25203
rect -4404 25183 -4402 25203
rect -4308 25183 -4306 25203
rect -4164 25183 -4162 25203
rect -4020 25183 -4018 25203
rect -3876 25183 -3874 25203
rect -3732 25183 -3730 25203
rect -3636 25183 -3634 25203
rect -3540 25183 -3538 25203
rect -3468 25183 -3466 25203
rect -3324 25183 -3322 25203
rect -3108 25183 -3106 25203
rect -3012 25183 -3010 25203
rect -2964 25183 -2962 25203
rect -2916 25183 -2914 25203
rect -2892 25183 -2890 25203
rect -2868 25183 -2866 25203
rect -2820 25183 -2818 25203
rect -2796 25184 -2794 25203
rect -2807 25183 -2773 25184
rect -2772 25183 -2770 25203
rect -2676 25183 -2674 25203
rect -2505 25200 -2491 25203
rect -2364 25183 -2362 25203
rect -2316 25183 -2314 25203
rect -2244 25184 -2242 25203
rect -2193 25200 -2179 25203
rect -2172 25200 -2169 25203
rect -2255 25183 -2221 25184
rect -2148 25183 -2146 25203
rect -2076 25183 -2074 25203
rect -2052 25183 -2050 25203
rect -1980 25183 -1978 25203
rect -1884 25183 -1882 25203
rect -1572 25183 -1570 25203
rect -1476 25183 -1474 25203
rect -1356 25183 -1354 25203
rect -1260 25183 -1258 25203
rect -1236 25183 -1234 25203
rect -1140 25183 -1138 25203
rect -876 25183 -874 25203
rect -660 25183 -658 25203
rect -537 25200 -523 25203
rect -492 25183 -490 25203
rect -444 25183 -442 25203
rect -396 25183 -394 25203
rect -348 25183 -346 25203
rect -276 25183 -274 25203
rect -225 25200 -211 25203
rect -12 25183 -10 25203
rect 156 25183 158 25203
rect 204 25183 206 25203
rect 252 25183 254 25203
rect 348 25183 350 25203
rect 468 25183 470 25203
rect 492 25183 494 25203
rect 564 25183 566 25203
rect 588 25183 590 25203
rect 636 25183 638 25203
rect 660 25183 662 25203
rect 732 25183 734 25203
rect 1092 25183 1094 25203
rect 1140 25183 1142 25203
rect 1236 25184 1238 25203
rect 1225 25183 1259 25184
rect 1308 25183 1310 25203
rect 1332 25183 1334 25203
rect 1380 25200 1382 25203
rect 1380 25183 1383 25200
rect 1428 25183 1430 25203
rect 1476 25183 1478 25203
rect 1692 25183 1694 25203
rect 1788 25184 1790 25203
rect 1753 25183 1811 25184
rect 2028 25183 2030 25203
rect 2076 25183 2078 25203
rect 2100 25183 2102 25203
rect 2124 25183 2126 25203
rect 2244 25183 2246 25203
rect 2412 25183 2414 25203
rect 2460 25183 2462 25203
rect 2508 25183 2510 25203
rect 2604 25183 2606 25203
rect 2772 25183 2774 25203
rect 2868 25183 2870 25203
rect 2940 25183 2942 25203
rect 3012 25183 3014 25203
rect 3108 25183 3110 25203
rect 3396 25183 3398 25203
rect 3564 25183 3566 25203
rect 3636 25183 3638 25203
rect 3660 25183 3662 25203
rect 3732 25183 3734 25203
rect 3780 25183 3782 25203
rect 3828 25183 3830 25203
rect 3924 25183 3926 25203
rect 4020 25183 4022 25203
rect 4092 25183 4094 25203
rect 4188 25183 4190 25203
rect 4308 25183 4310 25203
rect 4404 25183 4406 25203
rect 4500 25183 4502 25203
rect 4596 25183 4598 25203
rect 4692 25183 4694 25203
rect 4860 25183 4862 25203
rect 4956 25183 4958 25203
rect 4980 25183 4982 25203
rect 5052 25183 5054 25203
rect 5124 25183 5126 25203
rect 5220 25183 5222 25203
rect 5268 25183 5270 25203
rect 5388 25183 5390 25203
rect 5484 25183 5486 25203
rect 5508 25183 5510 25203
rect 5532 25183 5534 25203
rect 5628 25183 5630 25203
rect 5652 25183 5654 25203
rect 5748 25183 5750 25203
rect 5796 25183 5798 25203
rect 5844 25183 5846 25203
rect 5892 25183 5894 25203
rect 6132 25183 6134 25203
rect 6228 25183 6230 25203
rect 6252 25183 6254 25203
rect 6276 25183 6278 25203
rect 6324 25183 6326 25203
rect 6372 25183 6374 25203
rect 6420 25183 6422 25203
rect 6492 25183 6494 25203
rect 6516 25183 6518 25203
rect 6588 25183 6590 25203
rect 6612 25183 6614 25203
rect 6660 25183 6662 25203
rect 6684 25183 6686 25203
rect 6708 25183 6710 25203
rect 6780 25183 6782 25203
rect 6804 25183 6806 25203
rect 6900 25183 6902 25203
rect 6924 25183 6926 25203
rect 7020 25183 7022 25203
rect 7164 25183 7166 25203
rect 7236 25183 7238 25203
rect 7308 25183 7310 25203
rect 7380 25183 7382 25203
rect 7383 25200 7397 25203
rect 7407 25203 15965 25207
rect 7407 25200 7421 25203
rect 7428 25200 7431 25203
rect 7452 25183 7454 25203
rect 7476 25183 7478 25203
rect 7524 25183 7526 25203
rect 7548 25183 7550 25203
rect 7572 25183 7574 25203
rect 7620 25183 7622 25203
rect 7644 25183 7646 25203
rect 7668 25183 7670 25203
rect 7908 25183 7910 25203
rect 7956 25183 7958 25203
rect 8124 25183 8126 25203
rect 8209 25198 8212 25203
rect 8340 25200 8342 25203
rect 8219 25184 8222 25198
rect 8220 25183 8222 25184
rect 8340 25183 8343 25200
rect 8652 25183 8654 25203
rect 8700 25183 8702 25203
rect 8748 25183 8750 25203
rect 8820 25184 8822 25203
rect 8785 25183 8843 25184
rect 8844 25183 8846 25203
rect 8868 25183 8870 25203
rect 9516 25183 9518 25203
rect 9660 25183 9662 25203
rect 9684 25183 9686 25203
rect 9756 25183 9758 25203
rect 9780 25183 9782 25203
rect 9804 25183 9806 25203
rect 9852 25183 9854 25203
rect 9900 25183 9902 25203
rect 9948 25183 9950 25203
rect 10044 25183 10046 25203
rect 10116 25183 10118 25203
rect 10188 25183 10190 25203
rect 10212 25183 10214 25203
rect 10284 25183 10286 25203
rect 10332 25183 10334 25203
rect 10380 25183 10382 25203
rect 10428 25183 10430 25203
rect 10476 25183 10478 25203
rect 10500 25183 10502 25203
rect 10524 25183 10526 25203
rect 10572 25183 10574 25203
rect 10596 25183 10598 25203
rect 10620 25183 10622 25203
rect 10716 25183 10718 25203
rect 10956 25183 10958 25203
rect 11004 25183 11006 25203
rect 11052 25183 11054 25203
rect 11100 25183 11102 25203
rect 11172 25183 11174 25203
rect 11220 25183 11222 25203
rect 11340 25183 11342 25203
rect 11436 25183 11438 25203
rect 11532 25183 11534 25203
rect 11559 25200 11573 25203
rect 11580 25200 11583 25203
rect 11628 25183 11630 25203
rect 11676 25183 11678 25203
rect 11724 25183 11726 25203
rect 11772 25183 11774 25203
rect 11796 25183 11798 25203
rect 11892 25183 11894 25203
rect 11988 25183 11990 25203
rect 12060 25183 12062 25203
rect 12228 25183 12230 25203
rect 12276 25183 12278 25203
rect 12324 25183 12326 25203
rect 12420 25183 12422 25203
rect 12444 25183 12446 25203
rect 12481 25198 12484 25203
rect 12492 25198 12494 25203
rect 12491 25184 12494 25198
rect 12516 25183 12518 25203
rect 12540 25183 12542 25203
rect 12588 25200 12590 25203
rect 12588 25183 12591 25200
rect 12636 25183 12638 25203
rect 12732 25183 12734 25203
rect 12756 25183 12758 25203
rect 12804 25183 12806 25203
rect 12828 25183 12830 25203
rect 12972 25183 12974 25203
rect 13044 25183 13046 25203
rect 13068 25183 13070 25203
rect 13116 25183 13118 25203
rect 13284 25183 13286 25203
rect 13332 25183 13334 25203
rect 13572 25183 13574 25203
rect 13620 25183 13622 25203
rect 13668 25183 13670 25203
rect 13716 25183 13718 25203
rect 13764 25183 13766 25203
rect 13860 25183 13862 25203
rect 13956 25183 13958 25203
rect 14004 25183 14006 25203
rect 14100 25183 14102 25203
rect 14929 25183 14987 25184
rect 15180 25183 15182 25203
rect 15276 25183 15278 25203
rect 15420 25183 15422 25203
rect 15492 25183 15494 25203
rect 15660 25183 15662 25203
rect 15708 25183 15710 25203
rect 15732 25183 15734 25203
rect 15756 25183 15758 25203
rect 15804 25183 15806 25203
rect 15828 25183 15830 25203
rect 15852 25183 15854 25203
rect 15948 25183 15950 25203
rect 15951 25200 15965 25203
rect 15972 25203 19997 25207
rect 15972 25200 15989 25203
rect 15972 25183 15974 25200
rect 16044 25183 16046 25203
rect 16068 25183 16070 25203
rect 16164 25183 16166 25203
rect 16260 25183 16262 25203
rect 16332 25183 16334 25203
rect 16548 25183 16550 25203
rect 16572 25183 16574 25203
rect 16620 25183 16622 25203
rect 16668 25183 16670 25203
rect 16716 25183 16718 25203
rect 16764 25183 16766 25203
rect 16812 25183 16814 25203
rect 16884 25183 16886 25203
rect 16908 25183 16910 25203
rect 16980 25183 16982 25203
rect 17148 25183 17150 25203
rect 17196 25183 17198 25203
rect 17220 25183 17222 25203
rect 17292 25183 17294 25203
rect 17316 25183 17318 25203
rect 18132 25183 18134 25203
rect 18228 25183 18230 25203
rect 18492 25183 18494 25203
rect 18516 25183 18518 25203
rect 18564 25183 18566 25203
rect 18612 25183 18614 25203
rect 18660 25183 18662 25203
rect 18756 25183 18758 25203
rect 18900 25183 18902 25203
rect 18924 25183 18926 25203
rect 18996 25183 18998 25203
rect 19020 25183 19022 25203
rect 19092 25183 19094 25203
rect 19140 25183 19142 25203
rect 19188 25184 19190 25203
rect 19153 25183 19211 25184
rect 19236 25183 19238 25203
rect 19788 25183 19790 25203
rect 19836 25183 19838 25203
rect 19860 25183 19862 25203
rect 19884 25183 19886 25203
rect 19956 25183 19958 25203
rect 19980 25183 19982 25203
rect 19983 25200 19997 25203
rect 20007 25203 24755 25207
rect 20007 25200 20021 25203
rect 20028 25200 20031 25203
rect 20052 25183 20054 25203
rect 20076 25183 20078 25203
rect 20124 25183 20126 25203
rect 20172 25183 20174 25203
rect 20196 25183 20198 25203
rect 20268 25183 20270 25203
rect 20292 25183 20294 25203
rect 20388 25183 20390 25203
rect 20412 25183 20414 25203
rect 20508 25183 20510 25203
rect 20604 25183 20606 25203
rect 20964 25183 20966 25203
rect 21012 25183 21014 25203
rect 21108 25183 21110 25203
rect 21204 25183 21206 25203
rect 21300 25183 21302 25203
rect 21324 25183 21326 25203
rect 21444 25183 21446 25203
rect 21468 25183 21470 25203
rect 21564 25183 21566 25203
rect 21588 25183 21590 25203
rect 21684 25183 21686 25203
rect 21708 25183 21710 25203
rect 21828 25183 21830 25203
rect 21924 25183 21926 25203
rect 22068 25183 22070 25203
rect 22188 25183 22190 25203
rect 22212 25183 22214 25203
rect 22884 25183 22886 25203
rect 22980 25183 22982 25203
rect 23076 25183 23078 25203
rect 23100 25183 23102 25203
rect 23124 25183 23126 25203
rect 23244 25183 23246 25203
rect 23340 25183 23342 25203
rect 23412 25183 23414 25203
rect 23460 25183 23462 25203
rect 23508 25183 23510 25203
rect 23556 25183 23558 25203
rect 23604 25183 23606 25203
rect 23652 25183 23654 25203
rect 23676 25183 23678 25203
rect 23700 25183 23702 25203
rect 23772 25183 23774 25203
rect 23796 25183 23798 25203
rect 23916 25183 23918 25203
rect 24012 25183 24014 25203
rect 24060 25183 24062 25203
rect 24156 25183 24158 25203
rect 24492 25183 24494 25203
rect 24516 25183 24518 25203
rect 24588 25183 24590 25203
rect 24612 25184 24614 25203
rect 24673 25198 24676 25203
rect 24684 25198 24686 25203
rect 24683 25184 24686 25198
rect 24745 25190 24749 25198
rect 24735 25184 24745 25190
rect 24601 25183 24635 25184
rect -13799 25179 1349 25183
rect -13799 25176 -13795 25179
rect -13788 25176 -13785 25179
rect -13679 25159 -13645 25160
rect -13428 25159 -13426 25179
rect -12852 25159 -12850 25179
rect -12681 25176 -12667 25179
rect -12636 25159 -12634 25179
rect -12311 25174 -12308 25179
rect -12191 25174 -12188 25179
rect -12177 25176 -12163 25179
rect -12156 25176 -12153 25179
rect -12060 25176 -12058 25179
rect -12301 25160 -12298 25174
rect -12181 25160 -12177 25174
rect -12300 25159 -12298 25160
rect -12180 25159 -12177 25160
rect -12060 25159 -12057 25176
rect -11772 25159 -11770 25179
rect -11676 25159 -11674 25179
rect -11652 25159 -11650 25179
rect -11508 25159 -11506 25179
rect -11436 25159 -11434 25179
rect -11412 25159 -11410 25179
rect -11340 25159 -11338 25179
rect -11196 25159 -11194 25179
rect -11100 25159 -11098 25179
rect -10764 25159 -10762 25179
rect -10644 25159 -10642 25179
rect -9959 25159 -9925 25160
rect -9900 25159 -9898 25179
rect -9732 25159 -9730 25179
rect -9444 25159 -9442 25179
rect -9348 25159 -9346 25179
rect -9228 25159 -9226 25179
rect -9108 25159 -9106 25179
rect -8436 25159 -8434 25179
rect -8364 25159 -8362 25179
rect -8340 25159 -8338 25179
rect -8268 25159 -8266 25179
rect -8004 25159 -8002 25179
rect -7932 25159 -7930 25179
rect -7524 25159 -7522 25179
rect -7356 25159 -7354 25179
rect -7308 25159 -7306 25179
rect -7212 25159 -7210 25179
rect -7044 25159 -7042 25179
rect -6948 25159 -6946 25179
rect -6852 25159 -6850 25179
rect -6756 25159 -6754 25179
rect -6660 25159 -6658 25179
rect -6612 25159 -6610 25179
rect -6516 25159 -6514 25179
rect -6383 25174 -6380 25179
rect -6372 25176 -6370 25179
rect -5985 25176 -5971 25179
rect -6372 25174 -6369 25176
rect -6373 25160 -6369 25174
rect -5892 25159 -5890 25179
rect -5436 25159 -5434 25179
rect -5340 25159 -5338 25179
rect -5196 25159 -5194 25179
rect -5100 25159 -5098 25179
rect -4716 25159 -4714 25179
rect -4500 25159 -4498 25179
rect -4404 25159 -4402 25179
rect -4343 25159 -4309 25160
rect -4308 25159 -4306 25179
rect -4164 25159 -4162 25179
rect -4020 25159 -4018 25179
rect -3876 25159 -3874 25179
rect -3732 25159 -3730 25179
rect -3636 25159 -3634 25179
rect -3540 25159 -3538 25179
rect -3468 25159 -3466 25179
rect -3324 25159 -3322 25179
rect -3108 25159 -3106 25179
rect -3012 25159 -3010 25179
rect -2964 25159 -2962 25179
rect -2916 25159 -2914 25179
rect -2892 25159 -2890 25179
rect -2868 25159 -2866 25179
rect -2820 25159 -2818 25179
rect -2807 25174 -2804 25179
rect -2796 25174 -2794 25179
rect -2797 25160 -2794 25174
rect -2772 25159 -2770 25179
rect -2676 25159 -2674 25179
rect -2364 25159 -2362 25179
rect -2316 25159 -2314 25179
rect -2255 25174 -2252 25179
rect -2244 25174 -2242 25179
rect -2245 25160 -2242 25174
rect -2148 25176 -2146 25179
rect -2148 25159 -2145 25176
rect -2076 25159 -2074 25179
rect -2052 25159 -2050 25179
rect -1980 25159 -1978 25179
rect -1884 25159 -1882 25179
rect -1572 25159 -1570 25179
rect -1476 25159 -1474 25179
rect -1356 25159 -1354 25179
rect -1260 25159 -1258 25179
rect -1236 25159 -1234 25179
rect -1140 25159 -1138 25179
rect -876 25159 -874 25179
rect -660 25159 -658 25179
rect -492 25159 -490 25179
rect -444 25159 -442 25179
rect -396 25159 -394 25179
rect -348 25159 -346 25179
rect -276 25159 -274 25179
rect -12 25159 -10 25179
rect 156 25159 158 25179
rect 204 25159 206 25179
rect 252 25159 254 25179
rect 348 25159 350 25179
rect 468 25159 470 25179
rect 492 25159 494 25179
rect 564 25159 566 25179
rect 588 25159 590 25179
rect 636 25159 638 25179
rect 660 25159 662 25179
rect 732 25159 734 25179
rect 1092 25159 1094 25179
rect 1140 25159 1142 25179
rect 1225 25174 1228 25179
rect 1236 25174 1238 25179
rect 1235 25160 1238 25174
rect 1308 25159 1310 25179
rect 1332 25176 1334 25179
rect 1335 25176 1349 25179
rect 1359 25179 8309 25183
rect 1359 25176 1373 25179
rect 1380 25176 1383 25179
rect 1332 25159 1335 25176
rect 1428 25159 1430 25179
rect 1476 25159 1478 25179
rect 1692 25159 1694 25179
rect 1777 25174 1780 25179
rect 1788 25174 1790 25179
rect 1787 25160 1790 25174
rect 1860 25159 1863 25176
rect 2028 25159 2030 25179
rect 2076 25159 2078 25179
rect 2100 25159 2102 25179
rect 2124 25159 2126 25179
rect 2244 25159 2246 25179
rect 2412 25159 2414 25179
rect 2460 25159 2462 25179
rect 2508 25159 2510 25179
rect 2604 25159 2606 25179
rect 2772 25159 2774 25179
rect 2868 25159 2870 25179
rect 2940 25159 2942 25179
rect 3012 25159 3014 25179
rect 3108 25159 3110 25179
rect 3217 25159 3275 25160
rect 3396 25159 3398 25179
rect 3564 25159 3566 25179
rect 3636 25159 3638 25179
rect 3660 25159 3662 25179
rect 3732 25159 3734 25179
rect 3780 25159 3782 25179
rect 3828 25159 3830 25179
rect 3924 25159 3926 25179
rect 4020 25159 4022 25179
rect 4092 25159 4094 25179
rect 4188 25159 4190 25179
rect 4308 25159 4310 25179
rect 4404 25159 4406 25179
rect 4500 25159 4502 25179
rect 4596 25159 4598 25179
rect 4692 25159 4694 25179
rect 4719 25176 4733 25179
rect 4860 25159 4862 25179
rect 4956 25159 4958 25179
rect 4980 25159 4982 25179
rect 5052 25159 5054 25179
rect 5124 25159 5126 25179
rect 5220 25159 5222 25179
rect 5268 25159 5270 25179
rect 5388 25159 5390 25179
rect 5484 25159 5486 25179
rect 5508 25159 5510 25179
rect 5532 25159 5534 25179
rect 5628 25159 5630 25179
rect 5652 25159 5654 25179
rect 5748 25159 5750 25179
rect 5796 25159 5798 25179
rect 5844 25159 5846 25179
rect 5892 25159 5894 25179
rect 6132 25159 6134 25179
rect 6228 25159 6230 25179
rect 6252 25159 6254 25179
rect 6276 25159 6278 25179
rect 6324 25159 6326 25179
rect 6372 25159 6374 25179
rect 6420 25159 6422 25179
rect 6492 25159 6494 25179
rect 6516 25159 6518 25179
rect 6588 25159 6590 25179
rect 6612 25159 6614 25179
rect 6660 25159 6662 25179
rect 6684 25159 6686 25179
rect 6708 25159 6710 25179
rect 6780 25159 6782 25179
rect 6804 25159 6806 25179
rect 6900 25159 6902 25179
rect 6924 25159 6926 25179
rect 7020 25159 7022 25179
rect 7164 25159 7166 25179
rect 7236 25159 7238 25179
rect 7308 25159 7310 25179
rect 7380 25159 7382 25179
rect 7452 25159 7454 25179
rect 7476 25159 7478 25179
rect 7524 25159 7526 25179
rect 7548 25159 7550 25179
rect 7572 25159 7574 25179
rect 7620 25159 7622 25179
rect 7644 25159 7646 25179
rect 7668 25159 7670 25179
rect 7908 25159 7910 25179
rect 7956 25159 7958 25179
rect 8124 25159 8126 25179
rect 8220 25159 8222 25179
rect 8295 25176 8309 25179
rect 8319 25179 12557 25183
rect 8319 25176 8333 25179
rect 8340 25176 8343 25179
rect 8652 25159 8654 25179
rect 8700 25159 8702 25179
rect 8748 25159 8750 25179
rect 8785 25174 8788 25179
rect 8809 25174 8812 25179
rect 8820 25174 8822 25179
rect 8795 25160 8798 25174
rect 8819 25160 8822 25174
rect 8796 25159 8798 25160
rect 8844 25159 8846 25179
rect 8868 25159 8870 25179
rect 9516 25159 9518 25179
rect 9660 25159 9662 25179
rect 9684 25159 9686 25179
rect 9756 25159 9758 25179
rect 9780 25159 9782 25179
rect 9804 25159 9806 25179
rect 9852 25159 9854 25179
rect 9900 25159 9902 25179
rect 9948 25159 9950 25179
rect 10044 25159 10046 25179
rect 10116 25159 10118 25179
rect 10188 25159 10190 25179
rect 10212 25160 10214 25179
rect 10201 25159 10235 25160
rect 10284 25159 10286 25179
rect 10332 25159 10334 25179
rect 10380 25159 10382 25179
rect 10428 25159 10430 25179
rect 10476 25159 10478 25179
rect 10500 25159 10502 25179
rect 10524 25159 10526 25179
rect 10572 25160 10574 25179
rect 10537 25159 10595 25160
rect 10596 25159 10598 25179
rect 10620 25159 10622 25179
rect 10716 25159 10718 25179
rect 10956 25159 10958 25179
rect 11004 25159 11006 25179
rect 11052 25159 11054 25179
rect 11100 25159 11102 25179
rect 11172 25159 11174 25179
rect 11220 25159 11222 25179
rect 11340 25159 11342 25179
rect 11436 25159 11438 25179
rect 11532 25159 11534 25179
rect 11628 25159 11630 25179
rect 11676 25159 11678 25179
rect 11724 25159 11726 25179
rect 11772 25159 11774 25179
rect 11796 25159 11798 25179
rect 11892 25159 11894 25179
rect 11988 25159 11990 25179
rect 12060 25159 12062 25179
rect 12228 25159 12230 25179
rect 12276 25159 12278 25179
rect 12324 25159 12326 25179
rect 12420 25159 12422 25179
rect 12444 25159 12446 25179
rect 12516 25159 12518 25179
rect 12540 25159 12542 25179
rect 12543 25176 12557 25179
rect 12567 25179 24635 25183
rect 12567 25176 12581 25179
rect 12588 25176 12591 25179
rect 12636 25159 12638 25179
rect 12732 25159 12734 25179
rect 12756 25159 12758 25179
rect 12804 25159 12806 25179
rect 12828 25159 12830 25179
rect 12972 25159 12974 25179
rect 13044 25159 13046 25179
rect 13068 25159 13070 25179
rect 13116 25159 13118 25179
rect 13284 25159 13286 25179
rect 13332 25159 13334 25179
rect 13572 25159 13574 25179
rect 13620 25159 13622 25179
rect 13668 25159 13670 25179
rect 13716 25159 13718 25179
rect 13764 25159 13766 25179
rect 13860 25159 13862 25179
rect 13956 25159 13958 25179
rect 14004 25159 14006 25179
rect 14100 25159 14102 25179
rect 14929 25174 14932 25179
rect 14939 25160 14942 25174
rect 14940 25159 14942 25160
rect 15036 25159 15039 25176
rect 15180 25159 15182 25179
rect 15276 25159 15278 25179
rect 15420 25159 15422 25179
rect 15492 25159 15494 25179
rect 15660 25159 15662 25179
rect 15708 25159 15710 25179
rect 15732 25159 15734 25179
rect 15756 25159 15758 25179
rect 15804 25159 15806 25179
rect 15828 25159 15830 25179
rect 15852 25159 15854 25179
rect 15948 25159 15950 25179
rect 15972 25159 15974 25179
rect 16044 25159 16046 25179
rect 16068 25159 16070 25179
rect 16164 25159 16166 25179
rect 16260 25159 16262 25179
rect 16332 25159 16334 25179
rect 16548 25159 16550 25179
rect 16572 25159 16574 25179
rect 16620 25159 16622 25179
rect 16668 25159 16670 25179
rect 16716 25159 16718 25179
rect 16764 25159 16766 25179
rect 16812 25159 16814 25179
rect 16884 25159 16886 25179
rect 16908 25159 16910 25179
rect 16980 25159 16982 25179
rect 17148 25159 17150 25179
rect 17196 25159 17198 25179
rect 17220 25159 17222 25179
rect 17292 25159 17294 25179
rect 17316 25159 17318 25179
rect 18132 25159 18134 25179
rect 18228 25159 18230 25179
rect 18492 25159 18494 25179
rect 18516 25159 18518 25179
rect 18564 25159 18566 25179
rect 18612 25159 18614 25179
rect 18660 25159 18662 25179
rect 18756 25159 18758 25179
rect 18900 25159 18902 25179
rect 18924 25159 18926 25179
rect 18996 25159 18998 25179
rect 19020 25159 19022 25179
rect 19092 25159 19094 25179
rect 19140 25159 19142 25179
rect 19177 25174 19180 25179
rect 19188 25174 19190 25179
rect 19187 25160 19190 25174
rect 19236 25159 19238 25179
rect 19260 25159 19263 25176
rect 19788 25159 19790 25179
rect 19836 25159 19838 25179
rect 19860 25159 19862 25179
rect 19884 25159 19886 25179
rect 19956 25159 19958 25179
rect 19980 25159 19982 25179
rect 20052 25159 20054 25179
rect 20076 25159 20078 25179
rect 20124 25159 20126 25179
rect 20172 25159 20174 25179
rect 20196 25159 20198 25179
rect 20268 25159 20270 25179
rect 20292 25159 20294 25179
rect 20388 25159 20390 25179
rect 20412 25159 20414 25179
rect 20508 25159 20510 25179
rect 20604 25159 20606 25179
rect 20964 25159 20966 25179
rect 21012 25159 21014 25179
rect 21108 25159 21110 25179
rect 21204 25159 21206 25179
rect 21300 25159 21302 25179
rect 21324 25159 21326 25179
rect 21444 25159 21446 25179
rect 21468 25159 21470 25179
rect 21564 25159 21566 25179
rect 21588 25159 21590 25179
rect 21684 25159 21686 25179
rect 21708 25159 21710 25179
rect 21828 25159 21830 25179
rect 21924 25159 21926 25179
rect 22068 25159 22070 25179
rect 22188 25159 22190 25179
rect 22212 25159 22214 25179
rect 22884 25159 22886 25179
rect 22980 25159 22982 25179
rect 23076 25159 23078 25179
rect 23100 25159 23102 25179
rect 23124 25159 23126 25179
rect 23244 25159 23246 25179
rect 23340 25159 23342 25179
rect 23412 25159 23414 25179
rect 23460 25159 23462 25179
rect 23508 25159 23510 25179
rect 23556 25159 23558 25179
rect 23604 25159 23606 25179
rect 23652 25159 23654 25179
rect 23676 25159 23678 25179
rect 23700 25159 23702 25179
rect 23772 25159 23774 25179
rect 23796 25159 23798 25179
rect 23916 25159 23918 25179
rect 24012 25159 24014 25179
rect 24060 25159 24062 25179
rect 24156 25159 24158 25179
rect 24492 25159 24494 25179
rect 24516 25159 24518 25179
rect 24588 25160 24590 25179
rect 24601 25174 24604 25179
rect 24612 25174 24614 25179
rect 24611 25160 24614 25174
rect 24577 25159 24611 25160
rect -13679 25155 -12211 25159
rect -13535 25135 -13501 25136
rect -13428 25135 -13426 25155
rect -12852 25135 -12850 25155
rect -12636 25135 -12634 25155
rect -12300 25135 -12298 25155
rect -12225 25152 -12211 25155
rect -12201 25155 -12091 25159
rect -12201 25152 -12187 25155
rect -12180 25152 -12177 25155
rect -12105 25152 -12091 25155
rect -12081 25155 1853 25159
rect -12081 25152 -12067 25155
rect -12060 25152 -12057 25155
rect -11772 25135 -11770 25155
rect -11676 25135 -11674 25155
rect -11652 25135 -11650 25155
rect -11508 25135 -11506 25155
rect -11436 25135 -11434 25155
rect -11412 25135 -11410 25155
rect -11340 25135 -11338 25155
rect -11196 25135 -11194 25155
rect -11100 25135 -11098 25155
rect -10764 25135 -10762 25155
rect -10644 25135 -10642 25155
rect -9900 25135 -9898 25155
rect -9732 25135 -9730 25155
rect -9444 25135 -9442 25155
rect -9348 25135 -9346 25155
rect -9228 25135 -9226 25155
rect -9108 25135 -9106 25155
rect -8436 25135 -8434 25155
rect -8364 25135 -8362 25155
rect -8340 25135 -8338 25155
rect -8268 25135 -8266 25155
rect -8004 25135 -8002 25155
rect -7932 25135 -7930 25155
rect -7524 25135 -7522 25155
rect -7356 25135 -7354 25155
rect -7308 25135 -7306 25155
rect -7212 25135 -7210 25155
rect -7044 25135 -7042 25155
rect -6948 25135 -6946 25155
rect -6852 25135 -6850 25155
rect -6756 25135 -6754 25155
rect -6660 25135 -6658 25155
rect -6612 25135 -6610 25155
rect -6516 25135 -6514 25155
rect -6393 25152 -6379 25155
rect -6297 25152 -6283 25155
rect -5892 25135 -5890 25155
rect -5436 25135 -5434 25155
rect -5340 25135 -5338 25155
rect -5196 25135 -5194 25155
rect -5100 25135 -5098 25155
rect -4716 25135 -4714 25155
rect -4500 25135 -4498 25155
rect -4404 25135 -4402 25155
rect -4308 25135 -4306 25155
rect -4164 25135 -4162 25155
rect -4020 25135 -4018 25155
rect -3876 25135 -3874 25155
rect -3732 25135 -3730 25155
rect -3636 25135 -3634 25155
rect -3540 25135 -3538 25155
rect -3468 25135 -3466 25155
rect -3324 25135 -3322 25155
rect -3108 25135 -3106 25155
rect -3012 25135 -3010 25155
rect -2964 25135 -2962 25155
rect -2916 25135 -2914 25155
rect -2892 25135 -2890 25155
rect -2868 25135 -2866 25155
rect -2820 25135 -2818 25155
rect -2772 25135 -2770 25155
rect -2721 25152 -2707 25155
rect -2676 25135 -2674 25155
rect -2364 25135 -2362 25155
rect -2316 25135 -2314 25155
rect -2169 25152 -2155 25155
rect -2148 25152 -2145 25155
rect -2076 25135 -2074 25155
rect -2052 25135 -2050 25155
rect -1980 25135 -1978 25155
rect -1884 25135 -1882 25155
rect -1572 25135 -1570 25155
rect -1476 25135 -1474 25155
rect -1356 25135 -1354 25155
rect -1260 25135 -1258 25155
rect -1236 25135 -1234 25155
rect -1140 25135 -1138 25155
rect -876 25135 -874 25155
rect -660 25135 -658 25155
rect -492 25135 -490 25155
rect -444 25135 -442 25155
rect -396 25135 -394 25155
rect -348 25135 -346 25155
rect -276 25135 -274 25155
rect -12 25135 -10 25155
rect 156 25135 158 25155
rect 204 25135 206 25155
rect 252 25135 254 25155
rect 348 25135 350 25155
rect 468 25135 470 25155
rect 492 25135 494 25155
rect 564 25135 566 25155
rect 588 25135 590 25155
rect 636 25135 638 25155
rect 660 25135 662 25155
rect 732 25135 734 25155
rect 1092 25135 1094 25155
rect 1140 25135 1142 25155
rect 1308 25135 1310 25155
rect 1311 25152 1325 25155
rect 1332 25152 1335 25155
rect 1428 25135 1430 25155
rect 1476 25135 1478 25155
rect 1692 25135 1694 25155
rect 1839 25152 1853 25155
rect 1860 25155 8885 25159
rect 1860 25152 1877 25155
rect 1860 25135 1862 25152
rect 2028 25135 2030 25155
rect 2076 25135 2078 25155
rect 2100 25135 2102 25155
rect 2124 25135 2126 25155
rect 2244 25135 2246 25155
rect 2412 25135 2414 25155
rect 2460 25135 2462 25155
rect 2508 25135 2510 25155
rect 2604 25135 2606 25155
rect 2772 25135 2774 25155
rect 2868 25135 2870 25155
rect 2940 25135 2942 25155
rect 3012 25135 3014 25155
rect 3108 25135 3110 25155
rect 3324 25135 3327 25152
rect 3396 25135 3398 25155
rect 3564 25135 3566 25155
rect 3636 25135 3638 25155
rect 3660 25135 3662 25155
rect 3732 25135 3734 25155
rect 3780 25135 3782 25155
rect 3828 25135 3830 25155
rect 3924 25135 3926 25155
rect 4020 25135 4022 25155
rect 4092 25135 4094 25155
rect 4188 25135 4190 25155
rect 4308 25135 4310 25155
rect 4404 25135 4406 25155
rect 4500 25135 4502 25155
rect 4596 25135 4598 25155
rect 4692 25135 4694 25155
rect 4860 25135 4862 25155
rect 4956 25135 4958 25155
rect 4980 25135 4982 25155
rect 5052 25135 5054 25155
rect 5124 25135 5126 25155
rect 5220 25135 5222 25155
rect 5268 25135 5270 25155
rect 5388 25135 5390 25155
rect 5484 25135 5486 25155
rect 5508 25135 5510 25155
rect 5532 25135 5534 25155
rect 5628 25135 5630 25155
rect 5652 25135 5654 25155
rect 5748 25135 5750 25155
rect 5796 25135 5798 25155
rect 5844 25135 5846 25155
rect 5892 25135 5894 25155
rect 6132 25135 6134 25155
rect 6228 25135 6230 25155
rect 6252 25135 6254 25155
rect 6276 25135 6278 25155
rect 6324 25135 6326 25155
rect 6372 25135 6374 25155
rect 6420 25135 6422 25155
rect 6492 25135 6494 25155
rect 6516 25135 6518 25155
rect 6588 25135 6590 25155
rect 6612 25135 6614 25155
rect 6660 25135 6662 25155
rect 6684 25135 6686 25155
rect 6708 25135 6710 25155
rect 6780 25135 6782 25155
rect 6804 25135 6806 25155
rect 6900 25135 6902 25155
rect 6924 25135 6926 25155
rect 7020 25135 7022 25155
rect 7164 25135 7166 25155
rect 7236 25135 7238 25155
rect 7308 25135 7310 25155
rect 7380 25135 7382 25155
rect 7452 25135 7454 25155
rect 7476 25135 7478 25155
rect 7524 25135 7526 25155
rect 7548 25135 7550 25155
rect 7572 25135 7574 25155
rect 7620 25135 7622 25155
rect 7644 25135 7646 25155
rect 7668 25135 7670 25155
rect 7908 25135 7910 25155
rect 7956 25135 7958 25155
rect 8124 25135 8126 25155
rect 8220 25135 8222 25155
rect 8652 25135 8654 25155
rect 8700 25135 8702 25155
rect 8748 25135 8750 25155
rect 8796 25135 8798 25155
rect 8844 25135 8846 25155
rect 8868 25135 8870 25155
rect 8871 25152 8885 25155
rect 8895 25155 15029 25159
rect 8895 25152 8909 25155
rect 9516 25135 9518 25155
rect 9660 25135 9662 25155
rect 9684 25135 9686 25155
rect 9756 25135 9758 25155
rect 9780 25135 9782 25155
rect 9804 25135 9806 25155
rect 9852 25135 9854 25155
rect 9900 25135 9902 25155
rect 9948 25135 9950 25155
rect 10044 25135 10046 25155
rect 10116 25135 10118 25155
rect 10188 25135 10190 25155
rect 10201 25150 10204 25155
rect 10212 25150 10214 25155
rect 10211 25136 10214 25150
rect 10284 25135 10286 25155
rect 10332 25135 10334 25155
rect 10380 25135 10382 25155
rect 10428 25135 10430 25155
rect 10476 25135 10478 25155
rect 10500 25135 10502 25155
rect 10524 25135 10526 25155
rect 10561 25150 10564 25155
rect 10572 25150 10574 25155
rect 10571 25136 10574 25150
rect 10596 25135 10598 25155
rect 10620 25135 10622 25155
rect 10644 25135 10647 25152
rect 10716 25135 10718 25155
rect 10956 25135 10958 25155
rect 11004 25135 11006 25155
rect 11052 25135 11054 25155
rect 11100 25135 11102 25155
rect 11172 25135 11174 25155
rect 11220 25135 11222 25155
rect 11340 25135 11342 25155
rect 11436 25135 11438 25155
rect 11532 25135 11534 25155
rect 11628 25135 11630 25155
rect 11676 25135 11678 25155
rect 11724 25135 11726 25155
rect 11772 25135 11774 25155
rect 11796 25135 11798 25155
rect 11892 25135 11894 25155
rect 11988 25135 11990 25155
rect 12060 25135 12062 25155
rect 12228 25135 12230 25155
rect 12276 25135 12278 25155
rect 12324 25135 12326 25155
rect 12420 25135 12422 25155
rect 12444 25135 12446 25155
rect 12516 25135 12518 25155
rect 12540 25135 12542 25155
rect 12636 25135 12638 25155
rect 12732 25135 12734 25155
rect 12756 25135 12758 25155
rect 12804 25135 12806 25155
rect 12828 25135 12830 25155
rect 12972 25135 12974 25155
rect 13044 25135 13046 25155
rect 13068 25135 13070 25155
rect 13116 25135 13118 25155
rect 13284 25135 13286 25155
rect 13332 25135 13334 25155
rect 13572 25135 13574 25155
rect 13620 25135 13622 25155
rect 13668 25135 13670 25155
rect 13716 25135 13718 25155
rect 13764 25135 13766 25155
rect 13860 25135 13862 25155
rect 13956 25135 13958 25155
rect 14004 25135 14006 25155
rect 14100 25135 14102 25155
rect 14940 25135 14942 25155
rect 15015 25152 15029 25155
rect 15036 25155 19253 25159
rect 15036 25152 15053 25155
rect 15036 25135 15038 25152
rect 15180 25135 15182 25155
rect 15276 25135 15278 25155
rect 15420 25135 15422 25155
rect 15492 25135 15494 25155
rect 15660 25135 15662 25155
rect 15708 25135 15710 25155
rect 15732 25135 15734 25155
rect 15756 25135 15758 25155
rect 15804 25135 15806 25155
rect 15828 25135 15830 25155
rect 15852 25135 15854 25155
rect 15948 25135 15950 25155
rect 15972 25135 15974 25155
rect 16044 25135 16046 25155
rect 16068 25135 16070 25155
rect 16164 25135 16166 25155
rect 16260 25135 16262 25155
rect 16332 25135 16334 25155
rect 16548 25135 16550 25155
rect 16572 25135 16574 25155
rect 16620 25135 16622 25155
rect 16668 25135 16670 25155
rect 16716 25135 16718 25155
rect 16764 25135 16766 25155
rect 16812 25135 16814 25155
rect 16884 25135 16886 25155
rect 16908 25135 16910 25155
rect 16980 25135 16982 25155
rect 17148 25135 17150 25155
rect 17196 25135 17198 25155
rect 17220 25135 17222 25155
rect 17292 25135 17294 25155
rect 17316 25135 17318 25155
rect 18132 25135 18134 25155
rect 18228 25135 18230 25155
rect 18492 25135 18494 25155
rect 18516 25135 18518 25155
rect 18564 25135 18566 25155
rect 18612 25135 18614 25155
rect 18660 25135 18662 25155
rect 18756 25135 18758 25155
rect 18900 25135 18902 25155
rect 18924 25135 18926 25155
rect 18996 25135 18998 25155
rect 19020 25135 19022 25155
rect 19092 25135 19094 25155
rect 19140 25135 19142 25155
rect 19236 25135 19238 25155
rect 19239 25152 19253 25155
rect 19260 25155 24611 25159
rect 19260 25152 19277 25155
rect 19260 25135 19262 25152
rect 19788 25135 19790 25155
rect 19836 25135 19838 25155
rect 19860 25135 19862 25155
rect 19884 25135 19886 25155
rect 19956 25135 19958 25155
rect 19980 25135 19982 25155
rect 20052 25135 20054 25155
rect 20076 25135 20078 25155
rect 20124 25135 20126 25155
rect 20172 25135 20174 25155
rect 20196 25135 20198 25155
rect 20268 25136 20270 25155
rect 20257 25135 20291 25136
rect 20292 25135 20294 25155
rect 20388 25135 20390 25155
rect 20412 25135 20414 25155
rect 20508 25135 20510 25155
rect 20521 25135 20579 25136
rect 20604 25135 20606 25155
rect 20964 25135 20966 25155
rect 21012 25135 21014 25155
rect 21108 25135 21110 25155
rect 21204 25135 21206 25155
rect 21300 25135 21302 25155
rect 21324 25135 21326 25155
rect 21444 25135 21446 25155
rect 21468 25135 21470 25155
rect 21564 25135 21566 25155
rect 21588 25135 21590 25155
rect 21684 25135 21686 25155
rect 21708 25135 21710 25155
rect 21828 25135 21830 25155
rect 21924 25135 21926 25155
rect 22068 25135 22070 25155
rect 22188 25135 22190 25155
rect 22212 25135 22214 25155
rect 22884 25135 22886 25155
rect 22980 25135 22982 25155
rect 23076 25135 23078 25155
rect 23100 25135 23102 25155
rect 23124 25135 23126 25155
rect 23244 25135 23246 25155
rect 23340 25135 23342 25155
rect 23412 25135 23414 25155
rect 23460 25135 23462 25155
rect 23508 25135 23510 25155
rect 23556 25135 23558 25155
rect 23604 25135 23606 25155
rect 23652 25135 23654 25155
rect 23676 25135 23678 25155
rect 23700 25135 23702 25155
rect 23772 25135 23774 25155
rect 23796 25135 23798 25155
rect 23916 25135 23918 25155
rect 24012 25135 24014 25155
rect 24060 25135 24062 25155
rect 24156 25135 24158 25155
rect 24492 25135 24494 25155
rect 24516 25136 24518 25155
rect 24577 25150 24580 25155
rect 24588 25150 24590 25155
rect 24587 25136 24590 25150
rect 24505 25135 24539 25136
rect -13535 25131 3317 25135
rect -13428 25128 -13426 25131
rect -13428 25112 -13425 25128
rect -13439 25111 -13405 25112
rect -12852 25111 -12850 25131
rect -12636 25111 -12634 25131
rect -12300 25111 -12298 25131
rect -11772 25111 -11770 25131
rect -11676 25111 -11674 25131
rect -11652 25111 -11650 25131
rect -11508 25111 -11506 25131
rect -11436 25111 -11434 25131
rect -11412 25111 -11410 25131
rect -11340 25111 -11338 25131
rect -11196 25111 -11194 25131
rect -11100 25111 -11098 25131
rect -10764 25111 -10762 25131
rect -10644 25111 -10642 25131
rect -9900 25111 -9898 25131
rect -9873 25128 -9859 25131
rect -9732 25111 -9730 25131
rect -9444 25111 -9442 25131
rect -9348 25111 -9346 25131
rect -9228 25111 -9226 25131
rect -9108 25111 -9106 25131
rect -8436 25111 -8434 25131
rect -8364 25111 -8362 25131
rect -8340 25111 -8338 25131
rect -8268 25111 -8266 25131
rect -8135 25111 -8077 25112
rect -8004 25111 -8002 25131
rect -7932 25111 -7930 25131
rect -7775 25111 -7717 25112
rect -7524 25111 -7522 25131
rect -7356 25111 -7354 25131
rect -7308 25111 -7306 25131
rect -7212 25111 -7210 25131
rect -7044 25111 -7042 25131
rect -6948 25111 -6946 25131
rect -6852 25111 -6850 25131
rect -6756 25111 -6754 25131
rect -6660 25111 -6658 25131
rect -6612 25111 -6610 25131
rect -6516 25111 -6514 25131
rect -5892 25111 -5890 25131
rect -5436 25111 -5434 25131
rect -5340 25111 -5338 25131
rect -5196 25111 -5194 25131
rect -5100 25111 -5098 25131
rect -4716 25111 -4714 25131
rect -4500 25111 -4498 25131
rect -4404 25111 -4402 25131
rect -4308 25111 -4306 25131
rect -4257 25128 -4243 25131
rect -4164 25111 -4162 25131
rect -4020 25111 -4018 25131
rect -3876 25111 -3874 25131
rect -3732 25111 -3730 25131
rect -3636 25111 -3634 25131
rect -3540 25111 -3538 25131
rect -3468 25111 -3466 25131
rect -3324 25111 -3322 25131
rect -3108 25111 -3106 25131
rect -3012 25111 -3010 25131
rect -2964 25111 -2962 25131
rect -2916 25111 -2914 25131
rect -2892 25111 -2890 25131
rect -2868 25111 -2866 25131
rect -2820 25111 -2818 25131
rect -2772 25111 -2770 25131
rect -2676 25111 -2674 25131
rect -2364 25111 -2362 25131
rect -2316 25111 -2314 25131
rect -2076 25111 -2074 25131
rect -2052 25111 -2050 25131
rect -1980 25111 -1978 25131
rect -1884 25111 -1882 25131
rect -1572 25111 -1570 25131
rect -1476 25111 -1474 25131
rect -1356 25111 -1354 25131
rect -1260 25111 -1258 25131
rect -1236 25111 -1234 25131
rect -1140 25111 -1138 25131
rect -876 25111 -874 25131
rect -660 25111 -658 25131
rect -492 25111 -490 25131
rect -444 25111 -442 25131
rect -396 25111 -394 25131
rect -348 25111 -346 25131
rect -276 25111 -274 25131
rect -12 25111 -10 25131
rect 156 25111 158 25131
rect 204 25111 206 25131
rect 252 25111 254 25131
rect 348 25111 350 25131
rect 468 25111 470 25131
rect 492 25111 494 25131
rect 564 25111 566 25131
rect 588 25111 590 25131
rect 636 25111 638 25131
rect 660 25111 662 25131
rect 732 25111 734 25131
rect 1092 25111 1094 25131
rect 1140 25111 1142 25131
rect 1308 25111 1310 25131
rect 1345 25111 1403 25112
rect 1428 25111 1430 25131
rect 1476 25111 1478 25131
rect 1692 25111 1694 25131
rect 1860 25111 1862 25131
rect 2028 25111 2030 25131
rect 2076 25111 2078 25131
rect 2100 25111 2102 25131
rect 2124 25111 2126 25131
rect 2244 25111 2246 25131
rect 2412 25111 2414 25131
rect 2460 25111 2462 25131
rect 2508 25111 2510 25131
rect 2604 25111 2606 25131
rect 2772 25111 2774 25131
rect 2868 25111 2870 25131
rect 2940 25111 2942 25131
rect 3012 25111 3014 25131
rect 3108 25111 3110 25131
rect 3303 25128 3317 25131
rect 3324 25131 10637 25135
rect 3324 25128 3341 25131
rect 3324 25111 3326 25128
rect 3396 25111 3398 25131
rect 3564 25111 3566 25131
rect 3636 25111 3638 25131
rect 3660 25111 3662 25131
rect 3732 25111 3734 25131
rect 3780 25111 3782 25131
rect 3828 25111 3830 25131
rect 3924 25111 3926 25131
rect 4020 25111 4022 25131
rect 4092 25111 4094 25131
rect 4188 25111 4190 25131
rect 4308 25111 4310 25131
rect 4404 25111 4406 25131
rect 4500 25111 4502 25131
rect 4596 25111 4598 25131
rect 4692 25111 4694 25131
rect 4753 25111 4787 25112
rect 4860 25111 4862 25131
rect 4956 25111 4958 25131
rect 4980 25111 4982 25131
rect 5052 25111 5054 25131
rect 5124 25111 5126 25131
rect 5220 25111 5222 25131
rect 5268 25111 5270 25131
rect 5388 25111 5390 25131
rect 5484 25111 5486 25131
rect 5508 25111 5510 25131
rect 5532 25111 5534 25131
rect 5628 25111 5630 25131
rect 5652 25111 5654 25131
rect 5748 25111 5750 25131
rect 5796 25111 5798 25131
rect 5844 25111 5846 25131
rect 5892 25111 5894 25131
rect 6132 25111 6134 25131
rect 6228 25111 6230 25131
rect 6252 25111 6254 25131
rect 6276 25111 6278 25131
rect 6324 25111 6326 25131
rect 6372 25111 6374 25131
rect 6420 25111 6422 25131
rect 6492 25111 6494 25131
rect 6516 25111 6518 25131
rect 6588 25111 6590 25131
rect 6612 25111 6614 25131
rect 6660 25111 6662 25131
rect 6684 25111 6686 25131
rect 6708 25111 6710 25131
rect 6780 25111 6782 25131
rect 6804 25111 6806 25131
rect 6900 25111 6902 25131
rect 6924 25111 6926 25131
rect 7020 25111 7022 25131
rect 7164 25111 7166 25131
rect 7236 25111 7238 25131
rect 7308 25111 7310 25131
rect 7380 25111 7382 25131
rect 7393 25111 7451 25112
rect 7452 25111 7454 25131
rect 7476 25111 7478 25131
rect 7524 25111 7526 25131
rect 7548 25111 7550 25131
rect 7572 25111 7574 25131
rect 7620 25111 7622 25131
rect 7644 25111 7646 25131
rect 7668 25111 7670 25131
rect 7908 25111 7910 25131
rect 7956 25111 7958 25131
rect 8124 25111 8126 25131
rect 8220 25111 8222 25131
rect 8652 25111 8654 25131
rect 8700 25111 8702 25131
rect 8748 25111 8750 25131
rect 8796 25111 8798 25131
rect 8844 25111 8846 25131
rect 8868 25111 8870 25131
rect 9516 25111 9518 25131
rect 9660 25111 9662 25131
rect 9684 25111 9686 25131
rect 9756 25111 9758 25131
rect 9780 25111 9782 25131
rect 9804 25111 9806 25131
rect 9852 25111 9854 25131
rect 9900 25111 9902 25131
rect 9948 25111 9950 25131
rect 10044 25111 10046 25131
rect 10116 25111 10118 25131
rect 10188 25111 10190 25131
rect 10284 25111 10286 25131
rect 10287 25128 10301 25131
rect 10332 25111 10334 25131
rect 10380 25111 10382 25131
rect 10428 25111 10430 25131
rect 10476 25111 10478 25131
rect 10500 25111 10502 25131
rect 10524 25111 10526 25131
rect 10596 25111 10598 25131
rect 10620 25111 10622 25131
rect 10623 25128 10637 25131
rect 10644 25131 24539 25135
rect 10644 25128 10661 25131
rect 10644 25111 10646 25128
rect 10716 25111 10718 25131
rect 10956 25111 10958 25131
rect 11004 25111 11006 25131
rect 11052 25111 11054 25131
rect 11100 25111 11102 25131
rect 11172 25111 11174 25131
rect 11220 25111 11222 25131
rect 11340 25111 11342 25131
rect 11436 25111 11438 25131
rect 11532 25111 11534 25131
rect 11628 25111 11630 25131
rect 11676 25111 11678 25131
rect 11724 25111 11726 25131
rect 11772 25111 11774 25131
rect 11796 25111 11798 25131
rect 11892 25111 11894 25131
rect 11988 25111 11990 25131
rect 12060 25111 12062 25131
rect 12228 25111 12230 25131
rect 12276 25111 12278 25131
rect 12324 25111 12326 25131
rect 12420 25111 12422 25131
rect 12444 25111 12446 25131
rect 12516 25111 12518 25131
rect 12540 25111 12542 25131
rect 12636 25111 12638 25131
rect 12732 25111 12734 25131
rect 12756 25111 12758 25131
rect 12804 25111 12806 25131
rect 12828 25111 12830 25131
rect 12972 25111 12974 25131
rect 13044 25111 13046 25131
rect 13068 25111 13070 25131
rect 13116 25111 13118 25131
rect 13284 25111 13286 25131
rect 13332 25111 13334 25131
rect 13572 25111 13574 25131
rect 13620 25111 13622 25131
rect 13668 25111 13670 25131
rect 13716 25111 13718 25131
rect 13764 25111 13766 25131
rect 13860 25111 13862 25131
rect 13956 25111 13958 25131
rect 14004 25111 14006 25131
rect 14100 25111 14102 25131
rect 14940 25111 14942 25131
rect 15036 25111 15038 25131
rect 15180 25111 15182 25131
rect 15276 25111 15278 25131
rect 15420 25111 15422 25131
rect 15492 25111 15494 25131
rect 15660 25111 15662 25131
rect 15708 25111 15710 25131
rect 15732 25111 15734 25131
rect 15756 25111 15758 25131
rect 15804 25111 15806 25131
rect 15828 25111 15830 25131
rect 15852 25111 15854 25131
rect 15948 25111 15950 25131
rect 15972 25111 15974 25131
rect 16044 25111 16046 25131
rect 16068 25111 16070 25131
rect 16164 25111 16166 25131
rect 16260 25111 16262 25131
rect 16332 25111 16334 25131
rect 16548 25111 16550 25131
rect 16572 25111 16574 25131
rect 16620 25111 16622 25131
rect 16668 25111 16670 25131
rect 16716 25111 16718 25131
rect 16764 25111 16766 25131
rect 16812 25111 16814 25131
rect 16884 25111 16886 25131
rect 16908 25111 16910 25131
rect 16980 25111 16982 25131
rect 17148 25111 17150 25131
rect 17196 25111 17198 25131
rect 17220 25111 17222 25131
rect 17292 25111 17294 25131
rect 17316 25111 17318 25131
rect 18132 25111 18134 25131
rect 18228 25111 18230 25131
rect 18492 25111 18494 25131
rect 18516 25111 18518 25131
rect 18564 25111 18566 25131
rect 18612 25111 18614 25131
rect 18660 25111 18662 25131
rect 18756 25112 18758 25131
rect 18721 25111 18779 25112
rect 18900 25111 18902 25131
rect 18924 25111 18926 25131
rect 18996 25111 18998 25131
rect 19020 25111 19022 25131
rect 19092 25111 19094 25131
rect 19140 25111 19142 25131
rect 19236 25111 19238 25131
rect 19260 25111 19262 25131
rect 19788 25111 19790 25131
rect 19836 25111 19838 25131
rect 19860 25111 19862 25131
rect 19884 25111 19886 25131
rect 19956 25111 19958 25131
rect 19980 25111 19982 25131
rect 20052 25111 20054 25131
rect 20076 25111 20078 25131
rect 20124 25111 20126 25131
rect 20172 25111 20174 25131
rect 20196 25111 20198 25131
rect 20257 25126 20260 25131
rect 20268 25126 20270 25131
rect 20267 25112 20270 25126
rect 20292 25111 20294 25131
rect 20388 25111 20390 25131
rect 20412 25111 20414 25131
rect 20508 25111 20510 25131
rect 20521 25126 20524 25131
rect 20531 25112 20534 25126
rect 20532 25111 20534 25112
rect 20604 25111 20606 25131
rect 20628 25111 20631 25128
rect 20964 25111 20966 25131
rect 21012 25111 21014 25131
rect 21108 25111 21110 25131
rect 21204 25111 21206 25131
rect 21300 25111 21302 25131
rect 21324 25111 21326 25131
rect 21444 25111 21446 25131
rect 21468 25111 21470 25131
rect 21564 25111 21566 25131
rect 21588 25111 21590 25131
rect 21684 25111 21686 25131
rect 21708 25111 21710 25131
rect 21828 25111 21830 25131
rect 21924 25111 21926 25131
rect 22068 25111 22070 25131
rect 22188 25111 22190 25131
rect 22212 25111 22214 25131
rect 22884 25111 22886 25131
rect 22980 25111 22982 25131
rect 23076 25111 23078 25131
rect 23100 25111 23102 25131
rect 23124 25111 23126 25131
rect 23244 25111 23246 25131
rect 23340 25111 23342 25131
rect 23412 25111 23414 25131
rect 23460 25111 23462 25131
rect 23508 25111 23510 25131
rect 23556 25111 23558 25131
rect 23604 25111 23606 25131
rect 23652 25111 23654 25131
rect 23676 25111 23678 25131
rect 23700 25111 23702 25131
rect 23772 25111 23774 25131
rect 23796 25111 23798 25131
rect 23916 25111 23918 25131
rect 24012 25111 24014 25131
rect 24060 25111 24062 25131
rect 24156 25111 24158 25131
rect 24492 25112 24494 25131
rect 24505 25126 24508 25131
rect 24516 25126 24518 25131
rect 24515 25112 24518 25126
rect 24385 25111 24419 25112
rect 24481 25111 24515 25112
rect -13439 25107 20621 25111
rect -13439 25104 -13435 25107
rect -13428 25104 -13425 25107
rect -13319 25087 -13285 25088
rect -12852 25087 -12850 25107
rect -12636 25087 -12634 25107
rect -12300 25087 -12298 25107
rect -11772 25087 -11770 25107
rect -11676 25087 -11674 25107
rect -11652 25087 -11650 25107
rect -11508 25087 -11506 25107
rect -11436 25087 -11434 25107
rect -11412 25087 -11410 25107
rect -11340 25088 -11338 25107
rect -11351 25087 -11317 25088
rect -11196 25087 -11194 25107
rect -11100 25087 -11098 25107
rect -10764 25087 -10762 25107
rect -10644 25087 -10642 25107
rect -9900 25087 -9898 25107
rect -9791 25087 -9733 25088
rect -9732 25087 -9730 25107
rect -9444 25087 -9442 25107
rect -9348 25087 -9346 25107
rect -9228 25087 -9226 25107
rect -9108 25087 -9106 25107
rect -8436 25087 -8434 25107
rect -8364 25087 -8362 25107
rect -8340 25087 -8338 25107
rect -8268 25087 -8266 25107
rect -8135 25102 -8132 25107
rect -8004 25104 -8002 25107
rect -8125 25088 -8122 25102
rect -8124 25087 -8122 25088
rect -8028 25087 -8025 25104
rect -8004 25087 -8001 25104
rect -7932 25087 -7930 25107
rect -7775 25102 -7772 25107
rect -7765 25088 -7762 25102
rect -7764 25087 -7762 25088
rect -7524 25087 -7522 25107
rect -7356 25087 -7354 25107
rect -7308 25087 -7306 25107
rect -7212 25087 -7210 25107
rect -7044 25087 -7042 25107
rect -6948 25087 -6946 25107
rect -6852 25087 -6850 25107
rect -6756 25087 -6754 25107
rect -6660 25087 -6658 25107
rect -6612 25087 -6610 25107
rect -6516 25087 -6514 25107
rect -5892 25087 -5890 25107
rect -5436 25087 -5434 25107
rect -5340 25087 -5338 25107
rect -5196 25087 -5194 25107
rect -5100 25087 -5098 25107
rect -4716 25087 -4714 25107
rect -4500 25087 -4498 25107
rect -4404 25087 -4402 25107
rect -4308 25087 -4306 25107
rect -4164 25087 -4162 25107
rect -4020 25087 -4018 25107
rect -3876 25087 -3874 25107
rect -3732 25087 -3730 25107
rect -3636 25087 -3634 25107
rect -3540 25087 -3538 25107
rect -3468 25087 -3466 25107
rect -3324 25087 -3322 25107
rect -3108 25087 -3106 25107
rect -3012 25087 -3010 25107
rect -2964 25087 -2962 25107
rect -2916 25087 -2914 25107
rect -2892 25087 -2890 25107
rect -2868 25087 -2866 25107
rect -2820 25087 -2818 25107
rect -2772 25087 -2770 25107
rect -2676 25087 -2674 25107
rect -2364 25087 -2362 25107
rect -2316 25087 -2314 25107
rect -2076 25087 -2074 25107
rect -2052 25087 -2050 25107
rect -1980 25087 -1978 25107
rect -1884 25087 -1882 25107
rect -1572 25087 -1570 25107
rect -1476 25087 -1474 25107
rect -1356 25087 -1354 25107
rect -1260 25087 -1258 25107
rect -1236 25087 -1234 25107
rect -1140 25087 -1138 25107
rect -876 25087 -874 25107
rect -660 25087 -658 25107
rect -492 25087 -490 25107
rect -444 25087 -442 25107
rect -396 25087 -394 25107
rect -348 25087 -346 25107
rect -276 25087 -274 25107
rect -12 25087 -10 25107
rect 156 25087 158 25107
rect 204 25087 206 25107
rect 252 25087 254 25107
rect 348 25087 350 25107
rect 468 25087 470 25107
rect 492 25087 494 25107
rect 564 25087 566 25107
rect 588 25087 590 25107
rect 636 25087 638 25107
rect 660 25087 662 25107
rect 732 25087 734 25107
rect 1092 25087 1094 25107
rect 1140 25087 1142 25107
rect 1308 25087 1310 25107
rect 1345 25102 1348 25107
rect 1355 25088 1358 25102
rect 1356 25087 1358 25088
rect 1428 25087 1430 25107
rect 1476 25104 1478 25107
rect 1476 25087 1479 25104
rect 1692 25087 1694 25107
rect 1860 25087 1862 25107
rect 2028 25087 2030 25107
rect 2076 25087 2078 25107
rect 2100 25087 2102 25107
rect 2124 25087 2126 25107
rect 2244 25087 2246 25107
rect 2412 25087 2414 25107
rect 2460 25087 2462 25107
rect 2508 25087 2510 25107
rect 2604 25087 2606 25107
rect 2772 25087 2774 25107
rect 2868 25087 2870 25107
rect 2940 25087 2942 25107
rect 3012 25087 3014 25107
rect 3108 25087 3110 25107
rect 3324 25087 3326 25107
rect 3396 25087 3398 25107
rect 3564 25087 3566 25107
rect 3636 25087 3638 25107
rect 3660 25087 3662 25107
rect 3732 25087 3734 25107
rect 3780 25087 3782 25107
rect 3828 25087 3830 25107
rect 3924 25087 3926 25107
rect 4020 25087 4022 25107
rect 4092 25087 4094 25107
rect 4188 25087 4190 25107
rect 4308 25087 4310 25107
rect 4404 25087 4406 25107
rect 4500 25087 4502 25107
rect 4596 25087 4598 25107
rect 4692 25087 4694 25107
rect 4860 25104 4862 25107
rect 4860 25087 4863 25104
rect 4956 25087 4958 25107
rect 4980 25087 4982 25107
rect 5052 25087 5054 25107
rect 5124 25087 5126 25107
rect 5220 25087 5222 25107
rect 5268 25087 5270 25107
rect 5388 25087 5390 25107
rect 5484 25087 5486 25107
rect 5508 25087 5510 25107
rect 5532 25087 5534 25107
rect 5628 25087 5630 25107
rect 5652 25087 5654 25107
rect 5748 25087 5750 25107
rect 5796 25087 5798 25107
rect 5844 25087 5846 25107
rect 5892 25087 5894 25107
rect 6132 25087 6134 25107
rect 6228 25087 6230 25107
rect 6252 25087 6254 25107
rect 6276 25087 6278 25107
rect 6324 25087 6326 25107
rect 6372 25087 6374 25107
rect 6420 25087 6422 25107
rect 6492 25087 6494 25107
rect 6516 25087 6518 25107
rect 6588 25087 6590 25107
rect 6612 25087 6614 25107
rect 6660 25087 6662 25107
rect 6684 25087 6686 25107
rect 6708 25087 6710 25107
rect 6780 25087 6782 25107
rect 6804 25087 6806 25107
rect 6900 25087 6902 25107
rect 6924 25087 6926 25107
rect 7020 25087 7022 25107
rect 7164 25087 7166 25107
rect 7236 25087 7238 25107
rect 7308 25087 7310 25107
rect 7380 25087 7382 25107
rect 7393 25102 7396 25107
rect 7403 25088 7406 25102
rect 7404 25087 7406 25088
rect 7452 25087 7454 25107
rect 7476 25087 7478 25107
rect 7524 25104 7526 25107
rect 7524 25087 7527 25104
rect 7548 25087 7550 25107
rect 7572 25087 7574 25107
rect 7620 25087 7622 25107
rect 7644 25087 7646 25107
rect 7668 25087 7670 25107
rect 7908 25087 7910 25107
rect 7956 25087 7958 25107
rect 8124 25087 8126 25107
rect 8220 25087 8222 25107
rect 8652 25087 8654 25107
rect 8700 25087 8702 25107
rect 8748 25087 8750 25107
rect 8796 25087 8798 25107
rect 8844 25087 8846 25107
rect 8868 25087 8870 25107
rect 9516 25087 9518 25107
rect 9660 25087 9662 25107
rect 9684 25087 9686 25107
rect 9756 25087 9758 25107
rect 9780 25087 9782 25107
rect 9804 25087 9806 25107
rect 9852 25087 9854 25107
rect 9900 25087 9902 25107
rect 9948 25087 9950 25107
rect 10044 25087 10046 25107
rect 10116 25087 10118 25107
rect 10188 25087 10190 25107
rect 10284 25087 10286 25107
rect 10332 25087 10334 25107
rect 10380 25087 10382 25107
rect 10428 25087 10430 25107
rect 10476 25087 10478 25107
rect 10500 25087 10502 25107
rect 10524 25087 10526 25107
rect 10596 25087 10598 25107
rect 10620 25087 10622 25107
rect 10644 25087 10646 25107
rect 10716 25087 10718 25107
rect 10956 25087 10958 25107
rect 11004 25087 11006 25107
rect 11052 25087 11054 25107
rect 11100 25087 11102 25107
rect 11172 25087 11174 25107
rect 11220 25087 11222 25107
rect 11340 25087 11342 25107
rect 11436 25087 11438 25107
rect 11532 25087 11534 25107
rect 11628 25087 11630 25107
rect 11676 25087 11678 25107
rect 11724 25087 11726 25107
rect 11772 25087 11774 25107
rect 11796 25087 11798 25107
rect 11892 25087 11894 25107
rect 11988 25087 11990 25107
rect 12060 25087 12062 25107
rect 12228 25087 12230 25107
rect 12276 25087 12278 25107
rect 12324 25087 12326 25107
rect 12420 25087 12422 25107
rect 12444 25087 12446 25107
rect 12516 25087 12518 25107
rect 12540 25087 12542 25107
rect 12553 25087 12611 25088
rect 12636 25087 12638 25107
rect 12732 25087 12734 25107
rect 12756 25087 12758 25107
rect 12804 25087 12806 25107
rect 12828 25087 12830 25107
rect 12972 25087 12974 25107
rect 13044 25087 13046 25107
rect 13068 25087 13070 25107
rect 13116 25087 13118 25107
rect 13284 25087 13286 25107
rect 13332 25087 13334 25107
rect 13572 25087 13574 25107
rect 13620 25087 13622 25107
rect 13668 25087 13670 25107
rect 13716 25087 13718 25107
rect 13764 25087 13766 25107
rect 13860 25087 13862 25107
rect 13956 25087 13958 25107
rect 14004 25087 14006 25107
rect 14100 25087 14102 25107
rect 14940 25087 14942 25107
rect 15036 25087 15038 25107
rect 15180 25087 15182 25107
rect 15276 25087 15278 25107
rect 15420 25087 15422 25107
rect 15492 25087 15494 25107
rect 15660 25087 15662 25107
rect 15708 25087 15710 25107
rect 15732 25087 15734 25107
rect 15756 25087 15758 25107
rect 15804 25087 15806 25107
rect 15828 25087 15830 25107
rect 15852 25087 15854 25107
rect 15948 25087 15950 25107
rect 15972 25087 15974 25107
rect 16044 25087 16046 25107
rect 16068 25087 16070 25107
rect 16164 25087 16166 25107
rect 16260 25087 16262 25107
rect 16332 25087 16334 25107
rect 16548 25087 16550 25107
rect 16572 25087 16574 25107
rect 16620 25087 16622 25107
rect 16668 25087 16670 25107
rect 16716 25087 16718 25107
rect 16764 25087 16766 25107
rect 16812 25087 16814 25107
rect 16884 25087 16886 25107
rect 16908 25087 16910 25107
rect 16980 25087 16982 25107
rect 17148 25087 17150 25107
rect 17196 25087 17198 25107
rect 17220 25087 17222 25107
rect 17292 25087 17294 25107
rect 17316 25087 17318 25107
rect 18132 25087 18134 25107
rect 18228 25087 18230 25107
rect 18492 25087 18494 25107
rect 18516 25087 18518 25107
rect 18564 25088 18566 25107
rect 18529 25087 18587 25088
rect 18612 25087 18614 25107
rect 18660 25087 18662 25107
rect 18745 25102 18748 25107
rect 18756 25102 18758 25107
rect 18755 25088 18758 25102
rect 18828 25087 18831 25104
rect 18900 25087 18902 25107
rect 18924 25087 18926 25107
rect 18996 25087 18998 25107
rect 19020 25087 19022 25107
rect 19092 25087 19094 25107
rect 19140 25087 19142 25107
rect 19236 25087 19238 25107
rect 19260 25087 19262 25107
rect 19788 25087 19790 25107
rect 19836 25087 19838 25107
rect 19860 25087 19862 25107
rect 19884 25087 19886 25107
rect 19956 25087 19958 25107
rect 19980 25087 19982 25107
rect 20052 25087 20054 25107
rect 20076 25087 20078 25107
rect 20124 25087 20126 25107
rect 20172 25087 20174 25107
rect 20196 25087 20198 25107
rect 20292 25087 20294 25107
rect 20343 25104 20357 25107
rect 20388 25087 20390 25107
rect 20412 25087 20414 25107
rect 20508 25087 20510 25107
rect 20532 25087 20534 25107
rect 20604 25087 20606 25107
rect 20607 25104 20621 25107
rect 20628 25107 24515 25111
rect 20628 25104 20645 25107
rect 20628 25087 20630 25104
rect 20964 25087 20966 25107
rect 21012 25087 21014 25107
rect 21108 25087 21110 25107
rect 21204 25087 21206 25107
rect 21300 25087 21302 25107
rect 21324 25087 21326 25107
rect 21444 25087 21446 25107
rect 21468 25087 21470 25107
rect 21564 25087 21566 25107
rect 21588 25087 21590 25107
rect 21684 25087 21686 25107
rect 21708 25087 21710 25107
rect 21828 25087 21830 25107
rect 21924 25087 21926 25107
rect 22068 25087 22070 25107
rect 22188 25087 22190 25107
rect 22212 25087 22214 25107
rect 22884 25087 22886 25107
rect 22980 25087 22982 25107
rect 23076 25087 23078 25107
rect 23100 25087 23102 25107
rect 23124 25087 23126 25107
rect 23244 25087 23246 25107
rect 23340 25087 23342 25107
rect 23412 25087 23414 25107
rect 23460 25087 23462 25107
rect 23508 25087 23510 25107
rect 23556 25087 23558 25107
rect 23604 25087 23606 25107
rect 23652 25087 23654 25107
rect 23676 25087 23678 25107
rect 23700 25087 23702 25107
rect 23772 25087 23774 25107
rect 23796 25087 23798 25107
rect 23916 25087 23918 25107
rect 24012 25087 24014 25107
rect 24060 25087 24062 25107
rect 24156 25087 24158 25107
rect 24481 25102 24484 25107
rect 24492 25104 24494 25107
rect 24492 25102 24495 25104
rect 24491 25088 24495 25102
rect 24409 25087 24443 25088
rect -13319 25083 -8035 25087
rect -13199 25063 -13165 25064
rect -12852 25063 -12850 25083
rect -12636 25063 -12634 25083
rect -12300 25063 -12298 25083
rect -11772 25063 -11770 25083
rect -11676 25063 -11674 25083
rect -11652 25063 -11650 25083
rect -11508 25063 -11506 25083
rect -11436 25063 -11434 25083
rect -11412 25063 -11410 25083
rect -11351 25078 -11348 25083
rect -11340 25078 -11338 25083
rect -11341 25064 -11338 25078
rect -11196 25063 -11194 25083
rect -11100 25063 -11098 25083
rect -10764 25063 -10762 25083
rect -10644 25063 -10642 25083
rect -9900 25063 -9898 25083
rect -9732 25063 -9730 25083
rect -9444 25063 -9442 25083
rect -9348 25063 -9346 25083
rect -9228 25063 -9226 25083
rect -9108 25063 -9106 25083
rect -8436 25063 -8434 25083
rect -8364 25063 -8362 25083
rect -8340 25063 -8338 25083
rect -8268 25063 -8266 25083
rect -8124 25063 -8122 25083
rect -8049 25080 -8035 25083
rect -8028 25083 -7675 25087
rect -8028 25080 -8011 25083
rect -8004 25080 -8001 25083
rect -8028 25063 -8026 25080
rect -7932 25063 -7930 25083
rect -7764 25063 -7762 25083
rect -7689 25080 -7675 25083
rect -7665 25083 1445 25087
rect -7665 25080 -7651 25083
rect -7524 25063 -7522 25083
rect -7356 25063 -7354 25083
rect -7308 25063 -7306 25083
rect -7212 25063 -7210 25083
rect -7044 25063 -7042 25083
rect -6948 25063 -6946 25083
rect -6852 25063 -6850 25083
rect -6756 25063 -6754 25083
rect -6660 25063 -6658 25083
rect -6612 25063 -6610 25083
rect -6516 25063 -6514 25083
rect -5892 25063 -5890 25083
rect -5436 25063 -5434 25083
rect -5340 25063 -5338 25083
rect -5196 25063 -5194 25083
rect -5100 25063 -5098 25083
rect -4716 25063 -4714 25083
rect -4500 25063 -4498 25083
rect -4404 25063 -4402 25083
rect -4308 25063 -4306 25083
rect -4164 25063 -4162 25083
rect -4020 25063 -4018 25083
rect -3876 25063 -3874 25083
rect -3732 25063 -3730 25083
rect -3636 25063 -3634 25083
rect -3540 25063 -3538 25083
rect -3468 25063 -3466 25083
rect -3324 25063 -3322 25083
rect -3108 25063 -3106 25083
rect -3012 25063 -3010 25083
rect -2964 25063 -2962 25083
rect -2916 25063 -2914 25083
rect -2892 25063 -2890 25083
rect -2868 25063 -2866 25083
rect -2820 25063 -2818 25083
rect -2772 25063 -2770 25083
rect -2676 25063 -2674 25083
rect -2364 25063 -2362 25083
rect -2316 25063 -2314 25083
rect -2076 25063 -2074 25083
rect -2052 25063 -2050 25083
rect -1980 25063 -1978 25083
rect -1884 25063 -1882 25083
rect -1572 25063 -1570 25083
rect -1476 25063 -1474 25083
rect -1356 25063 -1354 25083
rect -1260 25063 -1258 25083
rect -1236 25063 -1234 25083
rect -1140 25063 -1138 25083
rect -876 25063 -874 25083
rect -660 25063 -658 25083
rect -492 25063 -490 25083
rect -444 25063 -442 25083
rect -396 25063 -394 25083
rect -348 25063 -346 25083
rect -276 25063 -274 25083
rect -12 25063 -10 25083
rect 156 25063 158 25083
rect 204 25063 206 25083
rect 252 25063 254 25083
rect 348 25063 350 25083
rect 468 25063 470 25083
rect 492 25063 494 25083
rect 564 25063 566 25083
rect 588 25063 590 25083
rect 636 25063 638 25083
rect 660 25063 662 25083
rect 732 25063 734 25083
rect 793 25063 827 25064
rect 1092 25063 1094 25083
rect 1140 25063 1142 25083
rect 1308 25063 1310 25083
rect 1356 25063 1358 25083
rect 1428 25063 1430 25083
rect 1431 25080 1445 25083
rect 1455 25083 7493 25087
rect 1455 25080 1469 25083
rect 1476 25080 1479 25083
rect 1692 25063 1694 25083
rect 1860 25063 1862 25083
rect 2028 25063 2030 25083
rect 2076 25063 2078 25083
rect 2100 25063 2102 25083
rect 2124 25063 2126 25083
rect 2244 25063 2246 25083
rect 2412 25063 2414 25083
rect 2460 25063 2462 25083
rect 2508 25063 2510 25083
rect 2604 25063 2606 25083
rect 2772 25063 2774 25083
rect 2868 25063 2870 25083
rect 2940 25063 2942 25083
rect 3012 25063 3014 25083
rect 3108 25063 3110 25083
rect 3324 25063 3326 25083
rect 3396 25063 3398 25083
rect 3564 25063 3566 25083
rect 3636 25063 3638 25083
rect 3660 25063 3662 25083
rect 3732 25063 3734 25083
rect 3780 25063 3782 25083
rect 3828 25063 3830 25083
rect 3924 25063 3926 25083
rect 4020 25063 4022 25083
rect 4092 25063 4094 25083
rect 4188 25063 4190 25083
rect 4308 25063 4310 25083
rect 4404 25063 4406 25083
rect 4500 25063 4502 25083
rect 4596 25063 4598 25083
rect 4692 25063 4694 25083
rect 4839 25080 4853 25083
rect 4860 25080 4863 25083
rect 4956 25063 4958 25083
rect 4980 25063 4982 25083
rect 5052 25063 5054 25083
rect 5124 25063 5126 25083
rect 5220 25063 5222 25083
rect 5268 25063 5270 25083
rect 5388 25063 5390 25083
rect 5484 25063 5486 25083
rect 5508 25063 5510 25083
rect 5532 25063 5534 25083
rect 5628 25063 5630 25083
rect 5652 25063 5654 25083
rect 5748 25063 5750 25083
rect 5796 25063 5798 25083
rect 5844 25063 5846 25083
rect 5892 25063 5894 25083
rect 6132 25063 6134 25083
rect 6228 25063 6230 25083
rect 6252 25063 6254 25083
rect 6276 25063 6278 25083
rect 6324 25063 6326 25083
rect 6372 25063 6374 25083
rect 6420 25063 6422 25083
rect 6492 25063 6494 25083
rect 6516 25063 6518 25083
rect 6588 25063 6590 25083
rect 6612 25063 6614 25083
rect 6660 25063 6662 25083
rect 6684 25063 6686 25083
rect 6708 25063 6710 25083
rect 6780 25063 6782 25083
rect 6804 25063 6806 25083
rect 6900 25063 6902 25083
rect 6924 25063 6926 25083
rect 7020 25063 7022 25083
rect 7164 25063 7166 25083
rect 7236 25063 7238 25083
rect 7308 25063 7310 25083
rect 7380 25063 7382 25083
rect 7404 25063 7406 25083
rect 7452 25064 7454 25083
rect 7441 25063 7475 25064
rect 7476 25063 7478 25083
rect 7479 25080 7493 25083
rect 7503 25083 18821 25087
rect 7503 25080 7517 25083
rect 7524 25080 7527 25083
rect 7548 25063 7550 25083
rect 7572 25063 7574 25083
rect 7620 25063 7622 25083
rect 7644 25063 7646 25083
rect 7668 25063 7670 25083
rect 7908 25063 7910 25083
rect 7956 25063 7958 25083
rect 8124 25063 8126 25083
rect 8220 25063 8222 25083
rect 8652 25063 8654 25083
rect 8700 25063 8702 25083
rect 8748 25063 8750 25083
rect 8796 25063 8798 25083
rect 8844 25063 8846 25083
rect 8868 25063 8870 25083
rect 9516 25063 9518 25083
rect 9660 25063 9662 25083
rect 9684 25063 9686 25083
rect 9756 25063 9758 25083
rect 9780 25063 9782 25083
rect 9804 25063 9806 25083
rect 9852 25063 9854 25083
rect 9900 25063 9902 25083
rect 9948 25063 9950 25083
rect 10044 25063 10046 25083
rect 10116 25063 10118 25083
rect 10188 25063 10190 25083
rect 10284 25063 10286 25083
rect 10332 25063 10334 25083
rect 10380 25063 10382 25083
rect 10428 25063 10430 25083
rect 10476 25063 10478 25083
rect 10500 25064 10502 25083
rect 10489 25063 10523 25064
rect 10524 25063 10526 25083
rect 10596 25064 10598 25083
rect 10585 25063 10619 25064
rect 10620 25063 10622 25083
rect 10644 25063 10646 25083
rect 10716 25063 10718 25083
rect 10956 25063 10958 25083
rect 11004 25063 11006 25083
rect 11052 25063 11054 25083
rect 11100 25063 11102 25083
rect 11172 25063 11174 25083
rect 11220 25063 11222 25083
rect 11340 25063 11342 25083
rect 11436 25063 11438 25083
rect 11532 25063 11534 25083
rect 11628 25063 11630 25083
rect 11676 25063 11678 25083
rect 11724 25063 11726 25083
rect 11772 25063 11774 25083
rect 11796 25063 11798 25083
rect 11892 25063 11894 25083
rect 11988 25063 11990 25083
rect 12060 25063 12062 25083
rect 12121 25063 12155 25064
rect 12228 25063 12230 25083
rect 12276 25063 12278 25083
rect 12324 25063 12326 25083
rect 12420 25063 12422 25083
rect 12444 25063 12446 25083
rect 12516 25063 12518 25083
rect 12540 25063 12542 25083
rect 12553 25078 12556 25083
rect 12563 25064 12566 25078
rect 12636 25064 12638 25083
rect 12564 25063 12566 25064
rect 12625 25063 12653 25064
rect -13199 25059 -9691 25063
rect -13079 25039 -13045 25040
rect -12852 25039 -12850 25059
rect -12636 25039 -12634 25059
rect -12431 25039 -12373 25040
rect -12300 25039 -12298 25059
rect -11772 25039 -11770 25059
rect -11676 25039 -11674 25059
rect -11652 25039 -11650 25059
rect -11508 25039 -11506 25059
rect -11436 25039 -11434 25059
rect -11412 25039 -11410 25059
rect -11265 25056 -11251 25059
rect -11196 25039 -11194 25059
rect -11100 25039 -11098 25059
rect -10895 25039 -10861 25040
rect -10764 25039 -10762 25059
rect -10644 25039 -10642 25059
rect -9900 25039 -9898 25059
rect -9732 25039 -9730 25059
rect -9705 25056 -9691 25059
rect -9681 25059 12653 25063
rect -9681 25056 -9667 25059
rect -9444 25039 -9442 25059
rect -9348 25039 -9346 25059
rect -9228 25039 -9226 25059
rect -9108 25039 -9106 25059
rect -8436 25039 -8434 25059
rect -8364 25039 -8362 25059
rect -8340 25039 -8338 25059
rect -8268 25039 -8266 25059
rect -8124 25039 -8122 25059
rect -8028 25039 -8026 25059
rect -7932 25039 -7930 25059
rect -7764 25039 -7762 25059
rect -7524 25039 -7522 25059
rect -7356 25039 -7354 25059
rect -7308 25039 -7306 25059
rect -7212 25039 -7210 25059
rect -7044 25039 -7042 25059
rect -6948 25039 -6946 25059
rect -6852 25039 -6850 25059
rect -6756 25039 -6754 25059
rect -6660 25039 -6658 25059
rect -6612 25039 -6610 25059
rect -6516 25039 -6514 25059
rect -5892 25039 -5890 25059
rect -5436 25039 -5434 25059
rect -5340 25039 -5338 25059
rect -5196 25039 -5194 25059
rect -5100 25039 -5098 25059
rect -4716 25039 -4714 25059
rect -4500 25039 -4498 25059
rect -4404 25039 -4402 25059
rect -4308 25039 -4306 25059
rect -4164 25039 -4162 25059
rect -4020 25039 -4018 25059
rect -3876 25039 -3874 25059
rect -3732 25039 -3730 25059
rect -3636 25039 -3634 25059
rect -3540 25039 -3538 25059
rect -3468 25039 -3466 25059
rect -3324 25039 -3322 25059
rect -3108 25039 -3106 25059
rect -3012 25039 -3010 25059
rect -2964 25039 -2962 25059
rect -2916 25039 -2914 25059
rect -2892 25039 -2890 25059
rect -2868 25039 -2866 25059
rect -2820 25039 -2818 25059
rect -2772 25039 -2770 25059
rect -2676 25039 -2674 25059
rect -2364 25039 -2362 25059
rect -2316 25039 -2314 25059
rect -2076 25039 -2074 25059
rect -2052 25039 -2050 25059
rect -1980 25039 -1978 25059
rect -1884 25039 -1882 25059
rect -1572 25039 -1570 25059
rect -1476 25039 -1474 25059
rect -1356 25039 -1354 25059
rect -1260 25039 -1258 25059
rect -1236 25039 -1234 25059
rect -1140 25039 -1138 25059
rect -876 25039 -874 25059
rect -660 25039 -658 25059
rect -492 25039 -490 25059
rect -444 25039 -442 25059
rect -396 25039 -394 25059
rect -348 25039 -346 25059
rect -276 25039 -274 25059
rect -12 25039 -10 25059
rect 156 25039 158 25059
rect 204 25039 206 25059
rect 252 25039 254 25059
rect 348 25039 350 25059
rect 468 25039 470 25059
rect 492 25039 494 25059
rect 564 25039 566 25059
rect 588 25039 590 25059
rect 636 25039 638 25059
rect 660 25039 662 25059
rect 732 25039 734 25059
rect 1092 25039 1094 25059
rect 1140 25039 1142 25059
rect 1308 25039 1310 25059
rect 1356 25039 1358 25059
rect 1428 25039 1430 25059
rect 1692 25039 1694 25059
rect 1860 25039 1862 25059
rect 2028 25039 2030 25059
rect 2076 25039 2078 25059
rect 2100 25039 2102 25059
rect 2124 25039 2126 25059
rect 2244 25039 2246 25059
rect 2412 25039 2414 25059
rect 2460 25039 2462 25059
rect 2508 25039 2510 25059
rect 2604 25039 2606 25059
rect 2772 25039 2774 25059
rect 2868 25039 2870 25059
rect 2940 25039 2942 25059
rect 3012 25039 3014 25059
rect 3108 25039 3110 25059
rect 3324 25039 3326 25059
rect 3396 25039 3398 25059
rect 3564 25039 3566 25059
rect 3636 25039 3638 25059
rect 3660 25039 3662 25059
rect 3732 25039 3734 25059
rect 3780 25039 3782 25059
rect 3828 25039 3830 25059
rect 3924 25039 3926 25059
rect 4020 25039 4022 25059
rect 4092 25039 4094 25059
rect 4188 25039 4190 25059
rect 4308 25039 4310 25059
rect 4404 25039 4406 25059
rect 4500 25039 4502 25059
rect 4596 25039 4598 25059
rect 4692 25039 4694 25059
rect 4956 25039 4958 25059
rect 4980 25039 4982 25059
rect 5052 25039 5054 25059
rect 5124 25039 5126 25059
rect 5220 25039 5222 25059
rect 5268 25039 5270 25059
rect 5388 25039 5390 25059
rect 5484 25039 5486 25059
rect 5508 25039 5510 25059
rect 5532 25039 5534 25059
rect 5628 25039 5630 25059
rect 5652 25039 5654 25059
rect 5748 25039 5750 25059
rect 5796 25039 5798 25059
rect 5844 25039 5846 25059
rect 5892 25039 5894 25059
rect 6132 25039 6134 25059
rect 6228 25039 6230 25059
rect 6252 25039 6254 25059
rect 6276 25039 6278 25059
rect 6324 25039 6326 25059
rect 6372 25039 6374 25059
rect 6420 25039 6422 25059
rect 6492 25039 6494 25059
rect 6516 25039 6518 25059
rect 6588 25039 6590 25059
rect 6612 25039 6614 25059
rect 6660 25039 6662 25059
rect 6684 25039 6686 25059
rect 6708 25039 6710 25059
rect 6780 25039 6782 25059
rect 6804 25039 6806 25059
rect 6900 25039 6902 25059
rect 6924 25039 6926 25059
rect 7020 25039 7022 25059
rect 7164 25039 7166 25059
rect 7236 25039 7238 25059
rect 7308 25039 7310 25059
rect 7380 25039 7382 25059
rect 7404 25039 7406 25059
rect 7441 25054 7444 25059
rect 7452 25054 7454 25059
rect 7451 25040 7454 25054
rect 7476 25039 7478 25059
rect 7548 25056 7550 25059
rect 7548 25039 7551 25056
rect 7572 25039 7574 25059
rect 7620 25039 7622 25059
rect 7644 25039 7646 25059
rect 7668 25039 7670 25059
rect 7908 25039 7910 25059
rect 7956 25039 7958 25059
rect 8124 25039 8126 25059
rect 8220 25039 8222 25059
rect 8652 25039 8654 25059
rect 8700 25039 8702 25059
rect 8748 25039 8750 25059
rect 8796 25039 8798 25059
rect 8844 25039 8846 25059
rect 8868 25039 8870 25059
rect 9516 25039 9518 25059
rect 9660 25039 9662 25059
rect 9684 25039 9686 25059
rect 9756 25039 9758 25059
rect 9780 25039 9782 25059
rect 9804 25039 9806 25059
rect 9852 25039 9854 25059
rect 9900 25039 9902 25059
rect 9948 25039 9950 25059
rect 10044 25039 10046 25059
rect 10116 25039 10118 25059
rect 10188 25039 10190 25059
rect 10284 25039 10286 25059
rect 10332 25039 10334 25059
rect 10380 25039 10382 25059
rect 10428 25039 10430 25059
rect 10476 25039 10478 25059
rect 10489 25054 10492 25059
rect 10500 25054 10502 25059
rect 10499 25040 10502 25054
rect 10524 25039 10526 25059
rect 10585 25054 10588 25059
rect 10596 25056 10598 25059
rect 10596 25054 10599 25056
rect 10595 25040 10599 25054
rect 10620 25039 10622 25059
rect 10644 25039 10646 25059
rect 10716 25039 10718 25059
rect 10956 25039 10958 25059
rect 11004 25039 11006 25059
rect 11052 25039 11054 25059
rect 11100 25039 11102 25059
rect 11172 25039 11174 25059
rect 11220 25039 11222 25059
rect 11340 25039 11342 25059
rect 11436 25039 11438 25059
rect 11532 25039 11534 25059
rect 11628 25039 11630 25059
rect 11676 25039 11678 25059
rect 11724 25039 11726 25059
rect 11772 25039 11774 25059
rect 11796 25039 11798 25059
rect 11892 25039 11894 25059
rect 11988 25039 11990 25059
rect 12060 25039 12062 25059
rect 12228 25056 12230 25059
rect 12228 25039 12231 25056
rect 12276 25039 12278 25059
rect 12324 25039 12326 25059
rect 12420 25039 12422 25059
rect 12444 25039 12446 25059
rect 12516 25039 12518 25059
rect 12540 25039 12542 25059
rect 12564 25039 12566 25059
rect 12625 25054 12628 25059
rect 12636 25054 12638 25059
rect 12639 25056 12653 25059
rect 12660 25063 12663 25080
rect 12732 25063 12734 25083
rect 12756 25063 12758 25083
rect 12804 25063 12806 25083
rect 12828 25063 12830 25083
rect 12972 25063 12974 25083
rect 13044 25063 13046 25083
rect 13068 25063 13070 25083
rect 13116 25063 13118 25083
rect 13284 25063 13286 25083
rect 13332 25063 13334 25083
rect 13489 25063 13547 25064
rect 13572 25063 13574 25083
rect 13620 25063 13622 25083
rect 13668 25063 13670 25083
rect 13716 25063 13718 25083
rect 13764 25063 13766 25083
rect 13860 25063 13862 25083
rect 13956 25063 13958 25083
rect 14004 25063 14006 25083
rect 14100 25063 14102 25083
rect 14940 25063 14942 25083
rect 15036 25063 15038 25083
rect 15180 25063 15182 25083
rect 15276 25063 15278 25083
rect 15420 25063 15422 25083
rect 15492 25063 15494 25083
rect 15660 25063 15662 25083
rect 15708 25063 15710 25083
rect 15732 25063 15734 25083
rect 15756 25063 15758 25083
rect 15804 25063 15806 25083
rect 15828 25063 15830 25083
rect 15852 25063 15854 25083
rect 15948 25063 15950 25083
rect 15972 25063 15974 25083
rect 16044 25063 16046 25083
rect 16068 25063 16070 25083
rect 16164 25063 16166 25083
rect 16260 25063 16262 25083
rect 16332 25063 16334 25083
rect 16548 25063 16550 25083
rect 16572 25063 16574 25083
rect 16620 25063 16622 25083
rect 16668 25063 16670 25083
rect 16716 25063 16718 25083
rect 16764 25063 16766 25083
rect 16812 25063 16814 25083
rect 16884 25063 16886 25083
rect 16908 25063 16910 25083
rect 16980 25063 16982 25083
rect 17148 25063 17150 25083
rect 17196 25063 17198 25083
rect 17220 25063 17222 25083
rect 17292 25063 17294 25083
rect 17316 25063 17318 25083
rect 18132 25063 18134 25083
rect 18228 25063 18230 25083
rect 18492 25063 18494 25083
rect 18516 25063 18518 25083
rect 18553 25078 18556 25083
rect 18564 25078 18566 25083
rect 18563 25064 18566 25078
rect 18612 25063 18614 25083
rect 18660 25080 18662 25083
rect 18807 25080 18821 25083
rect 18828 25083 24443 25087
rect 18828 25080 18845 25083
rect 18660 25063 18663 25080
rect 18828 25063 18830 25080
rect 18900 25063 18902 25083
rect 18924 25063 18926 25083
rect 18996 25063 18998 25083
rect 19020 25063 19022 25083
rect 19092 25063 19094 25083
rect 19140 25063 19142 25083
rect 19236 25063 19238 25083
rect 19260 25063 19262 25083
rect 19788 25063 19790 25083
rect 19836 25063 19838 25083
rect 19860 25063 19862 25083
rect 19884 25063 19886 25083
rect 19956 25063 19958 25083
rect 19980 25063 19982 25083
rect 20052 25063 20054 25083
rect 20076 25063 20078 25083
rect 20124 25063 20126 25083
rect 20172 25063 20174 25083
rect 20196 25063 20198 25083
rect 20292 25063 20294 25083
rect 20388 25063 20390 25083
rect 20412 25063 20414 25083
rect 20508 25063 20510 25083
rect 20532 25063 20534 25083
rect 20604 25063 20606 25083
rect 20628 25063 20630 25083
rect 20964 25063 20966 25083
rect 21012 25063 21014 25083
rect 21108 25063 21110 25083
rect 21204 25063 21206 25083
rect 21300 25063 21302 25083
rect 21324 25063 21326 25083
rect 21444 25063 21446 25083
rect 21468 25063 21470 25083
rect 21564 25063 21566 25083
rect 21588 25063 21590 25083
rect 21684 25063 21686 25083
rect 21708 25063 21710 25083
rect 21828 25063 21830 25083
rect 21924 25063 21926 25083
rect 22068 25063 22070 25083
rect 22188 25063 22190 25083
rect 22212 25063 22214 25083
rect 22884 25063 22886 25083
rect 22980 25063 22982 25083
rect 23076 25063 23078 25083
rect 23100 25063 23102 25083
rect 23124 25063 23126 25083
rect 23244 25063 23246 25083
rect 23340 25063 23342 25083
rect 23412 25063 23414 25083
rect 23460 25063 23462 25083
rect 23508 25063 23510 25083
rect 23556 25063 23558 25083
rect 23604 25063 23606 25083
rect 23652 25063 23654 25083
rect 23676 25063 23678 25083
rect 23700 25063 23702 25083
rect 23772 25063 23774 25083
rect 23796 25063 23798 25083
rect 23916 25063 23918 25083
rect 24012 25063 24014 25083
rect 24060 25063 24062 25083
rect 24156 25063 24158 25083
rect 24265 25063 24299 25064
rect 12660 25059 18629 25063
rect 12660 25056 12677 25059
rect 12732 25056 12734 25059
rect 12635 25040 12638 25054
rect 12660 25039 12662 25056
rect 12732 25039 12735 25056
rect 12756 25039 12758 25059
rect 12804 25040 12806 25059
rect 12769 25039 12827 25040
rect 12828 25039 12830 25059
rect 12972 25039 12974 25059
rect 13044 25039 13046 25059
rect 13068 25039 13070 25059
rect 13116 25039 13118 25059
rect 13284 25039 13286 25059
rect 13332 25039 13334 25059
rect 13489 25054 13492 25059
rect 13499 25040 13502 25054
rect 13500 25039 13502 25040
rect 13572 25039 13574 25059
rect 13620 25056 13622 25059
rect 13620 25039 13623 25056
rect 13668 25039 13670 25059
rect 13716 25039 13718 25059
rect 13764 25039 13766 25059
rect 13860 25039 13862 25059
rect 13956 25039 13958 25059
rect 14004 25039 14006 25059
rect 14100 25039 14102 25059
rect 14940 25039 14942 25059
rect 15036 25039 15038 25059
rect 15180 25039 15182 25059
rect 15276 25039 15278 25059
rect 15420 25039 15422 25059
rect 15492 25039 15494 25059
rect 15660 25039 15662 25059
rect 15708 25039 15710 25059
rect 15732 25039 15734 25059
rect 15756 25039 15758 25059
rect 15804 25039 15806 25059
rect 15828 25039 15830 25059
rect 15852 25039 15854 25059
rect 15948 25039 15950 25059
rect 15972 25039 15974 25059
rect 16044 25039 16046 25059
rect 16068 25039 16070 25059
rect 16164 25039 16166 25059
rect 16260 25039 16262 25059
rect 16332 25039 16334 25059
rect 16548 25039 16550 25059
rect 16572 25039 16574 25059
rect 16620 25039 16622 25059
rect 16668 25039 16670 25059
rect 16716 25039 16718 25059
rect 16764 25039 16766 25059
rect 16812 25039 16814 25059
rect 16884 25039 16886 25059
rect 16908 25039 16910 25059
rect 16980 25039 16982 25059
rect 17148 25039 17150 25059
rect 17196 25039 17198 25059
rect 17220 25039 17222 25059
rect 17292 25039 17294 25059
rect 17316 25039 17318 25059
rect 18132 25039 18134 25059
rect 18228 25039 18230 25059
rect 18492 25039 18494 25059
rect 18516 25039 18518 25059
rect 18612 25039 18614 25059
rect 18615 25056 18629 25059
rect 18639 25059 24299 25063
rect 18639 25056 18653 25059
rect 18660 25056 18663 25059
rect 18828 25039 18830 25059
rect 18900 25039 18902 25059
rect 18924 25039 18926 25059
rect 18996 25039 18998 25059
rect 19020 25039 19022 25059
rect 19092 25039 19094 25059
rect 19140 25039 19142 25059
rect 19236 25039 19238 25059
rect 19260 25039 19262 25059
rect 19788 25039 19790 25059
rect 19836 25039 19838 25059
rect 19860 25039 19862 25059
rect 19884 25039 19886 25059
rect 19956 25039 19958 25059
rect 19980 25039 19982 25059
rect 20052 25039 20054 25059
rect 20076 25039 20078 25059
rect 20124 25039 20126 25059
rect 20172 25039 20174 25059
rect 20196 25039 20198 25059
rect 20292 25039 20294 25059
rect 20388 25039 20390 25059
rect 20412 25039 20414 25059
rect 20508 25039 20510 25059
rect 20532 25039 20534 25059
rect 20604 25039 20606 25059
rect 20628 25039 20630 25059
rect 20881 25039 20939 25040
rect 20964 25039 20966 25059
rect 21012 25039 21014 25059
rect 21108 25039 21110 25059
rect 21204 25039 21206 25059
rect 21300 25039 21302 25059
rect 21324 25039 21326 25059
rect 21444 25039 21446 25059
rect 21468 25039 21470 25059
rect 21564 25039 21566 25059
rect 21588 25039 21590 25059
rect 21684 25039 21686 25059
rect 21708 25039 21710 25059
rect 21828 25039 21830 25059
rect 21924 25039 21926 25059
rect 22068 25039 22070 25059
rect 22188 25039 22190 25059
rect 22212 25039 22214 25059
rect 22884 25039 22886 25059
rect 22980 25039 22982 25059
rect 23076 25039 23078 25059
rect 23100 25039 23102 25059
rect 23124 25039 23126 25059
rect 23244 25039 23246 25059
rect 23340 25039 23342 25059
rect 23412 25039 23414 25059
rect 23460 25039 23462 25059
rect 23508 25039 23510 25059
rect 23556 25039 23558 25059
rect 23604 25039 23606 25059
rect 23652 25039 23654 25059
rect 23676 25039 23678 25059
rect 23700 25039 23702 25059
rect 23772 25039 23774 25059
rect 23796 25039 23798 25059
rect 23916 25039 23918 25059
rect 24012 25039 24014 25059
rect 24060 25040 24062 25059
rect 24156 25040 24158 25059
rect 24025 25039 24083 25040
rect 24145 25039 24179 25040
rect -13079 25035 13589 25039
rect -12959 25015 -12925 25016
rect -12852 25015 -12850 25035
rect -12636 25015 -12634 25035
rect -12431 25030 -12428 25035
rect -12300 25032 -12298 25035
rect -12421 25016 -12418 25030
rect -12420 25015 -12418 25016
rect -12300 25015 -12297 25032
rect -12095 25015 -12037 25016
rect -11772 25015 -11770 25035
rect -11676 25015 -11674 25035
rect -11652 25015 -11650 25035
rect -11508 25015 -11506 25035
rect -11436 25015 -11434 25035
rect -11412 25015 -11410 25035
rect -11196 25015 -11194 25035
rect -11100 25015 -11098 25035
rect -10764 25015 -10762 25035
rect -10644 25015 -10642 25035
rect -9900 25015 -9898 25035
rect -9732 25015 -9730 25035
rect -9444 25015 -9442 25035
rect -9348 25015 -9346 25035
rect -9228 25015 -9226 25035
rect -9108 25015 -9106 25035
rect -8436 25015 -8434 25035
rect -8364 25015 -8362 25035
rect -8340 25015 -8338 25035
rect -8268 25015 -8266 25035
rect -8124 25015 -8122 25035
rect -8028 25015 -8026 25035
rect -7932 25015 -7930 25035
rect -7764 25015 -7762 25035
rect -7583 25015 -7549 25016
rect -7524 25015 -7522 25035
rect -7356 25015 -7354 25035
rect -7308 25015 -7306 25035
rect -7212 25015 -7210 25035
rect -7044 25015 -7042 25035
rect -6948 25015 -6946 25035
rect -6852 25015 -6850 25035
rect -6756 25016 -6754 25035
rect -6767 25015 -6685 25016
rect -6660 25015 -6658 25035
rect -6612 25015 -6610 25035
rect -6516 25015 -6514 25035
rect -5892 25015 -5890 25035
rect -5436 25015 -5434 25035
rect -5340 25015 -5338 25035
rect -5196 25015 -5194 25035
rect -5100 25015 -5098 25035
rect -4716 25015 -4714 25035
rect -4500 25015 -4498 25035
rect -4404 25015 -4402 25035
rect -4308 25015 -4306 25035
rect -4164 25015 -4162 25035
rect -4020 25015 -4018 25035
rect -3876 25015 -3874 25035
rect -3732 25015 -3730 25035
rect -3636 25015 -3634 25035
rect -3540 25015 -3538 25035
rect -3468 25015 -3466 25035
rect -3324 25015 -3322 25035
rect -3108 25015 -3106 25035
rect -3012 25015 -3010 25035
rect -2964 25015 -2962 25035
rect -2916 25015 -2914 25035
rect -2892 25015 -2890 25035
rect -2868 25015 -2866 25035
rect -2820 25015 -2818 25035
rect -2772 25015 -2770 25035
rect -2676 25015 -2674 25035
rect -2364 25015 -2362 25035
rect -2316 25015 -2314 25035
rect -2159 25015 -2125 25016
rect -2076 25015 -2074 25035
rect -2052 25015 -2050 25035
rect -1980 25015 -1978 25035
rect -1884 25016 -1882 25035
rect -1919 25015 -1861 25016
rect -1572 25015 -1570 25035
rect -1476 25015 -1474 25035
rect -1356 25015 -1354 25035
rect -1260 25015 -1258 25035
rect -1236 25015 -1234 25035
rect -1140 25015 -1138 25035
rect -876 25015 -874 25035
rect -660 25015 -658 25035
rect -492 25015 -490 25035
rect -444 25015 -442 25035
rect -396 25015 -394 25035
rect -348 25015 -346 25035
rect -276 25015 -274 25035
rect -12 25015 -10 25035
rect 156 25015 158 25035
rect 204 25015 206 25035
rect 252 25015 254 25035
rect 348 25015 350 25035
rect 468 25015 470 25035
rect 492 25015 494 25035
rect 564 25015 566 25035
rect 588 25015 590 25035
rect 636 25015 638 25035
rect 660 25015 662 25035
rect 732 25015 734 25035
rect 879 25032 893 25035
rect 1092 25015 1094 25035
rect 1140 25015 1142 25035
rect 1308 25015 1310 25035
rect 1356 25015 1358 25035
rect 1428 25015 1430 25035
rect 1692 25015 1694 25035
rect 1860 25015 1862 25035
rect 2028 25016 2030 25035
rect 2017 25015 2051 25016
rect 2076 25015 2078 25035
rect 2100 25015 2102 25035
rect 2124 25015 2126 25035
rect 2244 25015 2246 25035
rect 2412 25016 2414 25035
rect 2305 25015 2339 25016
rect 2401 25015 2435 25016
rect 2460 25015 2462 25035
rect 2508 25015 2510 25035
rect 2604 25016 2606 25035
rect 2593 25015 2627 25016
rect 2772 25015 2774 25035
rect 2868 25015 2870 25035
rect 2940 25015 2942 25035
rect 3012 25015 3014 25035
rect 3108 25015 3110 25035
rect 3324 25015 3326 25035
rect 3396 25015 3398 25035
rect 3564 25015 3566 25035
rect 3636 25016 3638 25035
rect 3625 25015 3659 25016
rect 3660 25015 3662 25035
rect 3732 25015 3734 25035
rect 3780 25015 3782 25035
rect 3828 25015 3830 25035
rect 3924 25015 3926 25035
rect 4020 25015 4022 25035
rect 4092 25015 4094 25035
rect 4188 25015 4190 25035
rect 4308 25015 4310 25035
rect 4404 25015 4406 25035
rect 4500 25015 4502 25035
rect 4596 25015 4598 25035
rect 4692 25015 4694 25035
rect 4956 25015 4958 25035
rect 4980 25015 4982 25035
rect 5052 25015 5054 25035
rect 5124 25015 5126 25035
rect 5220 25015 5222 25035
rect 5268 25015 5270 25035
rect 5388 25015 5390 25035
rect 5484 25015 5486 25035
rect 5508 25015 5510 25035
rect 5532 25015 5534 25035
rect 5628 25015 5630 25035
rect 5652 25015 5654 25035
rect 5748 25015 5750 25035
rect 5796 25015 5798 25035
rect 5844 25015 5846 25035
rect 5892 25015 5894 25035
rect 6132 25015 6134 25035
rect 6228 25015 6230 25035
rect 6252 25015 6254 25035
rect 6276 25015 6278 25035
rect 6324 25015 6326 25035
rect 6372 25015 6374 25035
rect 6420 25015 6422 25035
rect 6492 25015 6494 25035
rect 6516 25015 6518 25035
rect 6588 25015 6590 25035
rect 6612 25015 6614 25035
rect 6660 25016 6662 25035
rect 6625 25015 6683 25016
rect 6684 25015 6686 25035
rect 6708 25015 6710 25035
rect 6780 25015 6782 25035
rect 6804 25015 6806 25035
rect 6900 25015 6902 25035
rect 6924 25015 6926 25035
rect 7020 25015 7022 25035
rect 7164 25015 7166 25035
rect 7236 25015 7238 25035
rect 7308 25015 7310 25035
rect 7380 25015 7382 25035
rect 7404 25015 7406 25035
rect 7476 25015 7478 25035
rect 7527 25032 7541 25035
rect 7548 25032 7551 25035
rect 7572 25015 7574 25035
rect 7620 25015 7622 25035
rect 7644 25015 7646 25035
rect 7668 25015 7670 25035
rect 7908 25015 7910 25035
rect 7956 25015 7958 25035
rect 8124 25015 8126 25035
rect 8220 25015 8222 25035
rect 8652 25015 8654 25035
rect 8700 25015 8702 25035
rect 8748 25015 8750 25035
rect 8796 25015 8798 25035
rect 8844 25015 8846 25035
rect 8868 25015 8870 25035
rect 9516 25015 9518 25035
rect 9660 25015 9662 25035
rect 9684 25015 9686 25035
rect 9756 25015 9758 25035
rect 9780 25015 9782 25035
rect 9804 25015 9806 25035
rect 9852 25015 9854 25035
rect 9900 25015 9902 25035
rect 9948 25015 9950 25035
rect 10044 25015 10046 25035
rect 10116 25015 10118 25035
rect 10188 25015 10190 25035
rect 10284 25015 10286 25035
rect 10332 25015 10334 25035
rect 10380 25015 10382 25035
rect 10428 25015 10430 25035
rect 10476 25015 10478 25035
rect 10524 25015 10526 25035
rect 10575 25032 10589 25035
rect 10620 25015 10622 25035
rect 10644 25015 10646 25035
rect 10671 25032 10685 25035
rect 10716 25015 10718 25035
rect 10956 25015 10958 25035
rect 11004 25015 11006 25035
rect 11052 25015 11054 25035
rect 11100 25015 11102 25035
rect 11172 25015 11174 25035
rect 11220 25015 11222 25035
rect 11340 25015 11342 25035
rect 11436 25015 11438 25035
rect 11532 25015 11534 25035
rect 11628 25015 11630 25035
rect 11676 25015 11678 25035
rect 11724 25015 11726 25035
rect 11772 25015 11774 25035
rect 11796 25015 11798 25035
rect 11892 25015 11894 25035
rect 11988 25015 11990 25035
rect 12060 25015 12062 25035
rect 12207 25032 12221 25035
rect 12228 25032 12231 25035
rect 12276 25015 12278 25035
rect 12324 25015 12326 25035
rect 12420 25015 12422 25035
rect 12444 25015 12446 25035
rect 12516 25015 12518 25035
rect 12540 25015 12542 25035
rect 12564 25015 12566 25035
rect 12660 25015 12662 25035
rect 12711 25032 12725 25035
rect 12732 25032 12735 25035
rect 12756 25015 12758 25035
rect 12793 25030 12796 25035
rect 12804 25030 12806 25035
rect 12803 25016 12806 25030
rect 12828 25015 12830 25035
rect 12876 25015 12879 25032
rect 12972 25015 12974 25035
rect 13044 25015 13046 25035
rect 13068 25015 13070 25035
rect 13116 25015 13118 25035
rect 13284 25015 13286 25035
rect 13332 25015 13334 25035
rect 13500 25015 13502 25035
rect 13572 25015 13574 25035
rect 13575 25032 13589 25035
rect 13599 25035 24179 25039
rect 13599 25032 13613 25035
rect 13620 25032 13623 25035
rect 13668 25015 13670 25035
rect 13716 25015 13718 25035
rect 13764 25015 13766 25035
rect 13860 25015 13862 25035
rect 13956 25015 13958 25035
rect 14004 25015 14006 25035
rect 14100 25015 14102 25035
rect 14940 25015 14942 25035
rect 15036 25015 15038 25035
rect 15180 25015 15182 25035
rect 15276 25015 15278 25035
rect 15420 25015 15422 25035
rect 15492 25015 15494 25035
rect 15660 25015 15662 25035
rect 15708 25015 15710 25035
rect 15732 25015 15734 25035
rect 15756 25015 15758 25035
rect 15804 25015 15806 25035
rect 15828 25015 15830 25035
rect 15852 25015 15854 25035
rect 15948 25015 15950 25035
rect 15972 25015 15974 25035
rect 16044 25015 16046 25035
rect 16068 25015 16070 25035
rect 16164 25015 16166 25035
rect 16260 25015 16262 25035
rect 16332 25015 16334 25035
rect 16548 25015 16550 25035
rect 16572 25015 16574 25035
rect 16620 25015 16622 25035
rect 16668 25015 16670 25035
rect 16716 25015 16718 25035
rect 16764 25015 16766 25035
rect 16812 25015 16814 25035
rect 16884 25015 16886 25035
rect 16908 25015 16910 25035
rect 16980 25015 16982 25035
rect 17148 25015 17150 25035
rect 17196 25015 17198 25035
rect 17220 25015 17222 25035
rect 17292 25015 17294 25035
rect 17316 25015 17318 25035
rect 18132 25015 18134 25035
rect 18228 25015 18230 25035
rect 18492 25015 18494 25035
rect 18516 25015 18518 25035
rect 18612 25015 18614 25035
rect 18828 25015 18830 25035
rect 18900 25015 18902 25035
rect 18924 25015 18926 25035
rect 18996 25015 18998 25035
rect 19020 25015 19022 25035
rect 19092 25015 19094 25035
rect 19140 25015 19142 25035
rect 19236 25015 19238 25035
rect 19260 25015 19262 25035
rect 19788 25015 19790 25035
rect 19836 25015 19838 25035
rect 19860 25015 19862 25035
rect 19884 25015 19886 25035
rect 19956 25015 19958 25035
rect 19980 25015 19982 25035
rect 20052 25015 20054 25035
rect 20076 25015 20078 25035
rect 20124 25015 20126 25035
rect 20172 25015 20174 25035
rect 20196 25015 20198 25035
rect 20292 25015 20294 25035
rect 20388 25015 20390 25035
rect 20412 25015 20414 25035
rect 20508 25015 20510 25035
rect 20532 25015 20534 25035
rect 20604 25015 20606 25035
rect 20628 25015 20630 25035
rect 20881 25030 20884 25035
rect 20891 25016 20894 25030
rect 20892 25015 20894 25016
rect 20964 25015 20966 25035
rect 21012 25032 21014 25035
rect 20988 25015 20991 25032
rect 21012 25015 21015 25032
rect 21108 25015 21110 25035
rect 21204 25015 21206 25035
rect 21300 25015 21302 25035
rect 21324 25015 21326 25035
rect 21444 25015 21446 25035
rect 21468 25015 21470 25035
rect 21564 25015 21566 25035
rect 21588 25015 21590 25035
rect 21684 25015 21686 25035
rect 21708 25015 21710 25035
rect 21828 25015 21830 25035
rect 21924 25015 21926 25035
rect 22068 25015 22070 25035
rect 22188 25015 22190 25035
rect 22212 25015 22214 25035
rect 22884 25015 22886 25035
rect 22980 25015 22982 25035
rect 23076 25015 23078 25035
rect 23100 25015 23102 25035
rect 23124 25015 23126 25035
rect 23244 25015 23246 25035
rect 23340 25015 23342 25035
rect 23412 25015 23414 25035
rect 23460 25015 23462 25035
rect 23508 25015 23510 25035
rect 23556 25015 23558 25035
rect 23604 25015 23606 25035
rect 23652 25015 23654 25035
rect 23676 25015 23678 25035
rect 23700 25015 23702 25035
rect 23772 25015 23774 25035
rect 23796 25015 23798 25035
rect 23916 25016 23918 25035
rect 24012 25016 24014 25035
rect 24049 25030 24052 25035
rect 24060 25030 24062 25035
rect 24145 25030 24148 25035
rect 24156 25032 24158 25035
rect 24156 25030 24159 25032
rect 24059 25016 24062 25030
rect 24155 25016 24159 25030
rect 23809 25015 23867 25016
rect 23905 25015 23939 25016
rect -12959 25011 -12331 25015
rect -12852 25008 -12850 25011
rect -12852 24992 -12849 25008
rect -12863 24991 -12829 24992
rect -12791 24991 -12757 24992
rect -12863 24987 -12757 24991
rect -12743 24991 -12709 24992
rect -12636 24991 -12634 25011
rect -12420 24991 -12418 25011
rect -12345 25008 -12331 25011
rect -12321 25011 12869 25015
rect -12321 25008 -12307 25011
rect -12300 25008 -12297 25011
rect -12095 25006 -12092 25011
rect -12085 24992 -12082 25006
rect -12084 24991 -12082 24992
rect -11772 24991 -11770 25011
rect -11676 24991 -11674 25011
rect -11652 24991 -11650 25011
rect -11508 24991 -11506 25011
rect -11436 24991 -11434 25011
rect -11412 24991 -11410 25011
rect -11196 24991 -11194 25011
rect -11100 24991 -11098 25011
rect -10809 25008 -10795 25011
rect -10764 24991 -10762 25011
rect -10644 24991 -10642 25011
rect -9900 24991 -9898 25011
rect -9732 24991 -9730 25011
rect -9444 24991 -9442 25011
rect -9348 24991 -9346 25011
rect -9228 24991 -9226 25011
rect -9108 24991 -9106 25011
rect -8436 24991 -8434 25011
rect -8364 24991 -8362 25011
rect -8340 24991 -8338 25011
rect -8268 24991 -8266 25011
rect -8124 24991 -8122 25011
rect -8028 24992 -8026 25011
rect -8039 24991 -8005 24992
rect -7932 24991 -7930 25011
rect -7764 24991 -7762 25011
rect -7524 24991 -7522 25011
rect -7356 24991 -7354 25011
rect -7308 24991 -7306 25011
rect -7212 24991 -7210 25011
rect -7044 24991 -7042 25011
rect -6948 24991 -6946 25011
rect -6852 24991 -6850 25011
rect -6767 25006 -6764 25011
rect -6756 25006 -6754 25011
rect -6743 25006 -6740 25011
rect -6660 25008 -6658 25011
rect -6612 25008 -6610 25011
rect -6757 24992 -6754 25006
rect -6733 24992 -6730 25006
rect -6732 24991 -6730 24992
rect -6660 24991 -6657 25008
rect -6612 24991 -6609 25008
rect -6516 24991 -6514 25011
rect -5892 24991 -5890 25011
rect -5436 24991 -5434 25011
rect -5340 24991 -5338 25011
rect -5196 24991 -5194 25011
rect -5100 24992 -5098 25011
rect -5111 24991 -5077 24992
rect -4716 24991 -4714 25011
rect -4500 24991 -4498 25011
rect -4404 24991 -4402 25011
rect -4308 24991 -4306 25011
rect -4164 24991 -4162 25011
rect -4127 24991 -4093 24992
rect -4020 24991 -4018 25011
rect -3876 24991 -3874 25011
rect -3732 24991 -3730 25011
rect -3636 24991 -3634 25011
rect -3540 24991 -3538 25011
rect -3468 24991 -3466 25011
rect -3324 24991 -3322 25011
rect -3108 24991 -3106 25011
rect -3012 24991 -3010 25011
rect -2964 24991 -2962 25011
rect -2916 24991 -2914 25011
rect -2892 24991 -2890 25011
rect -2868 24991 -2866 25011
rect -2820 24991 -2818 25011
rect -2772 24991 -2770 25011
rect -2676 24991 -2674 25011
rect -2364 24991 -2362 25011
rect -2316 24991 -2314 25011
rect -2076 24991 -2074 25011
rect -2052 25008 -2050 25011
rect -2052 24991 -2049 25008
rect -1980 24991 -1978 25011
rect -1895 25006 -1892 25011
rect -1884 25006 -1882 25011
rect -1885 24992 -1882 25006
rect -1812 24991 -1809 25008
rect -1572 24991 -1570 25011
rect -1476 24991 -1474 25011
rect -1356 24991 -1354 25011
rect -1260 24991 -1258 25011
rect -1236 24991 -1234 25011
rect -1140 24991 -1138 25011
rect -876 24991 -874 25011
rect -660 24991 -658 25011
rect -492 24991 -490 25011
rect -444 24991 -442 25011
rect -396 24991 -394 25011
rect -348 24991 -346 25011
rect -276 24991 -274 25011
rect -12 24991 -10 25011
rect 156 24991 158 25011
rect 204 24991 206 25011
rect 252 24991 254 25011
rect 348 24991 350 25011
rect 468 24991 470 25011
rect 492 24991 494 25011
rect 564 24991 566 25011
rect 588 24991 590 25011
rect 636 24991 638 25011
rect 660 24991 662 25011
rect 732 24991 734 25011
rect 1092 24991 1094 25011
rect 1140 24991 1142 25011
rect 1308 24991 1310 25011
rect 1356 24991 1358 25011
rect 1428 24991 1430 25011
rect 1692 24991 1694 25011
rect 1860 24991 1862 25011
rect 2017 25006 2020 25011
rect 2028 25006 2030 25011
rect 2027 24992 2030 25006
rect 2076 24991 2078 25011
rect 2100 24991 2102 25011
rect 2124 25008 2126 25011
rect 2124 24991 2127 25008
rect 2244 24991 2246 25011
rect 2401 25006 2404 25011
rect 2412 25008 2414 25011
rect 2412 25006 2415 25008
rect 2411 24992 2415 25006
rect 2460 24991 2462 25011
rect 2508 25008 2510 25011
rect 2508 24991 2511 25008
rect 2593 25006 2596 25011
rect 2604 25006 2606 25011
rect 2603 24992 2606 25006
rect 2772 24991 2774 25011
rect 2868 24991 2870 25011
rect 2940 24991 2942 25011
rect 3012 24991 3014 25011
rect 3108 24991 3110 25011
rect 3324 24991 3326 25011
rect 3396 24991 3398 25011
rect 3564 24991 3566 25011
rect 3625 25006 3628 25011
rect 3636 25006 3638 25011
rect 3635 24992 3638 25006
rect 3660 24991 3662 25011
rect 3732 25008 3734 25011
rect 3732 24991 3735 25008
rect 3780 24991 3782 25011
rect 3828 24992 3830 25011
rect 3924 24992 3926 25011
rect 3817 24991 3851 24992
rect 3913 24991 3947 24992
rect 4020 24991 4022 25011
rect 4092 24991 4094 25011
rect 4188 24991 4190 25011
rect 4308 24991 4310 25011
rect 4404 24991 4406 25011
rect 4500 24991 4502 25011
rect 4596 24991 4598 25011
rect 4692 24991 4694 25011
rect 4956 24991 4958 25011
rect 4980 24991 4982 25011
rect 5052 24991 5054 25011
rect 5124 24991 5126 25011
rect 5220 24991 5222 25011
rect 5268 24991 5270 25011
rect 5388 24991 5390 25011
rect 5484 24991 5486 25011
rect 5508 24991 5510 25011
rect 5532 24991 5534 25011
rect 5628 24991 5630 25011
rect 5652 24991 5654 25011
rect 5748 24991 5750 25011
rect 5796 24991 5798 25011
rect 5844 24991 5846 25011
rect 5892 24991 5894 25011
rect 6132 24991 6134 25011
rect 6228 24991 6230 25011
rect 6252 24991 6254 25011
rect 6276 24991 6278 25011
rect 6324 24991 6326 25011
rect 6372 24991 6374 25011
rect 6420 24991 6422 25011
rect 6492 24991 6494 25011
rect 6516 24991 6518 25011
rect 6588 24991 6590 25011
rect 6612 24991 6614 25011
rect 6649 25006 6652 25011
rect 6660 25006 6662 25011
rect 6659 24992 6662 25006
rect 6684 24991 6686 25011
rect 6708 24991 6710 25011
rect 6780 24991 6782 25011
rect 6804 24991 6806 25011
rect 6900 24991 6902 25011
rect 6924 24991 6926 25011
rect 7020 24991 7022 25011
rect 7164 24991 7166 25011
rect 7236 24991 7238 25011
rect 7308 24991 7310 25011
rect 7380 24991 7382 25011
rect 7404 24991 7406 25011
rect 7476 24991 7478 25011
rect 7572 24991 7574 25011
rect 7620 24991 7622 25011
rect 7644 24991 7646 25011
rect 7668 24991 7670 25011
rect 7849 24991 7883 24992
rect 7908 24991 7910 25011
rect 7956 24992 7958 25011
rect 7945 24991 7979 24992
rect 8124 24991 8126 25011
rect 8220 24991 8222 25011
rect 8652 24991 8654 25011
rect 8700 24991 8702 25011
rect 8748 24991 8750 25011
rect 8796 24991 8798 25011
rect 8844 24991 8846 25011
rect 8868 24991 8870 25011
rect 9516 24991 9518 25011
rect 9660 24991 9662 25011
rect 9684 24991 9686 25011
rect 9756 24991 9758 25011
rect 9780 24991 9782 25011
rect 9804 24991 9806 25011
rect 9852 24991 9854 25011
rect 9900 24991 9902 25011
rect 9948 24991 9950 25011
rect 10044 24991 10046 25011
rect 10116 24991 10118 25011
rect 10129 24991 10187 24992
rect 10188 24991 10190 25011
rect 10284 24991 10286 25011
rect 10332 24991 10334 25011
rect 10380 24991 10382 25011
rect 10428 24991 10430 25011
rect 10476 24991 10478 25011
rect 10524 24991 10526 25011
rect 10620 24991 10622 25011
rect 10644 24991 10646 25011
rect 10716 24991 10718 25011
rect 10956 24991 10958 25011
rect 11004 24991 11006 25011
rect 11052 24991 11054 25011
rect 11100 24991 11102 25011
rect 11172 24991 11174 25011
rect 11220 24991 11222 25011
rect 11340 24991 11342 25011
rect 11436 24991 11438 25011
rect 11532 24991 11534 25011
rect 11628 24991 11630 25011
rect 11676 24991 11678 25011
rect 11724 24991 11726 25011
rect 11772 24991 11774 25011
rect 11796 24991 11798 25011
rect 11892 24991 11894 25011
rect 11988 24991 11990 25011
rect 12060 24991 12062 25011
rect 12276 24991 12278 25011
rect 12324 24991 12326 25011
rect 12420 24991 12422 25011
rect 12444 24991 12446 25011
rect 12516 24991 12518 25011
rect 12540 24991 12542 25011
rect 12564 24991 12566 25011
rect 12660 24991 12662 25011
rect 12756 24991 12758 25011
rect 12828 24991 12830 25011
rect 12855 25008 12869 25011
rect 12876 25011 20981 25015
rect 12876 25008 12893 25011
rect 12876 24991 12878 25008
rect 12972 24991 12974 25011
rect 13044 24991 13046 25011
rect 13068 24991 13070 25011
rect 13116 24991 13118 25011
rect 13284 24991 13286 25011
rect 13332 24991 13334 25011
rect 13500 24991 13502 25011
rect 13572 24991 13574 25011
rect 13668 24991 13670 25011
rect 13716 24991 13718 25011
rect 13764 24991 13766 25011
rect 13860 24991 13862 25011
rect 13956 24991 13958 25011
rect 14004 24991 14006 25011
rect 14100 24991 14102 25011
rect 14940 24991 14942 25011
rect 15036 24991 15038 25011
rect 15180 24991 15182 25011
rect 15276 24991 15278 25011
rect 15420 24991 15422 25011
rect 15492 24991 15494 25011
rect 15660 24991 15662 25011
rect 15708 24991 15710 25011
rect 15732 24991 15734 25011
rect 15756 24991 15758 25011
rect 15804 24991 15806 25011
rect 15828 24991 15830 25011
rect 15852 24991 15854 25011
rect 15948 24991 15950 25011
rect 15972 24991 15974 25011
rect 16044 24991 16046 25011
rect 16068 24991 16070 25011
rect 16164 24991 16166 25011
rect 16260 24991 16262 25011
rect 16332 24991 16334 25011
rect 16548 24991 16550 25011
rect 16572 24991 16574 25011
rect 16620 24991 16622 25011
rect 16668 24991 16670 25011
rect 16716 24991 16718 25011
rect 16764 24991 16766 25011
rect 16812 24991 16814 25011
rect 16884 24991 16886 25011
rect 16908 24991 16910 25011
rect 16980 24991 16982 25011
rect 17148 24991 17150 25011
rect 17196 24991 17198 25011
rect 17220 24991 17222 25011
rect 17292 24991 17294 25011
rect 17316 24991 17318 25011
rect 18132 24991 18134 25011
rect 18228 24991 18230 25011
rect 18492 24991 18494 25011
rect 18516 24991 18518 25011
rect 18612 24991 18614 25011
rect 18828 24991 18830 25011
rect 18900 24991 18902 25011
rect 18924 24991 18926 25011
rect 18996 24991 18998 25011
rect 19020 24991 19022 25011
rect 19092 24991 19094 25011
rect 19140 24991 19142 25011
rect 19236 24991 19238 25011
rect 19260 24991 19262 25011
rect 19788 24991 19790 25011
rect 19836 24991 19838 25011
rect 19860 24991 19862 25011
rect 19884 24991 19886 25011
rect 19956 24991 19958 25011
rect 19980 24991 19982 25011
rect 20052 24991 20054 25011
rect 20076 24991 20078 25011
rect 20124 24991 20126 25011
rect 20172 24991 20174 25011
rect 20196 24991 20198 25011
rect 20292 24991 20294 25011
rect 20388 24991 20390 25011
rect 20412 24991 20414 25011
rect 20508 24991 20510 25011
rect 20532 24991 20534 25011
rect 20604 24991 20606 25011
rect 20628 24991 20630 25011
rect 20892 24991 20894 25011
rect 20964 24991 20966 25011
rect 20967 25008 20981 25011
rect 20988 25011 23939 25015
rect 23953 25015 23987 25016
rect 24001 25015 24035 25016
rect 23953 25011 24035 25015
rect 20988 25008 21005 25011
rect 21012 25008 21015 25011
rect 20988 24991 20990 25008
rect 21108 24991 21110 25011
rect 21204 24991 21206 25011
rect 21300 24991 21302 25011
rect 21324 24991 21326 25011
rect 21444 24991 21446 25011
rect 21468 24991 21470 25011
rect 21564 24991 21566 25011
rect 21588 24991 21590 25011
rect 21684 24991 21686 25011
rect 21708 24991 21710 25011
rect 21828 24991 21830 25011
rect 21924 24991 21926 25011
rect 22068 24991 22070 25011
rect 22188 24991 22190 25011
rect 22212 24991 22214 25011
rect 22884 24991 22886 25011
rect 22980 24991 22982 25011
rect 23076 24991 23078 25011
rect 23100 24991 23102 25011
rect 23124 24991 23126 25011
rect 23244 24991 23246 25011
rect 23340 24991 23342 25011
rect 23412 24991 23414 25011
rect 23460 24991 23462 25011
rect 23508 24991 23510 25011
rect 23556 24991 23558 25011
rect 23604 24991 23606 25011
rect 23652 24991 23654 25011
rect 23676 24991 23678 25011
rect 23700 24991 23702 25011
rect 23772 24991 23774 25011
rect 23796 24992 23798 25011
rect 23905 25006 23908 25011
rect 23916 25008 23918 25011
rect 23916 25006 23919 25008
rect 24001 25006 24004 25011
rect 24012 25008 24014 25011
rect 24012 25006 24015 25008
rect 23915 24998 23919 25006
rect 23929 24998 23933 25006
rect 23915 24992 23929 24998
rect 24011 24992 24015 25006
rect 23785 24991 23819 24992
rect -12743 24987 -11995 24991
rect -12863 24984 -12859 24987
rect -12852 24984 -12849 24987
rect -12636 24984 -12634 24987
rect -12767 24974 -12763 24982
rect -12777 24968 -12767 24974
rect -12636 24968 -12633 24984
rect -12647 24967 -12613 24968
rect -12455 24967 -12421 24968
rect -12420 24967 -12418 24987
rect -12084 24967 -12082 24987
rect -12009 24984 -11995 24987
rect -11985 24987 -6643 24991
rect -11985 24984 -11971 24987
rect -11772 24967 -11770 24987
rect -11676 24967 -11674 24987
rect -11652 24967 -11650 24987
rect -11508 24967 -11506 24987
rect -11436 24967 -11434 24987
rect -11412 24967 -11410 24987
rect -11196 24967 -11194 24987
rect -11100 24967 -11098 24987
rect -10764 24967 -10762 24987
rect -10644 24967 -10642 24987
rect -9900 24967 -9898 24987
rect -9732 24967 -9730 24987
rect -9647 24967 -9589 24968
rect -9444 24967 -9442 24987
rect -9348 24967 -9346 24987
rect -9228 24967 -9226 24987
rect -9108 24967 -9106 24987
rect -8436 24967 -8434 24987
rect -8364 24967 -8362 24987
rect -8340 24967 -8338 24987
rect -8268 24967 -8266 24987
rect -8124 24967 -8122 24987
rect -8039 24982 -8036 24987
rect -8028 24982 -8026 24987
rect -8029 24968 -8026 24982
rect -7932 24984 -7930 24987
rect -7932 24967 -7929 24984
rect -7764 24967 -7762 24987
rect -7524 24967 -7522 24987
rect -7497 24984 -7483 24987
rect -7356 24967 -7354 24987
rect -7308 24967 -7306 24987
rect -7212 24968 -7210 24987
rect -7247 24967 -7189 24968
rect -7044 24967 -7042 24987
rect -6948 24967 -6946 24987
rect -6852 24967 -6850 24987
rect -6732 24967 -6730 24987
rect -6681 24984 -6667 24987
rect -6660 24984 -6643 24987
rect -6633 24987 -1819 24991
rect -6633 24984 -6619 24987
rect -6612 24984 -6609 24987
rect -6516 24967 -6514 24987
rect -5892 24967 -5890 24987
rect -5436 24967 -5434 24987
rect -5340 24967 -5338 24987
rect -5196 24967 -5194 24987
rect -5111 24982 -5108 24987
rect -5100 24982 -5098 24987
rect -5101 24968 -5098 24982
rect -4716 24967 -4714 24987
rect -4500 24967 -4498 24987
rect -4404 24967 -4402 24987
rect -4308 24967 -4306 24987
rect -4164 24967 -4162 24987
rect -4020 24984 -4018 24987
rect -4020 24967 -4017 24984
rect -3876 24967 -3874 24987
rect -3732 24967 -3730 24987
rect -3636 24967 -3634 24987
rect -3540 24967 -3538 24987
rect -3468 24967 -3466 24987
rect -3324 24967 -3322 24987
rect -3108 24967 -3106 24987
rect -3012 24967 -3010 24987
rect -2964 24967 -2962 24987
rect -2916 24967 -2914 24987
rect -2892 24967 -2890 24987
rect -2868 24967 -2866 24987
rect -2820 24967 -2818 24987
rect -2772 24967 -2770 24987
rect -2676 24967 -2674 24987
rect -2364 24967 -2362 24987
rect -2316 24967 -2314 24987
rect -2076 24967 -2074 24987
rect -2073 24984 -2059 24987
rect -2052 24984 -2049 24987
rect -1980 24967 -1978 24987
rect -1833 24984 -1819 24987
rect -1812 24987 6725 24991
rect -1812 24984 -1795 24987
rect -1812 24967 -1810 24984
rect -1572 24967 -1570 24987
rect -1476 24967 -1474 24987
rect -1356 24967 -1354 24987
rect -1260 24967 -1258 24987
rect -1236 24967 -1234 24987
rect -1140 24967 -1138 24987
rect -876 24967 -874 24987
rect -660 24967 -658 24987
rect -492 24967 -490 24987
rect -444 24968 -442 24987
rect -479 24967 -421 24968
rect -396 24967 -394 24987
rect -348 24967 -346 24987
rect -276 24967 -274 24987
rect -12 24967 -10 24987
rect 156 24967 158 24987
rect 204 24967 206 24987
rect 252 24967 254 24987
rect 348 24967 350 24987
rect 468 24967 470 24987
rect 492 24967 494 24987
rect 564 24967 566 24987
rect 588 24967 590 24987
rect 636 24967 638 24987
rect 660 24967 662 24987
rect 732 24967 734 24987
rect 1092 24967 1094 24987
rect 1140 24967 1142 24987
rect 1308 24967 1310 24987
rect 1356 24967 1358 24987
rect 1428 24967 1430 24987
rect 1692 24967 1694 24987
rect 1860 24967 1862 24987
rect 2076 24967 2078 24987
rect 2100 24967 2102 24987
rect 2103 24984 2117 24987
rect 2124 24984 2127 24987
rect 2244 24967 2246 24987
rect 2391 24984 2405 24987
rect 2460 24967 2462 24987
rect 2487 24984 2501 24987
rect 2508 24984 2511 24987
rect 2679 24984 2693 24987
rect 2772 24967 2774 24987
rect 2868 24967 2870 24987
rect 2940 24967 2942 24987
rect 3012 24967 3014 24987
rect 3108 24967 3110 24987
rect 3324 24967 3326 24987
rect 3396 24967 3398 24987
rect 3564 24967 3566 24987
rect 3660 24967 3662 24987
rect 3711 24984 3725 24987
rect 3732 24984 3735 24987
rect 3780 24967 3782 24987
rect 3817 24982 3820 24987
rect 3828 24982 3830 24987
rect 3913 24982 3916 24987
rect 3924 24984 3926 24987
rect 4020 24984 4022 24987
rect 3924 24982 3927 24984
rect 3827 24968 3830 24982
rect 3923 24968 3927 24982
rect 4020 24967 4023 24984
rect 4092 24967 4094 24987
rect 4188 24967 4190 24987
rect 4308 24967 4310 24987
rect 4404 24967 4406 24987
rect 4500 24967 4502 24987
rect 4596 24967 4598 24987
rect 4692 24967 4694 24987
rect 4956 24967 4958 24987
rect 4980 24967 4982 24987
rect 5052 24967 5054 24987
rect 5124 24967 5126 24987
rect 5220 24967 5222 24987
rect 5268 24967 5270 24987
rect 5388 24967 5390 24987
rect 5484 24967 5486 24987
rect 5508 24967 5510 24987
rect 5532 24967 5534 24987
rect 5628 24967 5630 24987
rect 5652 24967 5654 24987
rect 5748 24967 5750 24987
rect 5796 24967 5798 24987
rect 5844 24967 5846 24987
rect 5892 24967 5894 24987
rect 6001 24967 6059 24968
rect 6132 24967 6134 24987
rect 6228 24967 6230 24987
rect 6252 24967 6254 24987
rect 6276 24967 6278 24987
rect 6324 24967 6326 24987
rect 6372 24967 6374 24987
rect 6420 24967 6422 24987
rect 6492 24967 6494 24987
rect 6516 24967 6518 24987
rect 6588 24967 6590 24987
rect 6612 24967 6614 24987
rect 6684 24967 6686 24987
rect 6708 24967 6710 24987
rect 6711 24984 6725 24987
rect 6735 24987 23819 24991
rect 6735 24984 6749 24987
rect 6780 24967 6782 24987
rect 6804 24967 6806 24987
rect 6900 24967 6902 24987
rect 6924 24967 6926 24987
rect 7020 24967 7022 24987
rect 7164 24967 7166 24987
rect 7236 24967 7238 24987
rect 7308 24967 7310 24987
rect 7380 24967 7382 24987
rect 7404 24967 7406 24987
rect 7476 24967 7478 24987
rect 7572 24967 7574 24987
rect 7620 24967 7622 24987
rect 7644 24967 7646 24987
rect 7668 24967 7670 24987
rect 7908 24967 7910 24987
rect 7945 24982 7948 24987
rect 7956 24984 7958 24987
rect 7956 24982 7959 24984
rect 7955 24968 7959 24982
rect 8124 24967 8126 24987
rect 8220 24967 8222 24987
rect 8652 24967 8654 24987
rect 8700 24967 8702 24987
rect 8748 24967 8750 24987
rect 8796 24967 8798 24987
rect 8844 24967 8846 24987
rect 8868 24967 8870 24987
rect 9516 24967 9518 24987
rect 9660 24967 9662 24987
rect 9684 24967 9686 24987
rect 9756 24967 9758 24987
rect 9780 24967 9782 24987
rect 9804 24967 9806 24987
rect 9852 24967 9854 24987
rect 9900 24968 9902 24987
rect 9889 24967 9923 24968
rect 9948 24967 9950 24987
rect 10044 24967 10046 24987
rect 10116 24967 10118 24987
rect 10129 24982 10132 24987
rect 10139 24968 10142 24982
rect 10140 24967 10142 24968
rect 10188 24967 10190 24987
rect 10236 24967 10239 24984
rect 10284 24967 10286 24987
rect 10332 24967 10334 24987
rect 10380 24967 10382 24987
rect 10428 24967 10430 24987
rect 10476 24967 10478 24987
rect 10524 24967 10526 24987
rect 10620 24967 10622 24987
rect 10644 24967 10646 24987
rect 10716 24967 10718 24987
rect 10956 24967 10958 24987
rect 11004 24967 11006 24987
rect 11052 24967 11054 24987
rect 11100 24967 11102 24987
rect 11172 24967 11174 24987
rect 11220 24967 11222 24987
rect 11340 24967 11342 24987
rect 11436 24967 11438 24987
rect 11532 24967 11534 24987
rect 11628 24967 11630 24987
rect 11676 24967 11678 24987
rect 11724 24967 11726 24987
rect 11772 24967 11774 24987
rect 11796 24967 11798 24987
rect 11892 24967 11894 24987
rect 11988 24967 11990 24987
rect 12060 24967 12062 24987
rect 12276 24967 12278 24987
rect 12324 24967 12326 24987
rect 12361 24967 12419 24968
rect 12420 24967 12422 24987
rect 12444 24967 12446 24987
rect 12516 24967 12518 24987
rect 12540 24967 12542 24987
rect 12564 24967 12566 24987
rect 12660 24967 12662 24987
rect 12756 24967 12758 24987
rect 12828 24967 12830 24987
rect 12876 24967 12878 24987
rect 12972 24967 12974 24987
rect 13044 24967 13046 24987
rect 13068 24967 13070 24987
rect 13116 24967 13118 24987
rect 13284 24967 13286 24987
rect 13332 24967 13334 24987
rect 13500 24967 13502 24987
rect 13572 24967 13574 24987
rect 13668 24967 13670 24987
rect 13716 24967 13718 24987
rect 13764 24967 13766 24987
rect 13860 24967 13862 24987
rect 13956 24967 13958 24987
rect 14004 24967 14006 24987
rect 14100 24967 14102 24987
rect 14940 24967 14942 24987
rect 15036 24967 15038 24987
rect 15180 24967 15182 24987
rect 15276 24967 15278 24987
rect 15420 24967 15422 24987
rect 15492 24967 15494 24987
rect 15660 24967 15662 24987
rect 15708 24967 15710 24987
rect 15732 24967 15734 24987
rect 15756 24967 15758 24987
rect 15804 24967 15806 24987
rect 15828 24967 15830 24987
rect 15852 24967 15854 24987
rect 15948 24967 15950 24987
rect 15972 24967 15974 24987
rect 16044 24967 16046 24987
rect 16068 24967 16070 24987
rect 16164 24967 16166 24987
rect 16260 24967 16262 24987
rect 16332 24967 16334 24987
rect 16548 24967 16550 24987
rect 16572 24967 16574 24987
rect 16620 24967 16622 24987
rect 16668 24967 16670 24987
rect 16716 24967 16718 24987
rect 16764 24967 16766 24987
rect 16812 24967 16814 24987
rect 16884 24967 16886 24987
rect 16908 24967 16910 24987
rect 16980 24967 16982 24987
rect 17148 24967 17150 24987
rect 17196 24967 17198 24987
rect 17220 24967 17222 24987
rect 17292 24967 17294 24987
rect 17316 24967 17318 24987
rect 18132 24967 18134 24987
rect 18228 24967 18230 24987
rect 18492 24967 18494 24987
rect 18516 24967 18518 24987
rect 18612 24967 18614 24987
rect 18625 24967 18683 24968
rect 18828 24967 18830 24987
rect 18900 24967 18902 24987
rect 18924 24967 18926 24987
rect 18996 24967 18998 24987
rect 19020 24967 19022 24987
rect 19092 24967 19094 24987
rect 19140 24967 19142 24987
rect 19236 24967 19238 24987
rect 19260 24967 19262 24987
rect 19788 24967 19790 24987
rect 19836 24967 19838 24987
rect 19860 24967 19862 24987
rect 19884 24967 19886 24987
rect 19956 24967 19958 24987
rect 19980 24967 19982 24987
rect 20052 24967 20054 24987
rect 20076 24967 20078 24987
rect 20124 24967 20126 24987
rect 20172 24967 20174 24987
rect 20196 24967 20198 24987
rect 20292 24967 20294 24987
rect 20388 24967 20390 24987
rect 20412 24967 20414 24987
rect 20508 24967 20510 24987
rect 20532 24967 20534 24987
rect 20604 24967 20606 24987
rect 20628 24967 20630 24987
rect 20892 24967 20894 24987
rect 20964 24967 20966 24987
rect 20988 24967 20990 24987
rect 21108 24967 21110 24987
rect 21204 24967 21206 24987
rect 21300 24967 21302 24987
rect 21324 24967 21326 24987
rect 21444 24967 21446 24987
rect 21468 24967 21470 24987
rect 21564 24967 21566 24987
rect 21588 24967 21590 24987
rect 21684 24967 21686 24987
rect 21708 24967 21710 24987
rect 21828 24967 21830 24987
rect 21924 24967 21926 24987
rect 22068 24967 22070 24987
rect 22188 24967 22190 24987
rect 22212 24967 22214 24987
rect 22884 24967 22886 24987
rect 22980 24967 22982 24987
rect 23076 24967 23078 24987
rect 23100 24967 23102 24987
rect 23124 24967 23126 24987
rect 23244 24967 23246 24987
rect 23340 24967 23342 24987
rect 23412 24967 23414 24987
rect 23460 24967 23462 24987
rect 23508 24967 23510 24987
rect 23556 24967 23558 24987
rect 23604 24967 23606 24987
rect 23652 24967 23654 24987
rect 23676 24968 23678 24987
rect 23700 24968 23702 24987
rect 23772 24968 23774 24987
rect 23785 24982 23788 24987
rect 23796 24982 23798 24987
rect 23795 24968 23798 24982
rect 23665 24967 23723 24968
rect 23761 24967 23795 24968
rect -12647 24963 10229 24967
rect -12647 24960 -12643 24963
rect -12636 24960 -12633 24963
rect -12527 24943 -12493 24944
rect -12420 24943 -12418 24963
rect -12084 24943 -12082 24963
rect -11903 24943 -11869 24944
rect -11772 24943 -11770 24963
rect -11676 24943 -11674 24963
rect -11652 24943 -11650 24963
rect -11508 24943 -11506 24963
rect -11436 24943 -11434 24963
rect -11412 24943 -11410 24963
rect -11196 24943 -11194 24963
rect -11100 24943 -11098 24963
rect -10764 24944 -10762 24963
rect -10644 24944 -10642 24963
rect -10775 24943 -10741 24944
rect -10655 24943 -10621 24944
rect -9900 24943 -9898 24963
rect -9732 24943 -9730 24963
rect -9647 24958 -9644 24963
rect -9637 24944 -9634 24958
rect -9636 24943 -9634 24944
rect -9540 24943 -9537 24960
rect -9444 24943 -9442 24963
rect -9348 24943 -9346 24963
rect -9228 24943 -9226 24963
rect -9108 24943 -9106 24963
rect -8639 24943 -8581 24944
rect -8436 24943 -8434 24963
rect -8364 24943 -8362 24963
rect -8340 24943 -8338 24963
rect -8268 24943 -8266 24963
rect -8124 24943 -8122 24963
rect -7953 24960 -7939 24963
rect -7932 24960 -7929 24963
rect -7764 24943 -7762 24963
rect -7524 24943 -7522 24963
rect -7356 24943 -7354 24963
rect -7308 24943 -7306 24963
rect -7223 24958 -7220 24963
rect -7212 24958 -7210 24963
rect -7213 24944 -7210 24958
rect -7140 24943 -7137 24960
rect -7044 24943 -7042 24963
rect -6948 24943 -6946 24963
rect -6852 24943 -6850 24963
rect -6732 24943 -6730 24963
rect -6516 24943 -6514 24963
rect -5892 24943 -5890 24963
rect -5436 24943 -5434 24963
rect -5375 24943 -5341 24944
rect -5340 24943 -5338 24963
rect -5196 24943 -5194 24963
rect -5025 24960 -5011 24963
rect -4716 24943 -4714 24963
rect -4500 24943 -4498 24963
rect -4404 24943 -4402 24963
rect -4308 24943 -4306 24963
rect -4164 24943 -4162 24963
rect -4041 24960 -4027 24963
rect -4020 24960 -4017 24963
rect -3876 24943 -3874 24963
rect -3732 24943 -3730 24963
rect -3636 24943 -3634 24963
rect -3540 24943 -3538 24963
rect -3468 24943 -3466 24963
rect -3324 24943 -3322 24963
rect -3108 24943 -3106 24963
rect -3012 24943 -3010 24963
rect -2964 24943 -2962 24963
rect -2916 24943 -2914 24963
rect -2892 24944 -2890 24963
rect -2903 24943 -2869 24944
rect -2868 24943 -2866 24963
rect -2820 24943 -2818 24963
rect -2772 24943 -2770 24963
rect -2676 24943 -2674 24963
rect -2364 24943 -2362 24963
rect -2316 24943 -2314 24963
rect -2076 24943 -2074 24963
rect -1980 24943 -1978 24963
rect -1812 24943 -1810 24963
rect -1572 24943 -1570 24963
rect -1476 24943 -1474 24963
rect -1356 24943 -1354 24963
rect -1260 24943 -1258 24963
rect -1236 24943 -1234 24963
rect -1140 24943 -1138 24963
rect -876 24943 -874 24963
rect -660 24943 -658 24963
rect -492 24943 -490 24963
rect -455 24958 -452 24963
rect -444 24958 -442 24963
rect -445 24944 -442 24958
rect -396 24943 -394 24963
rect -348 24960 -346 24963
rect -372 24943 -369 24960
rect -348 24943 -345 24960
rect -276 24943 -274 24963
rect -12 24943 -10 24963
rect 156 24943 158 24963
rect 204 24943 206 24963
rect 252 24943 254 24963
rect 348 24943 350 24963
rect 468 24943 470 24963
rect 492 24943 494 24963
rect 564 24943 566 24963
rect 588 24943 590 24963
rect 636 24943 638 24963
rect 660 24943 662 24963
rect 732 24943 734 24963
rect 1092 24943 1094 24963
rect 1140 24943 1142 24963
rect 1308 24943 1310 24963
rect 1356 24943 1358 24963
rect 1428 24943 1430 24963
rect 1692 24943 1694 24963
rect 1860 24943 1862 24963
rect 2076 24943 2078 24963
rect 2100 24943 2102 24963
rect 2244 24943 2246 24963
rect 2460 24943 2462 24963
rect 2772 24943 2774 24963
rect 2868 24943 2870 24963
rect 2940 24943 2942 24963
rect 3012 24943 3014 24963
rect 3108 24943 3110 24963
rect 3324 24943 3326 24963
rect 3396 24943 3398 24963
rect 3564 24943 3566 24963
rect 3660 24943 3662 24963
rect 3780 24943 3782 24963
rect 3903 24960 3917 24963
rect 3999 24960 4013 24963
rect 4020 24960 4023 24963
rect 4092 24943 4094 24963
rect 4188 24943 4190 24963
rect 4308 24943 4310 24963
rect 4404 24943 4406 24963
rect 4500 24943 4502 24963
rect 4596 24943 4598 24963
rect 4692 24943 4694 24963
rect 4956 24943 4958 24963
rect 4980 24943 4982 24963
rect 5052 24943 5054 24963
rect 5124 24943 5126 24963
rect 5220 24943 5222 24963
rect 5268 24943 5270 24963
rect 5388 24943 5390 24963
rect 5484 24943 5486 24963
rect 5508 24943 5510 24963
rect 5532 24943 5534 24963
rect 5628 24943 5630 24963
rect 5652 24943 5654 24963
rect 5748 24943 5750 24963
rect 5796 24943 5798 24963
rect 5844 24943 5846 24963
rect 5892 24943 5894 24963
rect 6132 24960 6134 24963
rect 6132 24943 6135 24960
rect 6228 24943 6230 24963
rect 6252 24944 6254 24963
rect 6241 24943 6275 24944
rect 6276 24943 6278 24963
rect 6324 24943 6326 24963
rect 6372 24943 6374 24963
rect 6420 24943 6422 24963
rect 6492 24943 6494 24963
rect 6516 24943 6518 24963
rect 6588 24943 6590 24963
rect 6612 24943 6614 24963
rect 6684 24943 6686 24963
rect 6708 24943 6710 24963
rect 6780 24943 6782 24963
rect 6804 24943 6806 24963
rect 6900 24943 6902 24963
rect 6924 24943 6926 24963
rect 7020 24943 7022 24963
rect 7164 24943 7166 24963
rect 7236 24943 7238 24963
rect 7308 24943 7310 24963
rect 7380 24943 7382 24963
rect 7404 24943 7406 24963
rect 7476 24943 7478 24963
rect 7572 24943 7574 24963
rect 7620 24943 7622 24963
rect 7644 24943 7646 24963
rect 7668 24943 7670 24963
rect 7908 24943 7910 24963
rect 7935 24960 7949 24963
rect 8031 24960 8045 24963
rect 8124 24943 8126 24963
rect 8220 24943 8222 24963
rect 8652 24943 8654 24963
rect 8700 24943 8702 24963
rect 8748 24943 8750 24963
rect 8796 24943 8798 24963
rect 8844 24943 8846 24963
rect 8868 24943 8870 24963
rect 9516 24943 9518 24963
rect 9660 24943 9662 24963
rect 9684 24943 9686 24963
rect 9756 24943 9758 24963
rect 9780 24943 9782 24963
rect 9804 24943 9806 24963
rect 9852 24943 9854 24963
rect 9889 24958 9892 24963
rect 9900 24958 9902 24963
rect 9899 24944 9902 24958
rect 9948 24943 9950 24963
rect 10044 24943 10046 24963
rect 10116 24943 10118 24963
rect 10140 24943 10142 24963
rect 10188 24943 10190 24963
rect 10215 24960 10229 24963
rect 10236 24963 23795 24967
rect 10236 24960 10253 24963
rect 10236 24943 10238 24960
rect 10284 24943 10286 24963
rect 10332 24943 10334 24963
rect 10380 24943 10382 24963
rect 10428 24943 10430 24963
rect 10476 24943 10478 24963
rect 10524 24943 10526 24963
rect 10620 24943 10622 24963
rect 10644 24943 10646 24963
rect 10716 24943 10718 24963
rect 10956 24943 10958 24963
rect 11004 24943 11006 24963
rect 11052 24943 11054 24963
rect 11100 24943 11102 24963
rect 11172 24943 11174 24963
rect 11220 24943 11222 24963
rect 11340 24943 11342 24963
rect 11436 24943 11438 24963
rect 11532 24943 11534 24963
rect 11628 24943 11630 24963
rect 11676 24943 11678 24963
rect 11724 24943 11726 24963
rect 11772 24943 11774 24963
rect 11796 24943 11798 24963
rect 11892 24943 11894 24963
rect 11988 24943 11990 24963
rect 12060 24943 12062 24963
rect 12276 24943 12278 24963
rect 12324 24943 12326 24963
rect 12361 24958 12364 24963
rect 12371 24944 12374 24958
rect 12372 24943 12374 24944
rect 12420 24943 12422 24963
rect 12444 24943 12446 24963
rect 12468 24943 12471 24960
rect 12516 24943 12518 24963
rect 12540 24943 12542 24963
rect 12564 24943 12566 24963
rect 12660 24943 12662 24963
rect 12756 24943 12758 24963
rect 12828 24943 12830 24963
rect 12876 24943 12878 24963
rect 12972 24943 12974 24963
rect 12985 24943 13043 24944
rect 13044 24943 13046 24963
rect 13068 24943 13070 24963
rect 13116 24943 13118 24963
rect 13284 24943 13286 24963
rect 13332 24943 13334 24963
rect 13500 24943 13502 24963
rect 13572 24943 13574 24963
rect 13668 24943 13670 24963
rect 13716 24943 13718 24963
rect 13764 24943 13766 24963
rect 13860 24943 13862 24963
rect 13956 24943 13958 24963
rect 14004 24943 14006 24963
rect 14100 24943 14102 24963
rect 14940 24943 14942 24963
rect 15036 24943 15038 24963
rect 15180 24943 15182 24963
rect 15276 24943 15278 24963
rect 15420 24943 15422 24963
rect 15492 24943 15494 24963
rect 15660 24943 15662 24963
rect 15708 24943 15710 24963
rect 15732 24943 15734 24963
rect 15756 24943 15758 24963
rect 15804 24943 15806 24963
rect 15828 24943 15830 24963
rect 15852 24943 15854 24963
rect 15948 24943 15950 24963
rect 15972 24943 15974 24963
rect 16044 24943 16046 24963
rect 16068 24943 16070 24963
rect 16164 24943 16166 24963
rect 16260 24943 16262 24963
rect 16332 24943 16334 24963
rect 16548 24943 16550 24963
rect 16572 24943 16574 24963
rect 16620 24943 16622 24963
rect 16668 24943 16670 24963
rect 16716 24943 16718 24963
rect 16764 24943 16766 24963
rect 16812 24943 16814 24963
rect 16884 24943 16886 24963
rect 16908 24943 16910 24963
rect 16980 24943 16982 24963
rect 17148 24943 17150 24963
rect 17196 24943 17198 24963
rect 17220 24943 17222 24963
rect 17292 24943 17294 24963
rect 17316 24943 17318 24963
rect 18132 24943 18134 24963
rect 18228 24943 18230 24963
rect 18492 24943 18494 24963
rect 18516 24943 18518 24963
rect 18612 24943 18614 24963
rect 18625 24958 18628 24963
rect 18635 24944 18638 24958
rect 18636 24943 18638 24944
rect 18732 24943 18735 24960
rect 18828 24943 18830 24963
rect 18900 24943 18902 24963
rect 18924 24943 18926 24963
rect 18996 24944 18998 24963
rect 18961 24943 19019 24944
rect 19020 24943 19022 24963
rect 19092 24943 19094 24963
rect 19140 24943 19142 24963
rect 19236 24943 19238 24963
rect 19260 24943 19262 24963
rect 19788 24943 19790 24963
rect 19836 24943 19838 24963
rect 19860 24943 19862 24963
rect 19884 24943 19886 24963
rect 19956 24943 19958 24963
rect 19980 24943 19982 24963
rect 20052 24943 20054 24963
rect 20076 24943 20078 24963
rect 20124 24943 20126 24963
rect 20172 24943 20174 24963
rect 20196 24943 20198 24963
rect 20292 24943 20294 24963
rect 20388 24943 20390 24963
rect 20412 24943 20414 24963
rect 20508 24943 20510 24963
rect 20532 24943 20534 24963
rect 20604 24943 20606 24963
rect 20628 24943 20630 24963
rect 20892 24943 20894 24963
rect 20964 24943 20966 24963
rect 20988 24943 20990 24963
rect 21108 24943 21110 24963
rect 21204 24943 21206 24963
rect 21300 24943 21302 24963
rect 21324 24943 21326 24963
rect 21444 24943 21446 24963
rect 21468 24943 21470 24963
rect 21564 24943 21566 24963
rect 21588 24943 21590 24963
rect 21684 24943 21686 24963
rect 21708 24943 21710 24963
rect 21828 24943 21830 24963
rect 21924 24943 21926 24963
rect 22068 24943 22070 24963
rect 22188 24943 22190 24963
rect 22212 24943 22214 24963
rect 22884 24943 22886 24963
rect 22980 24943 22982 24963
rect 23076 24943 23078 24963
rect 23100 24943 23102 24963
rect 23124 24943 23126 24963
rect 23244 24943 23246 24963
rect 23340 24943 23342 24963
rect 23412 24943 23414 24963
rect 23460 24943 23462 24963
rect 23508 24943 23510 24963
rect 23556 24943 23558 24963
rect 23604 24944 23606 24963
rect 23652 24944 23654 24963
rect 23665 24958 23668 24963
rect 23676 24958 23678 24963
rect 23689 24958 23692 24963
rect 23700 24958 23702 24963
rect 23761 24958 23764 24963
rect 23772 24960 23774 24963
rect 23772 24958 23775 24960
rect 23675 24944 23678 24958
rect 23699 24944 23702 24958
rect 23771 24950 23775 24958
rect 23785 24950 23789 24958
rect 23771 24944 23785 24950
rect 23569 24943 23627 24944
rect 23641 24943 23675 24944
rect -12527 24939 -9547 24943
rect -12420 24936 -12418 24939
rect -12369 24936 -12355 24939
rect -12420 24920 -12417 24936
rect -12431 24919 -12397 24920
rect -12084 24919 -12082 24939
rect -11772 24919 -11770 24939
rect -11676 24919 -11674 24939
rect -11652 24920 -11650 24939
rect -11663 24919 -11629 24920
rect -11508 24919 -11506 24939
rect -11436 24919 -11434 24939
rect -11412 24919 -11410 24939
rect -11196 24919 -11194 24939
rect -11100 24919 -11098 24939
rect -10775 24934 -10772 24939
rect -10764 24934 -10762 24939
rect -10655 24934 -10652 24939
rect -10644 24934 -10642 24939
rect -10765 24920 -10762 24934
rect -10645 24920 -10642 24934
rect -9900 24919 -9898 24939
rect -9732 24919 -9730 24939
rect -9636 24919 -9634 24939
rect -9561 24936 -9547 24939
rect -9540 24939 -7147 24943
rect -9540 24936 -9523 24939
rect -9540 24919 -9538 24936
rect -9444 24919 -9442 24939
rect -9348 24919 -9346 24939
rect -9228 24919 -9226 24939
rect -9108 24919 -9106 24939
rect -8639 24934 -8636 24939
rect -8629 24920 -8626 24934
rect -9023 24919 -8965 24920
rect -8628 24919 -8626 24920
rect -8532 24919 -8529 24936
rect -8436 24919 -8434 24939
rect -8364 24919 -8362 24939
rect -8340 24919 -8338 24939
rect -8268 24919 -8266 24939
rect -8124 24919 -8122 24939
rect -7764 24919 -7762 24939
rect -7524 24919 -7522 24939
rect -7356 24919 -7354 24939
rect -7308 24919 -7306 24939
rect -7161 24936 -7147 24939
rect -7140 24939 -379 24943
rect -7140 24936 -7123 24939
rect -7140 24919 -7138 24936
rect -7044 24919 -7042 24939
rect -6948 24919 -6946 24939
rect -6852 24919 -6850 24939
rect -6732 24919 -6730 24939
rect -6516 24919 -6514 24939
rect -5892 24919 -5890 24939
rect -5436 24919 -5434 24939
rect -5340 24919 -5338 24939
rect -5196 24919 -5194 24939
rect -4716 24919 -4714 24939
rect -4500 24919 -4498 24939
rect -4404 24919 -4402 24939
rect -4308 24919 -4306 24939
rect -4164 24919 -4162 24939
rect -3876 24919 -3874 24939
rect -3732 24920 -3730 24939
rect -3767 24919 -3709 24920
rect -3636 24919 -3634 24939
rect -3540 24919 -3538 24939
rect -3468 24919 -3466 24939
rect -3324 24919 -3322 24939
rect -3108 24919 -3106 24939
rect -3012 24919 -3010 24939
rect -2964 24919 -2962 24939
rect -2916 24919 -2914 24939
rect -2903 24934 -2900 24939
rect -2892 24934 -2890 24939
rect -2893 24920 -2890 24934
rect -2868 24919 -2866 24939
rect -2820 24919 -2818 24939
rect -2772 24919 -2770 24939
rect -2676 24919 -2674 24939
rect -2364 24919 -2362 24939
rect -2316 24919 -2314 24939
rect -2076 24919 -2074 24939
rect -1980 24919 -1978 24939
rect -1812 24919 -1810 24939
rect -1572 24919 -1570 24939
rect -1476 24919 -1474 24939
rect -1356 24919 -1354 24939
rect -1260 24919 -1258 24939
rect -1236 24919 -1234 24939
rect -1140 24919 -1138 24939
rect -876 24919 -874 24939
rect -660 24919 -658 24939
rect -492 24919 -490 24939
rect -396 24919 -394 24939
rect -393 24936 -379 24939
rect -372 24939 6101 24943
rect -372 24936 -355 24939
rect -348 24936 -345 24939
rect -372 24919 -370 24936
rect -276 24919 -274 24939
rect -12 24919 -10 24939
rect 73 24919 131 24920
rect 156 24919 158 24939
rect 204 24919 206 24939
rect 252 24919 254 24939
rect 348 24919 350 24939
rect 468 24919 470 24939
rect 492 24919 494 24939
rect 564 24919 566 24939
rect 588 24919 590 24939
rect 636 24919 638 24939
rect 660 24919 662 24939
rect 732 24919 734 24939
rect 1092 24919 1094 24939
rect 1140 24919 1142 24939
rect 1308 24919 1310 24939
rect 1356 24919 1358 24939
rect 1428 24919 1430 24939
rect 1692 24919 1694 24939
rect 1860 24919 1862 24939
rect 2076 24919 2078 24939
rect 2100 24919 2102 24939
rect 2244 24919 2246 24939
rect 2460 24919 2462 24939
rect 2772 24919 2774 24939
rect 2868 24919 2870 24939
rect 2940 24919 2942 24939
rect 3012 24919 3014 24939
rect 3108 24919 3110 24939
rect 3324 24919 3326 24939
rect 3396 24919 3398 24939
rect 3564 24919 3566 24939
rect 3660 24919 3662 24939
rect 3780 24919 3782 24939
rect 4092 24919 4094 24939
rect 4188 24919 4190 24939
rect 4308 24919 4310 24939
rect 4404 24919 4406 24939
rect 4500 24919 4502 24939
rect 4596 24919 4598 24939
rect 4692 24919 4694 24939
rect 4956 24919 4958 24939
rect 4980 24919 4982 24939
rect 5052 24919 5054 24939
rect 5124 24919 5126 24939
rect 5220 24919 5222 24939
rect 5268 24919 5270 24939
rect 5388 24919 5390 24939
rect 5484 24919 5486 24939
rect 5508 24919 5510 24939
rect 5532 24919 5534 24939
rect 5628 24919 5630 24939
rect 5652 24919 5654 24939
rect 5748 24919 5750 24939
rect 5796 24919 5798 24939
rect 5844 24919 5846 24939
rect 5892 24919 5894 24939
rect 6087 24936 6101 24939
rect 6111 24939 12461 24943
rect 6111 24936 6125 24939
rect 6132 24936 6135 24939
rect 6228 24920 6230 24939
rect 6241 24934 6244 24939
rect 6252 24934 6254 24939
rect 6251 24920 6254 24934
rect 6193 24919 6251 24920
rect 6276 24919 6278 24939
rect 6324 24919 6326 24939
rect 6372 24919 6374 24939
rect 6420 24919 6422 24939
rect 6492 24919 6494 24939
rect 6516 24919 6518 24939
rect 6588 24919 6590 24939
rect 6612 24919 6614 24939
rect 6684 24919 6686 24939
rect 6708 24919 6710 24939
rect 6780 24919 6782 24939
rect 6804 24919 6806 24939
rect 6900 24919 6902 24939
rect 6924 24919 6926 24939
rect 7020 24919 7022 24939
rect 7164 24919 7166 24939
rect 7236 24919 7238 24939
rect 7308 24919 7310 24939
rect 7380 24919 7382 24939
rect 7404 24919 7406 24939
rect 7476 24919 7478 24939
rect 7572 24919 7574 24939
rect 7620 24919 7622 24939
rect 7644 24919 7646 24939
rect 7668 24919 7670 24939
rect 7908 24919 7910 24939
rect 8124 24919 8126 24939
rect 8220 24919 8222 24939
rect 8652 24919 8654 24939
rect 8700 24919 8702 24939
rect 8748 24919 8750 24939
rect 8796 24919 8798 24939
rect 8844 24919 8846 24939
rect 8868 24919 8870 24939
rect 9516 24919 9518 24939
rect 9660 24919 9662 24939
rect 9684 24919 9686 24939
rect 9756 24919 9758 24939
rect 9780 24919 9782 24939
rect 9804 24919 9806 24939
rect 9852 24919 9854 24939
rect 9948 24919 9950 24939
rect 9975 24936 9989 24939
rect 10044 24919 10046 24939
rect 10116 24919 10118 24939
rect 10140 24919 10142 24939
rect 10188 24919 10190 24939
rect 10236 24919 10238 24939
rect 10284 24919 10286 24939
rect 10332 24919 10334 24939
rect 10380 24919 10382 24939
rect 10428 24919 10430 24939
rect 10476 24919 10478 24939
rect 10524 24919 10526 24939
rect 10620 24919 10622 24939
rect 10644 24919 10646 24939
rect 10716 24919 10718 24939
rect 10873 24919 10931 24920
rect 10956 24919 10958 24939
rect 11004 24919 11006 24939
rect 11052 24919 11054 24939
rect 11100 24919 11102 24939
rect 11172 24919 11174 24939
rect 11220 24919 11222 24939
rect 11340 24919 11342 24939
rect 11436 24919 11438 24939
rect 11532 24919 11534 24939
rect 11628 24919 11630 24939
rect 11676 24919 11678 24939
rect 11724 24919 11726 24939
rect 11772 24919 11774 24939
rect 11796 24919 11798 24939
rect 11892 24919 11894 24939
rect 11988 24919 11990 24939
rect 12060 24919 12062 24939
rect 12276 24919 12278 24939
rect 12324 24919 12326 24939
rect 12372 24919 12374 24939
rect 12420 24919 12422 24939
rect 12444 24919 12446 24939
rect 12447 24936 12461 24939
rect 12468 24939 18725 24943
rect 12468 24936 12485 24939
rect 12468 24919 12470 24936
rect 12516 24919 12518 24939
rect 12540 24919 12542 24939
rect 12564 24919 12566 24939
rect 12660 24919 12662 24939
rect 12756 24919 12758 24939
rect 12828 24919 12830 24939
rect 12876 24919 12878 24939
rect 12972 24919 12974 24939
rect 13044 24919 13046 24939
rect 13068 24919 13070 24939
rect 13116 24936 13118 24939
rect 13116 24919 13119 24936
rect 13284 24919 13286 24939
rect 13332 24919 13334 24939
rect 13500 24919 13502 24939
rect 13572 24919 13574 24939
rect 13668 24919 13670 24939
rect 13716 24919 13718 24939
rect 13764 24919 13766 24939
rect 13860 24919 13862 24939
rect 13956 24919 13958 24939
rect 14004 24919 14006 24939
rect 14100 24919 14102 24939
rect 14940 24919 14942 24939
rect 15036 24919 15038 24939
rect 15180 24919 15182 24939
rect 15276 24919 15278 24939
rect 15420 24919 15422 24939
rect 15492 24919 15494 24939
rect 15660 24919 15662 24939
rect 15708 24919 15710 24939
rect 15732 24919 15734 24939
rect 15756 24919 15758 24939
rect 15804 24919 15806 24939
rect 15828 24919 15830 24939
rect 15852 24919 15854 24939
rect 15948 24919 15950 24939
rect 15972 24919 15974 24939
rect 16044 24919 16046 24939
rect 16068 24919 16070 24939
rect 16164 24919 16166 24939
rect 16260 24919 16262 24939
rect 16332 24919 16334 24939
rect 16369 24919 16427 24920
rect 16548 24919 16550 24939
rect 16572 24919 16574 24939
rect 16620 24919 16622 24939
rect 16668 24919 16670 24939
rect 16716 24919 16718 24939
rect 16764 24919 16766 24939
rect 16812 24919 16814 24939
rect 16884 24919 16886 24939
rect 16908 24919 16910 24939
rect 16980 24919 16982 24939
rect 17148 24919 17150 24939
rect 17196 24919 17198 24939
rect 17220 24919 17222 24939
rect 17292 24919 17294 24939
rect 17316 24919 17318 24939
rect 18132 24919 18134 24939
rect 18228 24919 18230 24939
rect 18492 24919 18494 24939
rect 18516 24919 18518 24939
rect 18612 24919 18614 24939
rect 18636 24919 18638 24939
rect 18711 24936 18725 24939
rect 18732 24939 23675 24943
rect 18732 24936 18749 24939
rect 18732 24919 18734 24936
rect 18828 24919 18830 24939
rect 18900 24919 18902 24939
rect 18924 24919 18926 24939
rect 18961 24934 18964 24939
rect 18985 24934 18988 24939
rect 18996 24934 18998 24939
rect 18971 24920 18974 24934
rect 18995 24920 18998 24934
rect 18972 24919 18974 24920
rect 19020 24919 19022 24939
rect 19092 24936 19094 24939
rect 19092 24919 19095 24936
rect 19140 24919 19142 24939
rect 19236 24919 19238 24939
rect 19260 24919 19262 24939
rect 19788 24919 19790 24939
rect 19836 24919 19838 24939
rect 19860 24919 19862 24939
rect 19884 24919 19886 24939
rect 19956 24919 19958 24939
rect 19980 24919 19982 24939
rect 20052 24919 20054 24939
rect 20076 24919 20078 24939
rect 20124 24919 20126 24939
rect 20172 24919 20174 24939
rect 20196 24919 20198 24939
rect 20292 24919 20294 24939
rect 20388 24919 20390 24939
rect 20412 24919 20414 24939
rect 20508 24919 20510 24939
rect 20532 24919 20534 24939
rect 20604 24919 20606 24939
rect 20628 24919 20630 24939
rect 20892 24919 20894 24939
rect 20964 24919 20966 24939
rect 20988 24919 20990 24939
rect 21108 24919 21110 24939
rect 21204 24919 21206 24939
rect 21300 24919 21302 24939
rect 21324 24919 21326 24939
rect 21444 24919 21446 24939
rect 21468 24919 21470 24939
rect 21564 24919 21566 24939
rect 21588 24919 21590 24939
rect 21684 24919 21686 24939
rect 21708 24919 21710 24939
rect 21828 24919 21830 24939
rect 21924 24919 21926 24939
rect 22068 24919 22070 24939
rect 22188 24919 22190 24939
rect 22212 24919 22214 24939
rect 22884 24919 22886 24939
rect 22980 24919 22982 24939
rect 23076 24919 23078 24939
rect 23100 24919 23102 24939
rect 23124 24919 23126 24939
rect 23244 24919 23246 24939
rect 23340 24919 23342 24939
rect 23412 24919 23414 24939
rect 23460 24920 23462 24939
rect 23508 24920 23510 24939
rect 23556 24920 23558 24939
rect 23593 24934 23596 24939
rect 23604 24934 23606 24939
rect 23641 24934 23644 24939
rect 23652 24934 23654 24939
rect 23603 24920 23606 24934
rect 23651 24920 23654 24934
rect 23665 24926 23669 24934
rect 23655 24920 23665 24926
rect 23449 24919 23483 24920
rect -12431 24915 -8539 24919
rect -12431 24912 -12427 24915
rect -12420 24912 -12417 24915
rect -12311 24895 -12277 24896
rect -12239 24895 -12205 24896
rect -12311 24891 -12205 24895
rect -12191 24895 -12157 24896
rect -12084 24895 -12082 24915
rect -11817 24912 -11803 24915
rect -11975 24895 -11917 24896
rect -11772 24895 -11770 24915
rect -11676 24895 -11674 24915
rect -11663 24910 -11660 24915
rect -11652 24910 -11650 24915
rect -11653 24896 -11650 24910
rect -11508 24895 -11506 24915
rect -11436 24895 -11434 24915
rect -11412 24895 -11410 24915
rect -11196 24895 -11194 24915
rect -11100 24895 -11098 24915
rect -10689 24912 -10675 24915
rect -10569 24912 -10555 24915
rect -9900 24895 -9898 24915
rect -9732 24895 -9730 24915
rect -9636 24895 -9634 24915
rect -9540 24895 -9538 24915
rect -9444 24895 -9442 24915
rect -9348 24895 -9346 24915
rect -9228 24895 -9226 24915
rect -9108 24895 -9106 24915
rect -9023 24910 -9020 24915
rect -9013 24896 -9010 24910
rect -9012 24895 -9010 24896
rect -8916 24895 -8913 24912
rect -8628 24895 -8626 24915
rect -8553 24912 -8539 24915
rect -8532 24915 13085 24919
rect -8532 24912 -8515 24915
rect -8532 24895 -8530 24912
rect -8436 24895 -8434 24915
rect -8364 24895 -8362 24915
rect -8340 24895 -8338 24915
rect -8268 24895 -8266 24915
rect -8159 24895 -8125 24896
rect -8124 24895 -8122 24915
rect -7764 24895 -7762 24915
rect -7524 24895 -7522 24915
rect -7356 24895 -7354 24915
rect -7308 24895 -7306 24915
rect -7140 24895 -7138 24915
rect -7044 24895 -7042 24915
rect -6948 24895 -6946 24915
rect -6852 24895 -6850 24915
rect -6732 24895 -6730 24915
rect -6516 24895 -6514 24915
rect -5892 24895 -5890 24915
rect -5436 24895 -5434 24915
rect -5340 24895 -5338 24915
rect -5289 24912 -5275 24915
rect -5196 24895 -5194 24915
rect -4716 24895 -4714 24915
rect -4500 24895 -4498 24915
rect -4404 24895 -4402 24915
rect -4308 24895 -4306 24915
rect -4164 24895 -4162 24915
rect -3876 24895 -3874 24915
rect -3743 24910 -3740 24915
rect -3732 24910 -3730 24915
rect -3733 24896 -3730 24910
rect -3636 24912 -3634 24915
rect -3636 24895 -3633 24912
rect -3540 24895 -3538 24915
rect -3468 24895 -3466 24915
rect -3324 24895 -3322 24915
rect -3108 24895 -3106 24915
rect -3012 24895 -3010 24915
rect -2964 24895 -2962 24915
rect -2916 24895 -2914 24915
rect -2868 24895 -2866 24915
rect -2820 24895 -2818 24915
rect -2817 24912 -2803 24915
rect -2772 24895 -2770 24915
rect -2676 24895 -2674 24915
rect -2364 24895 -2362 24915
rect -2316 24895 -2314 24915
rect -2076 24895 -2074 24915
rect -1980 24895 -1978 24915
rect -1812 24895 -1810 24915
rect -1572 24895 -1570 24915
rect -1476 24895 -1474 24915
rect -1356 24895 -1354 24915
rect -1260 24895 -1258 24915
rect -1236 24895 -1234 24915
rect -1140 24895 -1138 24915
rect -876 24895 -874 24915
rect -660 24895 -658 24915
rect -492 24895 -490 24915
rect -396 24895 -394 24915
rect -372 24895 -370 24915
rect -276 24895 -274 24915
rect -12 24895 -10 24915
rect 73 24910 76 24915
rect 83 24896 86 24910
rect 84 24895 86 24896
rect 156 24895 158 24915
rect 204 24912 206 24915
rect 204 24895 207 24912
rect 252 24895 254 24915
rect 348 24895 350 24915
rect 468 24895 470 24915
rect 492 24895 494 24915
rect 564 24895 566 24915
rect 588 24895 590 24915
rect 636 24895 638 24915
rect 660 24895 662 24915
rect 732 24895 734 24915
rect 937 24895 995 24896
rect 1092 24895 1094 24915
rect 1140 24895 1142 24915
rect 1308 24895 1310 24915
rect 1356 24895 1358 24915
rect 1428 24895 1430 24915
rect 1692 24895 1694 24915
rect 1860 24895 1862 24915
rect 2076 24895 2078 24915
rect 2100 24895 2102 24915
rect 2244 24895 2246 24915
rect 2460 24895 2462 24915
rect 2772 24895 2774 24915
rect 2868 24895 2870 24915
rect 2940 24895 2942 24915
rect 3012 24895 3014 24915
rect 3108 24895 3110 24915
rect 3324 24895 3326 24915
rect 3396 24895 3398 24915
rect 3564 24895 3566 24915
rect 3660 24895 3662 24915
rect 3780 24895 3782 24915
rect 4092 24895 4094 24915
rect 4188 24895 4190 24915
rect 4308 24895 4310 24915
rect 4404 24895 4406 24915
rect 4500 24895 4502 24915
rect 4596 24895 4598 24915
rect 4692 24895 4694 24915
rect 4956 24895 4958 24915
rect 4980 24895 4982 24915
rect 5052 24895 5054 24915
rect 5124 24895 5126 24915
rect 5220 24895 5222 24915
rect 5268 24895 5270 24915
rect 5388 24895 5390 24915
rect 5484 24895 5486 24915
rect 5508 24895 5510 24915
rect 5532 24895 5534 24915
rect 5628 24895 5630 24915
rect 5652 24895 5654 24915
rect 5748 24895 5750 24915
rect 5796 24895 5798 24915
rect 5844 24895 5846 24915
rect 5892 24895 5894 24915
rect 6217 24910 6220 24915
rect 6228 24910 6230 24915
rect 6227 24896 6230 24910
rect 6276 24895 6278 24915
rect 6324 24912 6326 24915
rect 6327 24912 6341 24915
rect 6324 24895 6327 24912
rect 6372 24895 6374 24915
rect 6420 24895 6422 24915
rect 6492 24895 6494 24915
rect 6516 24895 6518 24915
rect 6588 24895 6590 24915
rect 6612 24895 6614 24915
rect 6684 24895 6686 24915
rect 6708 24895 6710 24915
rect 6780 24895 6782 24915
rect 6804 24895 6806 24915
rect 6900 24895 6902 24915
rect 6924 24895 6926 24915
rect 7020 24895 7022 24915
rect 7164 24895 7166 24915
rect 7236 24895 7238 24915
rect 7308 24895 7310 24915
rect 7380 24895 7382 24915
rect 7404 24895 7406 24915
rect 7476 24895 7478 24915
rect 7489 24895 7547 24896
rect 7572 24895 7574 24915
rect 7620 24895 7622 24915
rect 7644 24895 7646 24915
rect 7668 24895 7670 24915
rect 7908 24895 7910 24915
rect 8124 24895 8126 24915
rect 8220 24895 8222 24915
rect 8652 24895 8654 24915
rect 8700 24895 8702 24915
rect 8748 24895 8750 24915
rect 8796 24895 8798 24915
rect 8844 24895 8846 24915
rect 8868 24895 8870 24915
rect 9516 24895 9518 24915
rect 9660 24895 9662 24915
rect 9684 24895 9686 24915
rect 9756 24895 9758 24915
rect 9780 24895 9782 24915
rect 9804 24895 9806 24915
rect 9852 24895 9854 24915
rect 9948 24895 9950 24915
rect 10044 24895 10046 24915
rect 10116 24895 10118 24915
rect 10140 24895 10142 24915
rect 10188 24895 10190 24915
rect 10236 24895 10238 24915
rect 10284 24895 10286 24915
rect 10332 24895 10334 24915
rect 10380 24895 10382 24915
rect 10428 24895 10430 24915
rect 10476 24895 10478 24915
rect 10524 24895 10526 24915
rect 10620 24895 10622 24915
rect 10644 24895 10646 24915
rect 10716 24895 10718 24915
rect 10873 24910 10876 24915
rect 10883 24896 10886 24910
rect 10884 24895 10886 24896
rect 10956 24895 10958 24915
rect 11004 24912 11006 24915
rect 11004 24895 11007 24912
rect 11052 24895 11054 24915
rect 11100 24895 11102 24915
rect 11172 24895 11174 24915
rect 11220 24895 11222 24915
rect 11340 24895 11342 24915
rect 11436 24895 11438 24915
rect 11532 24895 11534 24915
rect 11628 24895 11630 24915
rect 11676 24895 11678 24915
rect 11724 24895 11726 24915
rect 11772 24895 11774 24915
rect 11796 24895 11798 24915
rect 11892 24895 11894 24915
rect 11988 24895 11990 24915
rect 12060 24895 12062 24915
rect 12276 24895 12278 24915
rect 12324 24895 12326 24915
rect 12372 24895 12374 24915
rect 12420 24895 12422 24915
rect 12444 24895 12446 24915
rect 12468 24895 12470 24915
rect 12516 24895 12518 24915
rect 12540 24895 12542 24915
rect 12564 24895 12566 24915
rect 12660 24895 12662 24915
rect 12756 24895 12758 24915
rect 12828 24895 12830 24915
rect 12876 24895 12878 24915
rect 12972 24895 12974 24915
rect 13044 24895 13046 24915
rect 13068 24895 13070 24915
rect 13071 24912 13085 24915
rect 13095 24915 19061 24919
rect 13095 24912 13109 24915
rect 13116 24912 13119 24915
rect 13284 24895 13286 24915
rect 13332 24895 13334 24915
rect 13500 24895 13502 24915
rect 13572 24895 13574 24915
rect 13668 24895 13670 24915
rect 13716 24895 13718 24915
rect 13764 24895 13766 24915
rect 13860 24895 13862 24915
rect 13956 24895 13958 24915
rect 14004 24895 14006 24915
rect 14100 24895 14102 24915
rect 14940 24895 14942 24915
rect 15036 24895 15038 24915
rect 15049 24895 15107 24896
rect 15180 24895 15182 24915
rect 15276 24895 15278 24915
rect 15420 24895 15422 24915
rect 15492 24895 15494 24915
rect 15660 24895 15662 24915
rect 15708 24895 15710 24915
rect 15732 24895 15734 24915
rect 15756 24895 15758 24915
rect 15804 24895 15806 24915
rect 15828 24895 15830 24915
rect 15852 24895 15854 24915
rect 15948 24895 15950 24915
rect 15972 24895 15974 24915
rect 16044 24895 16046 24915
rect 16068 24895 16070 24915
rect 16164 24895 16166 24915
rect 16260 24895 16262 24915
rect 16332 24895 16334 24915
rect 16369 24910 16372 24915
rect 16379 24896 16382 24910
rect 16380 24895 16382 24896
rect 16476 24895 16479 24912
rect 16548 24895 16550 24915
rect 16572 24895 16574 24915
rect 16620 24895 16622 24915
rect 16668 24895 16670 24915
rect 16716 24895 16718 24915
rect 16764 24895 16766 24915
rect 16812 24895 16814 24915
rect 16884 24895 16886 24915
rect 16908 24895 16910 24915
rect 16980 24895 16982 24915
rect 17148 24895 17150 24915
rect 17196 24895 17198 24915
rect 17220 24895 17222 24915
rect 17292 24895 17294 24915
rect 17316 24895 17318 24915
rect 18132 24895 18134 24915
rect 18228 24895 18230 24915
rect 18409 24895 18443 24896
rect 18492 24895 18494 24915
rect 18516 24896 18518 24915
rect 18505 24895 18539 24896
rect 18612 24895 18614 24915
rect 18636 24895 18638 24915
rect 18732 24895 18734 24915
rect 18793 24895 18827 24896
rect 18828 24895 18830 24915
rect 18900 24895 18902 24915
rect 18924 24895 18926 24915
rect 18972 24895 18974 24915
rect 19020 24895 19022 24915
rect 19047 24912 19061 24915
rect 19071 24915 23483 24919
rect 23497 24919 23531 24920
rect 23545 24919 23579 24920
rect 23497 24915 23579 24919
rect 19071 24912 19085 24915
rect 19092 24912 19095 24915
rect 19057 24895 19115 24896
rect 19140 24895 19142 24915
rect 19236 24895 19238 24915
rect 19260 24895 19262 24915
rect 19788 24895 19790 24915
rect 19836 24895 19838 24915
rect 19860 24895 19862 24915
rect 19884 24895 19886 24915
rect 19956 24895 19958 24915
rect 19980 24895 19982 24915
rect 20052 24895 20054 24915
rect 20076 24895 20078 24915
rect 20124 24895 20126 24915
rect 20172 24895 20174 24915
rect 20196 24895 20198 24915
rect 20292 24895 20294 24915
rect 20388 24895 20390 24915
rect 20412 24895 20414 24915
rect 20508 24895 20510 24915
rect 20532 24895 20534 24915
rect 20604 24895 20606 24915
rect 20628 24895 20630 24915
rect 20737 24895 20771 24896
rect 20892 24895 20894 24915
rect 20964 24895 20966 24915
rect 20988 24895 20990 24915
rect 21108 24895 21110 24915
rect 21204 24895 21206 24915
rect 21300 24895 21302 24915
rect 21324 24895 21326 24915
rect 21444 24895 21446 24915
rect 21468 24895 21470 24915
rect 21564 24895 21566 24915
rect 21588 24895 21590 24915
rect 21684 24895 21686 24915
rect 21708 24895 21710 24915
rect 21828 24895 21830 24915
rect 21924 24895 21926 24915
rect 22068 24895 22070 24915
rect 22188 24895 22190 24915
rect 22212 24895 22214 24915
rect 22884 24895 22886 24915
rect 22980 24895 22982 24915
rect 23076 24895 23078 24915
rect 23100 24895 23102 24915
rect 23124 24895 23126 24915
rect 23244 24895 23246 24915
rect 23340 24896 23342 24915
rect 23412 24896 23414 24915
rect 23449 24910 23452 24915
rect 23460 24910 23462 24915
rect 23497 24910 23500 24915
rect 23508 24910 23510 24915
rect 23545 24910 23548 24915
rect 23556 24912 23558 24915
rect 23556 24910 23559 24912
rect 23459 24896 23462 24910
rect 23507 24896 23510 24910
rect 23555 24896 23559 24910
rect 23329 24895 23387 24896
rect 23401 24895 23435 24896
rect -12191 24891 -8923 24895
rect -12084 24888 -12082 24891
rect -12215 24878 -12211 24886
rect -12225 24872 -12215 24878
rect -12084 24872 -12081 24888
rect -12095 24871 -12061 24872
rect -11868 24871 -11865 24888
rect -11772 24871 -11770 24891
rect -11676 24871 -11674 24891
rect -11577 24888 -11563 24891
rect -11508 24871 -11506 24891
rect -11436 24871 -11434 24891
rect -11412 24871 -11410 24891
rect -11196 24871 -11194 24891
rect -11100 24871 -11098 24891
rect -9900 24871 -9898 24891
rect -9732 24871 -9730 24891
rect -9636 24871 -9634 24891
rect -9540 24871 -9538 24891
rect -9444 24871 -9442 24891
rect -9348 24871 -9346 24891
rect -9228 24871 -9226 24891
rect -9108 24871 -9106 24891
rect -9012 24871 -9010 24891
rect -8937 24888 -8923 24891
rect -8916 24891 -3667 24895
rect -8916 24888 -8899 24891
rect -8916 24871 -8914 24888
rect -8628 24871 -8626 24891
rect -8532 24871 -8530 24891
rect -8436 24871 -8434 24891
rect -8364 24871 -8362 24891
rect -8340 24871 -8338 24891
rect -8268 24871 -8266 24891
rect -8124 24871 -8122 24891
rect -7764 24871 -7762 24891
rect -7524 24871 -7522 24891
rect -7356 24871 -7354 24891
rect -7308 24871 -7306 24891
rect -7140 24871 -7138 24891
rect -7044 24871 -7042 24891
rect -6948 24871 -6946 24891
rect -6852 24871 -6850 24891
rect -6732 24871 -6730 24891
rect -6516 24871 -6514 24891
rect -5892 24871 -5890 24891
rect -5436 24871 -5434 24891
rect -5340 24871 -5338 24891
rect -5196 24871 -5194 24891
rect -4716 24871 -4714 24891
rect -4500 24871 -4498 24891
rect -4404 24871 -4402 24891
rect -4308 24871 -4306 24891
rect -4164 24871 -4162 24891
rect -3876 24871 -3874 24891
rect -3681 24888 -3667 24891
rect -3657 24891 173 24895
rect -3657 24888 -3643 24891
rect -3636 24888 -3633 24891
rect -3540 24871 -3538 24891
rect -3468 24871 -3466 24891
rect -3324 24871 -3322 24891
rect -3108 24871 -3106 24891
rect -3012 24871 -3010 24891
rect -2964 24871 -2962 24891
rect -2916 24871 -2914 24891
rect -2868 24871 -2866 24891
rect -2820 24871 -2818 24891
rect -2772 24871 -2770 24891
rect -2676 24871 -2674 24891
rect -2364 24871 -2362 24891
rect -2316 24871 -2314 24891
rect -2076 24871 -2074 24891
rect -1980 24871 -1978 24891
rect -1812 24871 -1810 24891
rect -1572 24871 -1570 24891
rect -1476 24871 -1474 24891
rect -1356 24871 -1354 24891
rect -1260 24871 -1258 24891
rect -1236 24871 -1234 24891
rect -1140 24871 -1138 24891
rect -876 24871 -874 24891
rect -660 24871 -658 24891
rect -492 24871 -490 24891
rect -396 24871 -394 24891
rect -372 24871 -370 24891
rect -276 24871 -274 24891
rect -12 24871 -10 24891
rect 84 24871 86 24891
rect 156 24871 158 24891
rect 159 24888 173 24891
rect 183 24891 6293 24895
rect 183 24888 197 24891
rect 204 24888 207 24891
rect 252 24871 254 24891
rect 348 24871 350 24891
rect 468 24871 470 24891
rect 492 24871 494 24891
rect 564 24871 566 24891
rect 588 24871 590 24891
rect 636 24871 638 24891
rect 660 24871 662 24891
rect 732 24871 734 24891
rect 937 24886 940 24891
rect 947 24872 950 24886
rect 948 24871 950 24872
rect 1044 24871 1047 24888
rect 1092 24871 1094 24891
rect 1140 24871 1142 24891
rect 1308 24871 1310 24891
rect 1356 24871 1358 24891
rect 1428 24871 1430 24891
rect 1692 24871 1694 24891
rect 1860 24871 1862 24891
rect 2076 24871 2078 24891
rect 2100 24871 2102 24891
rect 2244 24871 2246 24891
rect 2460 24871 2462 24891
rect 2772 24871 2774 24891
rect 2868 24871 2870 24891
rect 2940 24871 2942 24891
rect 3012 24871 3014 24891
rect 3108 24871 3110 24891
rect 3324 24871 3326 24891
rect 3396 24871 3398 24891
rect 3564 24871 3566 24891
rect 3660 24871 3662 24891
rect 3780 24871 3782 24891
rect 4092 24871 4094 24891
rect 4188 24871 4190 24891
rect 4308 24871 4310 24891
rect 4404 24871 4406 24891
rect 4500 24871 4502 24891
rect 4596 24871 4598 24891
rect 4692 24871 4694 24891
rect 4956 24871 4958 24891
rect 4980 24871 4982 24891
rect 5052 24871 5054 24891
rect 5124 24871 5126 24891
rect 5220 24871 5222 24891
rect 5268 24871 5270 24891
rect 5388 24871 5390 24891
rect 5484 24871 5486 24891
rect 5508 24871 5510 24891
rect 5532 24871 5534 24891
rect 5628 24871 5630 24891
rect 5652 24871 5654 24891
rect 5748 24871 5750 24891
rect 5796 24871 5798 24891
rect 5844 24871 5846 24891
rect 5892 24871 5894 24891
rect 6276 24871 6278 24891
rect 6279 24888 6293 24891
rect 6303 24891 10973 24895
rect 6303 24888 6317 24891
rect 6324 24888 6327 24891
rect 6372 24871 6374 24891
rect 6420 24871 6422 24891
rect 6492 24871 6494 24891
rect 6516 24871 6518 24891
rect 6588 24871 6590 24891
rect 6612 24871 6614 24891
rect 6684 24871 6686 24891
rect 6708 24871 6710 24891
rect 6780 24871 6782 24891
rect 6804 24871 6806 24891
rect 6900 24871 6902 24891
rect 6924 24871 6926 24891
rect 7020 24871 7022 24891
rect 7164 24871 7166 24891
rect 7236 24871 7238 24891
rect 7308 24871 7310 24891
rect 7380 24871 7382 24891
rect 7404 24871 7406 24891
rect 7476 24871 7478 24891
rect 7489 24886 7492 24891
rect 7499 24872 7502 24886
rect 7500 24871 7502 24872
rect 7572 24871 7574 24891
rect 7620 24888 7622 24891
rect 7620 24871 7623 24888
rect 7644 24871 7646 24891
rect 7668 24871 7670 24891
rect 7908 24871 7910 24891
rect 8124 24871 8126 24891
rect 8220 24871 8222 24891
rect 8652 24871 8654 24891
rect 8700 24871 8702 24891
rect 8748 24871 8750 24891
rect 8796 24871 8798 24891
rect 8844 24871 8846 24891
rect 8868 24871 8870 24891
rect 9516 24871 9518 24891
rect 9660 24871 9662 24891
rect 9684 24871 9686 24891
rect 9756 24871 9758 24891
rect 9780 24871 9782 24891
rect 9804 24871 9806 24891
rect 9852 24871 9854 24891
rect 9948 24871 9950 24891
rect 10044 24871 10046 24891
rect 10116 24871 10118 24891
rect 10140 24871 10142 24891
rect 10188 24871 10190 24891
rect 10236 24871 10238 24891
rect 10284 24871 10286 24891
rect 10332 24871 10334 24891
rect 10380 24871 10382 24891
rect 10428 24871 10430 24891
rect 10476 24871 10478 24891
rect 10524 24871 10526 24891
rect 10620 24871 10622 24891
rect 10644 24871 10646 24891
rect 10716 24871 10718 24891
rect 10884 24871 10886 24891
rect 10956 24871 10958 24891
rect 10959 24888 10973 24891
rect 10983 24891 16469 24895
rect 10983 24888 10997 24891
rect 11004 24888 11007 24891
rect 11052 24871 11054 24891
rect 11100 24871 11102 24891
rect 11172 24871 11174 24891
rect 11220 24871 11222 24891
rect 11340 24871 11342 24891
rect 11436 24871 11438 24891
rect 11532 24871 11534 24891
rect 11628 24871 11630 24891
rect 11676 24871 11678 24891
rect 11724 24871 11726 24891
rect 11772 24871 11774 24891
rect 11796 24871 11798 24891
rect 11892 24871 11894 24891
rect 11988 24871 11990 24891
rect 12060 24871 12062 24891
rect 12276 24871 12278 24891
rect 12324 24871 12326 24891
rect 12372 24871 12374 24891
rect 12420 24871 12422 24891
rect 12444 24871 12446 24891
rect 12468 24871 12470 24891
rect 12516 24871 12518 24891
rect 12540 24871 12542 24891
rect 12564 24871 12566 24891
rect 12660 24871 12662 24891
rect 12756 24871 12758 24891
rect 12828 24871 12830 24891
rect 12876 24871 12878 24891
rect 12972 24871 12974 24891
rect 13044 24871 13046 24891
rect 13068 24871 13070 24891
rect 13284 24871 13286 24891
rect 13332 24871 13334 24891
rect 13500 24871 13502 24891
rect 13572 24871 13574 24891
rect 13668 24871 13670 24891
rect 13716 24871 13718 24891
rect 13764 24871 13766 24891
rect 13860 24871 13862 24891
rect 13956 24871 13958 24891
rect 14004 24871 14006 24891
rect 14100 24871 14102 24891
rect 14940 24871 14942 24891
rect 15036 24871 15038 24891
rect 15180 24888 15182 24891
rect 15180 24871 15183 24888
rect 15276 24871 15278 24891
rect 15420 24871 15422 24891
rect 15492 24871 15494 24891
rect 15660 24871 15662 24891
rect 15708 24871 15710 24891
rect 15732 24871 15734 24891
rect 15756 24871 15758 24891
rect 15804 24871 15806 24891
rect 15828 24871 15830 24891
rect 15852 24871 15854 24891
rect 15948 24871 15950 24891
rect 15972 24871 15974 24891
rect 16044 24871 16046 24891
rect 16068 24871 16070 24891
rect 16164 24871 16166 24891
rect 16260 24871 16262 24891
rect 16332 24871 16334 24891
rect 16380 24871 16382 24891
rect 16455 24888 16469 24891
rect 16476 24891 23435 24895
rect 16476 24888 16493 24891
rect 16476 24871 16478 24888
rect 16548 24871 16550 24891
rect 16572 24871 16574 24891
rect 16620 24871 16622 24891
rect 16668 24871 16670 24891
rect 16716 24871 16718 24891
rect 16764 24871 16766 24891
rect 16812 24871 16814 24891
rect 16884 24871 16886 24891
rect 16908 24871 16910 24891
rect 16980 24871 16982 24891
rect 17148 24871 17150 24891
rect 17196 24871 17198 24891
rect 17220 24871 17222 24891
rect 17292 24871 17294 24891
rect 17316 24871 17318 24891
rect 18132 24871 18134 24891
rect 18228 24871 18230 24891
rect 18492 24871 18494 24891
rect 18505 24886 18508 24891
rect 18516 24888 18518 24891
rect 18612 24888 18614 24891
rect 18516 24886 18519 24888
rect 18515 24872 18519 24886
rect 18612 24871 18615 24888
rect 18636 24871 18638 24891
rect 18732 24871 18734 24891
rect 18828 24871 18830 24891
rect 18900 24888 18902 24891
rect 18900 24871 18903 24888
rect 18924 24871 18926 24891
rect 18972 24871 18974 24891
rect 19020 24871 19022 24891
rect 19057 24886 19060 24891
rect 19067 24872 19070 24886
rect 19068 24871 19070 24872
rect 19140 24871 19142 24891
rect 19164 24871 19167 24888
rect 19236 24871 19238 24891
rect 19260 24871 19262 24891
rect 19788 24871 19790 24891
rect 19836 24871 19838 24891
rect 19860 24871 19862 24891
rect 19884 24871 19886 24891
rect 19956 24871 19958 24891
rect 19980 24871 19982 24891
rect 19993 24871 20051 24872
rect 20052 24871 20054 24891
rect 20076 24871 20078 24891
rect 20124 24871 20126 24891
rect 20172 24871 20174 24891
rect 20196 24871 20198 24891
rect 20292 24871 20294 24891
rect 20388 24871 20390 24891
rect 20412 24871 20414 24891
rect 20508 24871 20510 24891
rect 20532 24871 20534 24891
rect 20604 24871 20606 24891
rect 20628 24871 20630 24891
rect 20892 24871 20894 24891
rect 20964 24871 20966 24891
rect 20988 24871 20990 24891
rect 21108 24871 21110 24891
rect 21204 24871 21206 24891
rect 21300 24871 21302 24891
rect 21324 24871 21326 24891
rect 21444 24871 21446 24891
rect 21468 24871 21470 24891
rect 21564 24871 21566 24891
rect 21588 24871 21590 24891
rect 21684 24871 21686 24891
rect 21708 24871 21710 24891
rect 21828 24871 21830 24891
rect 21924 24871 21926 24891
rect 22068 24871 22070 24891
rect 22188 24871 22190 24891
rect 22212 24871 22214 24891
rect 22884 24871 22886 24891
rect 22980 24871 22982 24891
rect 23076 24871 23078 24891
rect 23100 24871 23102 24891
rect 23124 24871 23126 24891
rect 23244 24871 23246 24891
rect 23329 24886 23332 24891
rect 23340 24886 23342 24891
rect 23401 24886 23404 24891
rect 23412 24886 23414 24891
rect 23339 24872 23342 24886
rect 23411 24872 23414 24886
rect 23425 24878 23429 24886
rect 23415 24872 23425 24878
rect 23305 24871 23339 24872
rect -12095 24867 -11875 24871
rect -12095 24864 -12091 24867
rect -12084 24864 -12081 24867
rect -11889 24864 -11875 24867
rect -11868 24867 1037 24871
rect -11868 24864 -11851 24867
rect -11975 24847 -11941 24848
rect -11868 24847 -11866 24864
rect -11772 24847 -11770 24867
rect -11676 24847 -11674 24867
rect -11508 24847 -11506 24867
rect -11436 24847 -11434 24867
rect -11412 24847 -11410 24867
rect -11196 24847 -11194 24867
rect -11100 24847 -11098 24867
rect -9900 24847 -9898 24867
rect -9732 24847 -9730 24867
rect -9636 24847 -9634 24867
rect -9540 24847 -9538 24867
rect -9444 24847 -9442 24867
rect -9348 24847 -9346 24867
rect -9228 24847 -9226 24867
rect -9108 24847 -9106 24867
rect -9012 24847 -9010 24867
rect -8916 24847 -8914 24867
rect -8628 24847 -8626 24867
rect -8532 24847 -8530 24867
rect -8436 24847 -8434 24867
rect -8364 24847 -8362 24867
rect -8340 24847 -8338 24867
rect -8268 24847 -8266 24867
rect -8124 24847 -8122 24867
rect -8073 24864 -8059 24867
rect -7764 24847 -7762 24867
rect -7524 24847 -7522 24867
rect -7356 24847 -7354 24867
rect -7308 24847 -7306 24867
rect -7140 24847 -7138 24867
rect -7044 24847 -7042 24867
rect -6948 24847 -6946 24867
rect -6852 24847 -6850 24867
rect -6732 24847 -6730 24867
rect -6516 24847 -6514 24867
rect -5892 24847 -5890 24867
rect -5436 24847 -5434 24867
rect -5340 24847 -5338 24867
rect -5196 24847 -5194 24867
rect -4716 24847 -4714 24867
rect -4500 24847 -4498 24867
rect -4404 24847 -4402 24867
rect -4308 24847 -4306 24867
rect -4164 24847 -4162 24867
rect -3876 24847 -3874 24867
rect -3540 24847 -3538 24867
rect -3468 24847 -3466 24867
rect -3324 24847 -3322 24867
rect -3108 24847 -3106 24867
rect -3012 24847 -3010 24867
rect -2964 24847 -2962 24867
rect -2916 24847 -2914 24867
rect -2868 24847 -2866 24867
rect -2820 24847 -2818 24867
rect -2772 24847 -2770 24867
rect -2676 24847 -2674 24867
rect -2364 24847 -2362 24867
rect -2316 24847 -2314 24867
rect -2076 24847 -2074 24867
rect -1980 24847 -1978 24867
rect -1812 24847 -1810 24867
rect -1572 24847 -1570 24867
rect -1476 24847 -1474 24867
rect -1356 24847 -1354 24867
rect -1260 24847 -1258 24867
rect -1236 24847 -1234 24867
rect -1140 24847 -1138 24867
rect -876 24847 -874 24867
rect -660 24847 -658 24867
rect -492 24847 -490 24867
rect -396 24847 -394 24867
rect -372 24847 -370 24867
rect -276 24847 -274 24867
rect -12 24847 -10 24867
rect 84 24847 86 24867
rect 156 24847 158 24867
rect 252 24847 254 24867
rect 348 24847 350 24867
rect 468 24847 470 24867
rect 492 24847 494 24867
rect 564 24847 566 24867
rect 588 24847 590 24867
rect 636 24847 638 24867
rect 660 24847 662 24867
rect 732 24847 734 24867
rect 948 24847 950 24867
rect 1023 24864 1037 24867
rect 1044 24867 7589 24871
rect 1044 24864 1061 24867
rect 1044 24847 1046 24864
rect 1092 24847 1094 24867
rect 1140 24847 1142 24867
rect 1308 24847 1310 24867
rect 1356 24847 1358 24867
rect 1428 24847 1430 24867
rect 1692 24847 1694 24867
rect 1860 24847 1862 24867
rect 2076 24847 2078 24867
rect 2100 24847 2102 24867
rect 2244 24847 2246 24867
rect 2460 24847 2462 24867
rect 2772 24847 2774 24867
rect 2868 24847 2870 24867
rect 2940 24847 2942 24867
rect 3012 24847 3014 24867
rect 3108 24847 3110 24867
rect 3324 24847 3326 24867
rect 3396 24847 3398 24867
rect 3564 24847 3566 24867
rect 3660 24847 3662 24867
rect 3780 24847 3782 24867
rect 4092 24847 4094 24867
rect 4188 24847 4190 24867
rect 4308 24847 4310 24867
rect 4404 24847 4406 24867
rect 4500 24847 4502 24867
rect 4596 24847 4598 24867
rect 4692 24847 4694 24867
rect 4956 24847 4958 24867
rect 4980 24847 4982 24867
rect 5052 24847 5054 24867
rect 5124 24847 5126 24867
rect 5220 24847 5222 24867
rect 5268 24848 5270 24867
rect 5233 24847 5291 24848
rect 5388 24847 5390 24867
rect 5484 24847 5486 24867
rect 5508 24847 5510 24867
rect 5532 24847 5534 24867
rect 5628 24847 5630 24867
rect 5652 24847 5654 24867
rect 5748 24847 5750 24867
rect 5796 24847 5798 24867
rect 5844 24847 5846 24867
rect 5892 24847 5894 24867
rect 6276 24847 6278 24867
rect 6372 24847 6374 24867
rect 6420 24847 6422 24867
rect 6492 24847 6494 24867
rect 6516 24847 6518 24867
rect 6588 24847 6590 24867
rect 6612 24847 6614 24867
rect 6684 24847 6686 24867
rect 6708 24847 6710 24867
rect 6780 24847 6782 24867
rect 6804 24847 6806 24867
rect 6900 24847 6902 24867
rect 6924 24847 6926 24867
rect 7020 24847 7022 24867
rect 7164 24847 7166 24867
rect 7236 24847 7238 24867
rect 7308 24847 7310 24867
rect 7380 24847 7382 24867
rect 7404 24847 7406 24867
rect 7476 24847 7478 24867
rect 7500 24847 7502 24867
rect 7572 24847 7574 24867
rect 7575 24864 7589 24867
rect 7599 24867 15149 24871
rect 7599 24864 7613 24867
rect 7620 24864 7623 24867
rect 7644 24847 7646 24867
rect 7668 24847 7670 24867
rect 7908 24847 7910 24867
rect 8124 24847 8126 24867
rect 8220 24847 8222 24867
rect 8652 24847 8654 24867
rect 8700 24847 8702 24867
rect 8748 24847 8750 24867
rect 8796 24847 8798 24867
rect 8844 24847 8846 24867
rect 8868 24847 8870 24867
rect 9516 24847 9518 24867
rect 9660 24847 9662 24867
rect 9684 24847 9686 24867
rect 9756 24847 9758 24867
rect 9780 24847 9782 24867
rect 9804 24847 9806 24867
rect 9852 24847 9854 24867
rect 9948 24847 9950 24867
rect 10044 24847 10046 24867
rect 10116 24847 10118 24867
rect 10140 24847 10142 24867
rect 10188 24847 10190 24867
rect 10236 24847 10238 24867
rect 10284 24847 10286 24867
rect 10332 24847 10334 24867
rect 10380 24847 10382 24867
rect 10428 24847 10430 24867
rect 10476 24847 10478 24867
rect 10524 24847 10526 24867
rect 10620 24847 10622 24867
rect 10644 24847 10646 24867
rect 10716 24847 10718 24867
rect 10884 24847 10886 24867
rect 10956 24847 10958 24867
rect 11052 24847 11054 24867
rect 11100 24847 11102 24867
rect 11172 24847 11174 24867
rect 11220 24847 11222 24867
rect 11340 24847 11342 24867
rect 11436 24847 11438 24867
rect 11532 24847 11534 24867
rect 11628 24847 11630 24867
rect 11676 24847 11678 24867
rect 11724 24847 11726 24867
rect 11772 24847 11774 24867
rect 11796 24847 11798 24867
rect 11892 24847 11894 24867
rect 11988 24847 11990 24867
rect 12060 24847 12062 24867
rect 12276 24847 12278 24867
rect 12324 24847 12326 24867
rect 12372 24847 12374 24867
rect 12420 24847 12422 24867
rect 12444 24847 12446 24867
rect 12468 24847 12470 24867
rect 12516 24847 12518 24867
rect 12540 24847 12542 24867
rect 12564 24847 12566 24867
rect 12660 24847 12662 24867
rect 12756 24847 12758 24867
rect 12828 24847 12830 24867
rect 12876 24847 12878 24867
rect 12972 24847 12974 24867
rect 13044 24847 13046 24867
rect 13068 24847 13070 24867
rect 13284 24847 13286 24867
rect 13332 24847 13334 24867
rect 13500 24847 13502 24867
rect 13572 24847 13574 24867
rect 13668 24847 13670 24867
rect 13716 24847 13718 24867
rect 13764 24847 13766 24867
rect 13860 24847 13862 24867
rect 13956 24847 13958 24867
rect 14004 24847 14006 24867
rect 14100 24847 14102 24867
rect 14940 24847 14942 24867
rect 15036 24847 15038 24867
rect 15135 24864 15149 24867
rect 15159 24867 19157 24871
rect 15159 24864 15173 24867
rect 15180 24864 15183 24867
rect 15276 24847 15278 24867
rect 15420 24847 15422 24867
rect 15492 24847 15494 24867
rect 15660 24847 15662 24867
rect 15708 24847 15710 24867
rect 15732 24847 15734 24867
rect 15756 24847 15758 24867
rect 15804 24847 15806 24867
rect 15828 24847 15830 24867
rect 15852 24847 15854 24867
rect 15948 24847 15950 24867
rect 15972 24847 15974 24867
rect 16044 24847 16046 24867
rect 16068 24847 16070 24867
rect 16164 24847 16166 24867
rect 16260 24847 16262 24867
rect 16332 24847 16334 24867
rect 16380 24847 16382 24867
rect 16476 24847 16478 24867
rect 16548 24847 16550 24867
rect 16572 24847 16574 24867
rect 16620 24847 16622 24867
rect 16668 24847 16670 24867
rect 16716 24847 16718 24867
rect 16764 24847 16766 24867
rect 16812 24847 16814 24867
rect 16884 24847 16886 24867
rect 16908 24847 16910 24867
rect 16980 24847 16982 24867
rect 17148 24847 17150 24867
rect 17196 24847 17198 24867
rect 17220 24847 17222 24867
rect 17292 24847 17294 24867
rect 17316 24847 17318 24867
rect 18132 24847 18134 24867
rect 18228 24847 18230 24867
rect 18433 24847 18491 24848
rect 18492 24847 18494 24867
rect 18495 24864 18509 24867
rect 18591 24864 18605 24867
rect 18612 24864 18615 24867
rect 18636 24847 18638 24867
rect 18732 24847 18734 24867
rect 18828 24847 18830 24867
rect 18879 24864 18893 24867
rect 18900 24864 18903 24867
rect 18924 24847 18926 24867
rect 18972 24847 18974 24867
rect 19020 24847 19022 24867
rect 19068 24847 19070 24867
rect 19140 24847 19142 24867
rect 19143 24864 19157 24867
rect 19164 24867 23339 24871
rect 19164 24864 19181 24867
rect 19164 24847 19166 24864
rect 19236 24847 19238 24867
rect 19260 24847 19262 24867
rect 19788 24847 19790 24867
rect 19836 24847 19838 24867
rect 19860 24847 19862 24867
rect 19884 24847 19886 24867
rect 19956 24847 19958 24867
rect 19980 24847 19982 24867
rect 19993 24862 19996 24867
rect 20003 24848 20006 24862
rect 20004 24847 20006 24848
rect 20052 24847 20054 24867
rect 20076 24847 20078 24867
rect 20124 24864 20126 24867
rect 20100 24847 20103 24864
rect 20124 24847 20127 24864
rect 20172 24847 20174 24867
rect 20196 24847 20198 24867
rect 20292 24847 20294 24867
rect 20388 24847 20390 24867
rect 20412 24847 20414 24867
rect 20508 24847 20510 24867
rect 20532 24847 20534 24867
rect 20604 24847 20606 24867
rect 20628 24847 20630 24867
rect 20823 24864 20837 24867
rect 20892 24847 20894 24867
rect 20964 24847 20966 24867
rect 20988 24847 20990 24867
rect 21108 24847 21110 24867
rect 21204 24847 21206 24867
rect 21300 24847 21302 24867
rect 21324 24847 21326 24867
rect 21444 24847 21446 24867
rect 21468 24847 21470 24867
rect 21564 24847 21566 24867
rect 21588 24847 21590 24867
rect 21684 24847 21686 24867
rect 21708 24847 21710 24867
rect 21828 24847 21830 24867
rect 21924 24847 21926 24867
rect 22068 24847 22070 24867
rect 22188 24847 22190 24867
rect 22212 24847 22214 24867
rect 22884 24847 22886 24867
rect 22980 24847 22982 24867
rect 23076 24847 23078 24867
rect 23100 24847 23102 24867
rect 23124 24847 23126 24867
rect 23244 24848 23246 24867
rect 23233 24847 23267 24848
rect -11975 24843 20093 24847
rect -11868 24840 -11866 24843
rect -11868 24824 -11865 24840
rect -11772 24824 -11770 24843
rect -11676 24824 -11674 24843
rect -11879 24823 -11845 24824
rect -11783 24823 -11725 24824
rect -11687 24823 -11653 24824
rect -11615 24823 -11581 24824
rect -11508 24823 -11506 24843
rect -11436 24823 -11434 24843
rect -11412 24823 -11410 24843
rect -11196 24823 -11194 24843
rect -11100 24823 -11098 24843
rect -9900 24823 -9898 24843
rect -9732 24823 -9730 24843
rect -9636 24823 -9634 24843
rect -9540 24823 -9538 24843
rect -9444 24823 -9442 24843
rect -9348 24823 -9346 24843
rect -9228 24823 -9226 24843
rect -9108 24823 -9106 24843
rect -9012 24823 -9010 24843
rect -8916 24823 -8914 24843
rect -8628 24823 -8626 24843
rect -8532 24823 -8530 24843
rect -8436 24823 -8434 24843
rect -8364 24823 -8362 24843
rect -8340 24823 -8338 24843
rect -8268 24823 -8266 24843
rect -8124 24823 -8122 24843
rect -7764 24823 -7762 24843
rect -7524 24823 -7522 24843
rect -7356 24823 -7354 24843
rect -7308 24823 -7306 24843
rect -7140 24823 -7138 24843
rect -7044 24823 -7042 24843
rect -6948 24823 -6946 24843
rect -6852 24823 -6850 24843
rect -6732 24823 -6730 24843
rect -6516 24823 -6514 24843
rect -5892 24823 -5890 24843
rect -5436 24823 -5434 24843
rect -5340 24823 -5338 24843
rect -5196 24823 -5194 24843
rect -4716 24823 -4714 24843
rect -4500 24823 -4498 24843
rect -4404 24823 -4402 24843
rect -4308 24823 -4306 24843
rect -4164 24823 -4162 24843
rect -3876 24823 -3874 24843
rect -3540 24823 -3538 24843
rect -3468 24823 -3466 24843
rect -3324 24823 -3322 24843
rect -3108 24823 -3106 24843
rect -3012 24823 -3010 24843
rect -2964 24823 -2962 24843
rect -2916 24823 -2914 24843
rect -2868 24823 -2866 24843
rect -2820 24823 -2818 24843
rect -2772 24823 -2770 24843
rect -2676 24823 -2674 24843
rect -2364 24823 -2362 24843
rect -2316 24823 -2314 24843
rect -2076 24823 -2074 24843
rect -1980 24823 -1978 24843
rect -1812 24823 -1810 24843
rect -1572 24823 -1570 24843
rect -1476 24823 -1474 24843
rect -1356 24823 -1354 24843
rect -1260 24823 -1258 24843
rect -1236 24823 -1234 24843
rect -1140 24823 -1138 24843
rect -876 24823 -874 24843
rect -660 24823 -658 24843
rect -492 24823 -490 24843
rect -396 24823 -394 24843
rect -372 24823 -370 24843
rect -276 24823 -274 24843
rect -12 24823 -10 24843
rect 84 24823 86 24843
rect 156 24823 158 24843
rect 252 24823 254 24843
rect 348 24823 350 24843
rect 468 24823 470 24843
rect 492 24823 494 24843
rect 564 24823 566 24843
rect 588 24823 590 24843
rect 636 24823 638 24843
rect 660 24823 662 24843
rect 732 24823 734 24843
rect 948 24823 950 24843
rect 1044 24823 1046 24843
rect 1092 24823 1094 24843
rect 1140 24823 1142 24843
rect 1308 24823 1310 24843
rect 1356 24823 1358 24843
rect 1428 24823 1430 24843
rect 1692 24823 1694 24843
rect 1860 24823 1862 24843
rect 2076 24823 2078 24843
rect 2100 24823 2102 24843
rect 2244 24823 2246 24843
rect 2460 24823 2462 24843
rect 2772 24823 2774 24843
rect 2868 24823 2870 24843
rect 2940 24823 2942 24843
rect 3012 24823 3014 24843
rect 3108 24823 3110 24843
rect 3324 24823 3326 24843
rect 3396 24823 3398 24843
rect 3564 24823 3566 24843
rect 3660 24823 3662 24843
rect 3780 24823 3782 24843
rect 4092 24823 4094 24843
rect 4188 24823 4190 24843
rect 4308 24823 4310 24843
rect 4404 24823 4406 24843
rect 4500 24823 4502 24843
rect 4596 24823 4598 24843
rect 4692 24823 4694 24843
rect 4956 24823 4958 24843
rect 4980 24823 4982 24843
rect 5052 24823 5054 24843
rect 5124 24823 5126 24843
rect 5220 24823 5222 24843
rect 5257 24838 5260 24843
rect 5268 24838 5270 24843
rect 5267 24824 5270 24838
rect 5388 24823 5390 24843
rect 5484 24823 5486 24843
rect 5508 24823 5510 24843
rect 5532 24823 5534 24843
rect 5628 24823 5630 24843
rect 5652 24823 5654 24843
rect 5748 24823 5750 24843
rect 5796 24823 5798 24843
rect 5844 24823 5846 24843
rect 5892 24823 5894 24843
rect 6276 24823 6278 24843
rect 6372 24823 6374 24843
rect 6420 24823 6422 24843
rect 6492 24823 6494 24843
rect 6516 24823 6518 24843
rect 6588 24823 6590 24843
rect 6612 24823 6614 24843
rect 6684 24823 6686 24843
rect 6708 24823 6710 24843
rect 6780 24823 6782 24843
rect 6804 24823 6806 24843
rect 6900 24823 6902 24843
rect 6924 24823 6926 24843
rect 7020 24823 7022 24843
rect 7164 24823 7166 24843
rect 7177 24823 7235 24824
rect 7236 24823 7238 24843
rect 7308 24823 7310 24843
rect 7380 24823 7382 24843
rect 7404 24823 7406 24843
rect 7476 24823 7478 24843
rect 7500 24823 7502 24843
rect 7572 24823 7574 24843
rect 7644 24823 7646 24843
rect 7668 24823 7670 24843
rect 7908 24823 7910 24843
rect 8124 24823 8126 24843
rect 8220 24823 8222 24843
rect 8652 24823 8654 24843
rect 8700 24823 8702 24843
rect 8748 24823 8750 24843
rect 8796 24823 8798 24843
rect 8844 24823 8846 24843
rect 8868 24823 8870 24843
rect 9516 24823 9518 24843
rect 9660 24823 9662 24843
rect 9684 24823 9686 24843
rect 9756 24823 9758 24843
rect 9780 24823 9782 24843
rect 9804 24823 9806 24843
rect 9852 24823 9854 24843
rect 9948 24823 9950 24843
rect 10044 24823 10046 24843
rect 10116 24823 10118 24843
rect 10140 24823 10142 24843
rect 10188 24823 10190 24843
rect 10236 24823 10238 24843
rect 10284 24823 10286 24843
rect 10332 24823 10334 24843
rect 10380 24823 10382 24843
rect 10428 24823 10430 24843
rect 10476 24823 10478 24843
rect 10524 24823 10526 24843
rect 10620 24823 10622 24843
rect 10644 24823 10646 24843
rect 10716 24823 10718 24843
rect 10884 24823 10886 24843
rect 10956 24823 10958 24843
rect 11052 24823 11054 24843
rect 11100 24823 11102 24843
rect 11172 24823 11174 24843
rect 11220 24823 11222 24843
rect 11340 24823 11342 24843
rect 11436 24823 11438 24843
rect 11532 24823 11534 24843
rect 11628 24823 11630 24843
rect 11676 24823 11678 24843
rect 11724 24823 11726 24843
rect 11772 24823 11774 24843
rect 11796 24823 11798 24843
rect 11892 24823 11894 24843
rect 11988 24823 11990 24843
rect 12060 24823 12062 24843
rect 12276 24823 12278 24843
rect 12324 24823 12326 24843
rect 12372 24823 12374 24843
rect 12420 24823 12422 24843
rect 12444 24823 12446 24843
rect 12468 24823 12470 24843
rect 12516 24823 12518 24843
rect 12540 24823 12542 24843
rect 12564 24823 12566 24843
rect 12660 24823 12662 24843
rect 12756 24823 12758 24843
rect 12828 24823 12830 24843
rect 12876 24823 12878 24843
rect 12972 24823 12974 24843
rect 13044 24823 13046 24843
rect 13068 24823 13070 24843
rect 13284 24823 13286 24843
rect 13332 24823 13334 24843
rect 13500 24823 13502 24843
rect 13572 24823 13574 24843
rect 13668 24823 13670 24843
rect 13716 24823 13718 24843
rect 13764 24823 13766 24843
rect 13860 24823 13862 24843
rect 13956 24823 13958 24843
rect 14004 24823 14006 24843
rect 14100 24823 14102 24843
rect 14940 24823 14942 24843
rect 15036 24823 15038 24843
rect 15276 24823 15278 24843
rect 15420 24823 15422 24843
rect 15492 24824 15494 24843
rect 15457 24823 15515 24824
rect 15660 24823 15662 24843
rect 15708 24823 15710 24843
rect 15732 24823 15734 24843
rect 15756 24823 15758 24843
rect 15804 24823 15806 24843
rect 15828 24823 15830 24843
rect 15852 24823 15854 24843
rect 15948 24823 15950 24843
rect 15972 24823 15974 24843
rect 16044 24823 16046 24843
rect 16068 24823 16070 24843
rect 16164 24823 16166 24843
rect 16260 24823 16262 24843
rect 16332 24823 16334 24843
rect 16380 24823 16382 24843
rect 16476 24823 16478 24843
rect 16548 24823 16550 24843
rect 16572 24823 16574 24843
rect 16620 24823 16622 24843
rect 16668 24823 16670 24843
rect 16716 24823 16718 24843
rect 16764 24823 16766 24843
rect 16812 24823 16814 24843
rect 16884 24823 16886 24843
rect 16908 24823 16910 24843
rect 16980 24823 16982 24843
rect 17148 24823 17150 24843
rect 17196 24823 17198 24843
rect 17220 24823 17222 24843
rect 17292 24823 17294 24843
rect 17316 24823 17318 24843
rect 18132 24823 18134 24843
rect 18228 24823 18230 24843
rect 18492 24823 18494 24843
rect 18540 24823 18543 24840
rect 18636 24823 18638 24843
rect 18732 24823 18734 24843
rect 18828 24823 18830 24843
rect 18924 24823 18926 24843
rect 18972 24823 18974 24843
rect 19020 24823 19022 24843
rect 19068 24823 19070 24843
rect 19140 24823 19142 24843
rect 19164 24823 19166 24843
rect 19236 24823 19238 24843
rect 19260 24823 19262 24843
rect 19788 24823 19790 24843
rect 19836 24823 19838 24843
rect 19860 24823 19862 24843
rect 19884 24823 19886 24843
rect 19956 24823 19958 24843
rect 19980 24823 19982 24843
rect 20004 24823 20006 24843
rect 20052 24823 20054 24843
rect 20076 24823 20078 24843
rect 20079 24840 20093 24843
rect 20100 24843 23267 24847
rect 20100 24840 20117 24843
rect 20124 24840 20127 24843
rect 20100 24823 20102 24840
rect 20172 24823 20174 24843
rect 20196 24823 20198 24843
rect 20292 24823 20294 24843
rect 20388 24823 20390 24843
rect 20412 24823 20414 24843
rect 20508 24823 20510 24843
rect 20532 24823 20534 24843
rect 20604 24823 20606 24843
rect 20628 24823 20630 24843
rect 20892 24823 20894 24843
rect 20964 24823 20966 24843
rect 20988 24823 20990 24843
rect 21108 24823 21110 24843
rect 21204 24823 21206 24843
rect 21300 24823 21302 24843
rect 21324 24823 21326 24843
rect 21444 24823 21446 24843
rect 21468 24823 21470 24843
rect 21564 24823 21566 24843
rect 21588 24823 21590 24843
rect 21684 24823 21686 24843
rect 21708 24823 21710 24843
rect 21828 24824 21830 24843
rect 21817 24823 21851 24824
rect 21924 24823 21926 24843
rect 22068 24823 22070 24843
rect 22188 24823 22190 24843
rect 22212 24823 22214 24843
rect 22884 24823 22886 24843
rect 22980 24823 22982 24843
rect 23076 24823 23078 24843
rect 23100 24823 23102 24843
rect 23124 24823 23126 24843
rect 23233 24838 23236 24843
rect 23244 24838 23246 24843
rect 23243 24824 23246 24838
rect 23137 24823 23171 24824
rect -11879 24819 5333 24823
rect -11879 24816 -11875 24819
rect -11868 24816 -11865 24819
rect -11783 24814 -11780 24819
rect -11772 24816 -11770 24819
rect -11772 24814 -11769 24816
rect -11687 24814 -11684 24819
rect -11676 24816 -11674 24819
rect -11508 24816 -11506 24819
rect -11676 24814 -11673 24816
rect -11773 24800 -11769 24814
rect -11677 24806 -11673 24814
rect -11663 24806 -11659 24814
rect -11591 24806 -11587 24814
rect -11677 24800 -11663 24806
rect -11601 24800 -11591 24806
rect -11508 24800 -11505 24816
rect -11436 24800 -11434 24819
rect -11412 24800 -11410 24819
rect -11616 24795 -11550 24799
rect -11601 24792 -11587 24795
rect -11543 24790 -11540 24800
rect -11529 24799 -11485 24800
rect -11447 24799 -11389 24800
rect -11196 24799 -11194 24819
rect -11100 24799 -11098 24819
rect -9900 24799 -9898 24819
rect -9732 24799 -9730 24819
rect -9636 24799 -9634 24819
rect -9540 24799 -9538 24819
rect -9444 24799 -9442 24819
rect -9348 24799 -9346 24819
rect -9228 24799 -9226 24819
rect -9108 24799 -9106 24819
rect -9012 24799 -9010 24819
rect -8916 24799 -8914 24819
rect -8628 24799 -8626 24819
rect -8532 24799 -8530 24819
rect -8436 24799 -8434 24819
rect -8364 24799 -8362 24819
rect -8340 24799 -8338 24819
rect -8268 24799 -8266 24819
rect -8124 24799 -8122 24819
rect -7764 24799 -7762 24819
rect -7524 24799 -7522 24819
rect -7356 24799 -7354 24819
rect -7308 24799 -7306 24819
rect -7140 24799 -7138 24819
rect -7044 24799 -7042 24819
rect -6948 24799 -6946 24819
rect -6852 24799 -6850 24819
rect -6732 24799 -6730 24819
rect -6516 24799 -6514 24819
rect -5892 24799 -5890 24819
rect -5436 24799 -5434 24819
rect -5340 24799 -5338 24819
rect -5196 24799 -5194 24819
rect -4716 24799 -4714 24819
rect -4500 24799 -4498 24819
rect -4404 24799 -4402 24819
rect -4308 24799 -4306 24819
rect -4164 24799 -4162 24819
rect -3876 24799 -3874 24819
rect -3540 24799 -3538 24819
rect -3468 24799 -3466 24819
rect -3324 24799 -3322 24819
rect -3108 24799 -3106 24819
rect -3012 24799 -3010 24819
rect -2964 24799 -2962 24819
rect -2916 24799 -2914 24819
rect -2868 24799 -2866 24819
rect -2820 24799 -2818 24819
rect -2772 24799 -2770 24819
rect -2676 24799 -2674 24819
rect -2364 24799 -2362 24819
rect -2316 24799 -2314 24819
rect -2135 24799 -2077 24800
rect -2076 24799 -2074 24819
rect -1980 24799 -1978 24819
rect -1812 24799 -1810 24819
rect -1572 24799 -1570 24819
rect -1476 24799 -1474 24819
rect -1356 24799 -1354 24819
rect -1260 24799 -1258 24819
rect -1236 24799 -1234 24819
rect -1140 24799 -1138 24819
rect -876 24799 -874 24819
rect -660 24799 -658 24819
rect -492 24799 -490 24819
rect -396 24799 -394 24819
rect -372 24799 -370 24819
rect -276 24799 -274 24819
rect -12 24799 -10 24819
rect 84 24799 86 24819
rect 156 24799 158 24819
rect 252 24799 254 24819
rect 348 24799 350 24819
rect 468 24799 470 24819
rect 492 24799 494 24819
rect 564 24799 566 24819
rect 588 24799 590 24819
rect 636 24799 638 24819
rect 660 24799 662 24819
rect 732 24799 734 24819
rect 948 24799 950 24819
rect 1044 24799 1046 24819
rect 1092 24799 1094 24819
rect 1140 24799 1142 24819
rect 1308 24799 1310 24819
rect 1356 24799 1358 24819
rect 1428 24799 1430 24819
rect 1692 24799 1694 24819
rect 1860 24799 1862 24819
rect 2076 24800 2078 24819
rect 2041 24799 2099 24800
rect 2100 24799 2102 24819
rect 2244 24799 2246 24819
rect 2460 24799 2462 24819
rect 2772 24799 2774 24819
rect 2868 24799 2870 24819
rect 2940 24799 2942 24819
rect 3012 24800 3014 24819
rect 2977 24799 3035 24800
rect 3108 24799 3110 24819
rect 3324 24799 3326 24819
rect 3396 24799 3398 24819
rect 3564 24799 3566 24819
rect 3660 24799 3662 24819
rect 3780 24799 3782 24819
rect 4092 24799 4094 24819
rect 4188 24799 4190 24819
rect 4308 24799 4310 24819
rect 4404 24799 4406 24819
rect 4500 24799 4502 24819
rect 4596 24799 4598 24819
rect 4692 24799 4694 24819
rect 4956 24799 4958 24819
rect 4980 24799 4982 24819
rect 5052 24799 5054 24819
rect 5124 24799 5126 24819
rect 5220 24799 5222 24819
rect 5319 24816 5333 24819
rect 5343 24819 18533 24823
rect 5343 24816 5357 24819
rect 5388 24799 5390 24819
rect 5484 24799 5486 24819
rect 5508 24799 5510 24819
rect 5532 24799 5534 24819
rect 5628 24799 5630 24819
rect 5652 24799 5654 24819
rect 5748 24799 5750 24819
rect 5796 24799 5798 24819
rect 5844 24799 5846 24819
rect 5892 24799 5894 24819
rect 6276 24799 6278 24819
rect 6372 24799 6374 24819
rect 6420 24799 6422 24819
rect 6492 24799 6494 24819
rect 6516 24799 6518 24819
rect 6588 24799 6590 24819
rect 6612 24799 6614 24819
rect 6684 24799 6686 24819
rect 6708 24799 6710 24819
rect 6780 24799 6782 24819
rect 6804 24799 6806 24819
rect 6900 24799 6902 24819
rect 6924 24799 6926 24819
rect 7020 24799 7022 24819
rect 7164 24799 7166 24819
rect 7236 24799 7238 24819
rect 7308 24816 7310 24819
rect 7284 24799 7287 24816
rect 7308 24799 7311 24816
rect 7380 24799 7382 24819
rect 7404 24799 7406 24819
rect 7476 24799 7478 24819
rect 7500 24799 7502 24819
rect 7572 24799 7574 24819
rect 7644 24799 7646 24819
rect 7668 24799 7670 24819
rect 7908 24799 7910 24819
rect 8124 24799 8126 24819
rect 8220 24799 8222 24819
rect 8652 24799 8654 24819
rect 8700 24799 8702 24819
rect 8748 24799 8750 24819
rect 8796 24799 8798 24819
rect 8844 24799 8846 24819
rect 8868 24799 8870 24819
rect 9516 24799 9518 24819
rect 9660 24799 9662 24819
rect 9684 24799 9686 24819
rect 9756 24799 9758 24819
rect 9780 24799 9782 24819
rect 9804 24799 9806 24819
rect 9852 24799 9854 24819
rect 9948 24799 9950 24819
rect 10044 24799 10046 24819
rect 10116 24800 10118 24819
rect 10105 24799 10139 24800
rect 10140 24799 10142 24819
rect 10188 24799 10190 24819
rect 10236 24799 10238 24819
rect 10284 24799 10286 24819
rect 10332 24799 10334 24819
rect 10380 24799 10382 24819
rect 10428 24799 10430 24819
rect 10476 24800 10478 24819
rect 10441 24799 10499 24800
rect 10524 24799 10526 24819
rect 10620 24799 10622 24819
rect 10644 24799 10646 24819
rect 10716 24799 10718 24819
rect 10884 24799 10886 24819
rect 10956 24799 10958 24819
rect 11052 24799 11054 24819
rect 11100 24799 11102 24819
rect 11172 24799 11174 24819
rect 11220 24799 11222 24819
rect 11340 24799 11342 24819
rect 11436 24799 11438 24819
rect 11532 24799 11534 24819
rect 11628 24799 11630 24819
rect 11676 24799 11678 24819
rect 11724 24799 11726 24819
rect 11772 24799 11774 24819
rect 11796 24799 11798 24819
rect 11892 24799 11894 24819
rect 11988 24799 11990 24819
rect 12060 24799 12062 24819
rect 12276 24799 12278 24819
rect 12324 24799 12326 24819
rect 12372 24799 12374 24819
rect 12420 24799 12422 24819
rect 12444 24799 12446 24819
rect 12468 24799 12470 24819
rect 12516 24799 12518 24819
rect 12540 24799 12542 24819
rect 12564 24799 12566 24819
rect 12660 24799 12662 24819
rect 12756 24799 12758 24819
rect 12828 24799 12830 24819
rect 12876 24799 12878 24819
rect 12972 24799 12974 24819
rect 13044 24799 13046 24819
rect 13068 24799 13070 24819
rect 13284 24799 13286 24819
rect 13332 24799 13334 24819
rect 13500 24799 13502 24819
rect 13572 24799 13574 24819
rect 13668 24799 13670 24819
rect 13716 24799 13718 24819
rect 13764 24799 13766 24819
rect 13860 24799 13862 24819
rect 13956 24799 13958 24819
rect 14004 24799 14006 24819
rect 14100 24799 14102 24819
rect 14940 24799 14942 24819
rect 15036 24799 15038 24819
rect 15276 24799 15278 24819
rect 15420 24799 15422 24819
rect 15481 24814 15484 24819
rect 15492 24814 15494 24819
rect 15491 24800 15494 24814
rect 15564 24799 15567 24816
rect 15660 24799 15662 24819
rect 15708 24799 15710 24819
rect 15732 24799 15734 24819
rect 15756 24799 15758 24819
rect 15804 24799 15806 24819
rect 15828 24799 15830 24819
rect 15852 24799 15854 24819
rect 15948 24799 15950 24819
rect 15972 24799 15974 24819
rect 16044 24799 16046 24819
rect 16068 24799 16070 24819
rect 16164 24799 16166 24819
rect 16260 24799 16262 24819
rect 16332 24799 16334 24819
rect 16380 24799 16382 24819
rect 16476 24799 16478 24819
rect 16548 24799 16550 24819
rect 16572 24799 16574 24819
rect 16620 24799 16622 24819
rect 16668 24799 16670 24819
rect 16716 24799 16718 24819
rect 16764 24799 16766 24819
rect 16812 24799 16814 24819
rect 16884 24799 16886 24819
rect 16908 24799 16910 24819
rect 16980 24799 16982 24819
rect 17017 24799 17075 24800
rect 17148 24799 17150 24819
rect 17196 24799 17198 24819
rect 17220 24799 17222 24819
rect 17292 24799 17294 24819
rect 17316 24799 17318 24819
rect 18132 24799 18134 24819
rect 18228 24799 18230 24819
rect 18492 24799 18494 24819
rect 18519 24816 18533 24819
rect 18540 24819 23171 24823
rect 18540 24816 18557 24819
rect 18540 24799 18542 24816
rect 18636 24799 18638 24819
rect 18732 24799 18734 24819
rect 18828 24799 18830 24819
rect 18924 24799 18926 24819
rect 18972 24799 18974 24819
rect 19020 24799 19022 24819
rect 19068 24799 19070 24819
rect 19140 24799 19142 24819
rect 19164 24799 19166 24819
rect 19236 24799 19238 24819
rect 19260 24799 19262 24819
rect 19788 24799 19790 24819
rect 19836 24799 19838 24819
rect 19860 24799 19862 24819
rect 19884 24799 19886 24819
rect 19956 24799 19958 24819
rect 19980 24799 19982 24819
rect 20004 24799 20006 24819
rect 20052 24799 20054 24819
rect 20076 24799 20078 24819
rect 20100 24799 20102 24819
rect 20172 24799 20174 24819
rect 20196 24799 20198 24819
rect 20292 24799 20294 24819
rect 20388 24799 20390 24819
rect 20412 24799 20414 24819
rect 20508 24799 20510 24819
rect 20532 24799 20534 24819
rect 20604 24799 20606 24819
rect 20628 24799 20630 24819
rect 20892 24799 20894 24819
rect 20964 24799 20966 24819
rect 20988 24799 20990 24819
rect 21108 24799 21110 24819
rect 21204 24799 21206 24819
rect 21300 24799 21302 24819
rect 21324 24799 21326 24819
rect 21444 24799 21446 24819
rect 21468 24799 21470 24819
rect 21564 24799 21566 24819
rect 21588 24799 21590 24819
rect 21684 24799 21686 24819
rect 21708 24799 21710 24819
rect 21817 24814 21820 24819
rect 21828 24814 21830 24819
rect 21827 24800 21830 24814
rect 21924 24816 21926 24819
rect 21924 24799 21927 24816
rect 22068 24799 22070 24819
rect 22188 24799 22190 24819
rect 22212 24799 22214 24819
rect 22884 24799 22886 24819
rect 22980 24799 22982 24819
rect 23076 24799 23078 24819
rect 23100 24799 23102 24819
rect 23124 24800 23126 24819
rect 23113 24799 23147 24800
rect -11529 24795 7277 24799
rect -11529 24792 -11515 24795
rect -11508 24792 -11505 24795
rect -11447 24790 -11444 24795
rect -11436 24792 -11434 24795
rect -11436 24790 -11433 24792
rect -11533 24789 -11530 24790
rect -11437 24782 -11433 24790
rect -11423 24790 -11420 24795
rect -11412 24792 -11410 24795
rect -11412 24790 -11409 24792
rect -11423 24782 -11419 24790
rect -11437 24776 -11423 24782
rect -11413 24776 -11409 24790
rect -11303 24775 -11269 24776
rect -11196 24775 -11194 24795
rect -11100 24775 -11098 24795
rect -9900 24775 -9898 24795
rect -9732 24775 -9730 24795
rect -9636 24775 -9634 24795
rect -9540 24775 -9538 24795
rect -9444 24775 -9442 24795
rect -9348 24775 -9346 24795
rect -9228 24775 -9226 24795
rect -9108 24775 -9106 24795
rect -9012 24775 -9010 24795
rect -8916 24775 -8914 24795
rect -8628 24775 -8626 24795
rect -8532 24775 -8530 24795
rect -8436 24775 -8434 24795
rect -8364 24776 -8362 24795
rect -8375 24775 -8341 24776
rect -8340 24775 -8338 24795
rect -8268 24775 -8266 24795
rect -8124 24775 -8122 24795
rect -7764 24775 -7762 24795
rect -7524 24775 -7522 24795
rect -7356 24775 -7354 24795
rect -7308 24775 -7306 24795
rect -7140 24775 -7138 24795
rect -7044 24775 -7042 24795
rect -6948 24775 -6946 24795
rect -6852 24775 -6850 24795
rect -6732 24775 -6730 24795
rect -6516 24775 -6514 24795
rect -5892 24775 -5890 24795
rect -5436 24775 -5434 24795
rect -5340 24775 -5338 24795
rect -5196 24775 -5194 24795
rect -4716 24775 -4714 24795
rect -4500 24775 -4498 24795
rect -4404 24775 -4402 24795
rect -4308 24775 -4306 24795
rect -4164 24775 -4162 24795
rect -3876 24775 -3874 24795
rect -3540 24775 -3538 24795
rect -3468 24775 -3466 24795
rect -3324 24775 -3322 24795
rect -3108 24775 -3106 24795
rect -3012 24775 -3010 24795
rect -2964 24775 -2962 24795
rect -2916 24775 -2914 24795
rect -2868 24775 -2866 24795
rect -2820 24775 -2818 24795
rect -2772 24775 -2770 24795
rect -2676 24775 -2674 24795
rect -2364 24775 -2362 24795
rect -2316 24775 -2314 24795
rect -2076 24775 -2074 24795
rect -1980 24775 -1978 24795
rect -1812 24775 -1810 24795
rect -1572 24775 -1570 24795
rect -1476 24775 -1474 24795
rect -1356 24775 -1354 24795
rect -1260 24775 -1258 24795
rect -1236 24775 -1234 24795
rect -1140 24775 -1138 24795
rect -876 24775 -874 24795
rect -660 24775 -658 24795
rect -492 24775 -490 24795
rect -396 24775 -394 24795
rect -372 24775 -370 24795
rect -276 24775 -274 24795
rect -12 24775 -10 24795
rect 84 24775 86 24795
rect 156 24775 158 24795
rect 252 24775 254 24795
rect 348 24775 350 24795
rect 468 24775 470 24795
rect 492 24775 494 24795
rect 564 24775 566 24795
rect 588 24775 590 24795
rect 636 24775 638 24795
rect 660 24775 662 24795
rect 732 24775 734 24795
rect 948 24775 950 24795
rect 1044 24775 1046 24795
rect 1092 24775 1094 24795
rect 1140 24775 1142 24795
rect 1308 24775 1310 24795
rect 1356 24775 1358 24795
rect 1428 24775 1430 24795
rect 1692 24775 1694 24795
rect 1860 24775 1862 24795
rect 2065 24790 2068 24795
rect 2076 24790 2078 24795
rect 2075 24776 2078 24790
rect 1993 24775 2027 24776
rect 2100 24775 2102 24795
rect 2148 24775 2151 24792
rect 2244 24775 2246 24795
rect 2460 24775 2462 24795
rect 2772 24775 2774 24795
rect 2868 24775 2870 24795
rect 2940 24775 2942 24795
rect 2977 24790 2980 24795
rect 3001 24790 3004 24795
rect 3012 24790 3014 24795
rect 2987 24776 2990 24790
rect 3011 24776 3014 24790
rect 3108 24792 3110 24795
rect 2988 24775 2990 24776
rect 3108 24775 3111 24792
rect 3324 24775 3326 24795
rect 3396 24775 3398 24795
rect 3564 24775 3566 24795
rect 3660 24775 3662 24795
rect 3780 24775 3782 24795
rect 4092 24775 4094 24795
rect 4188 24775 4190 24795
rect 4308 24775 4310 24795
rect 4404 24775 4406 24795
rect 4500 24775 4502 24795
rect 4596 24775 4598 24795
rect 4692 24775 4694 24795
rect 4897 24775 4931 24776
rect 4956 24775 4958 24795
rect 4980 24775 4982 24795
rect 5052 24775 5054 24795
rect 5124 24775 5126 24795
rect 5220 24775 5222 24795
rect 5388 24775 5390 24795
rect 5484 24775 5486 24795
rect 5508 24775 5510 24795
rect 5532 24775 5534 24795
rect 5628 24775 5630 24795
rect 5652 24775 5654 24795
rect 5748 24775 5750 24795
rect 5796 24775 5798 24795
rect 5844 24775 5846 24795
rect 5892 24775 5894 24795
rect 6276 24775 6278 24795
rect 6372 24775 6374 24795
rect 6420 24775 6422 24795
rect 6492 24775 6494 24795
rect 6516 24775 6518 24795
rect 6588 24775 6590 24795
rect 6612 24775 6614 24795
rect 6684 24775 6686 24795
rect 6708 24775 6710 24795
rect 6780 24775 6782 24795
rect 6804 24775 6806 24795
rect 6900 24775 6902 24795
rect 6924 24775 6926 24795
rect 7020 24775 7022 24795
rect 7164 24775 7166 24795
rect 7236 24775 7238 24795
rect 7263 24792 7277 24795
rect 7284 24795 15557 24799
rect 7284 24792 7301 24795
rect 7308 24792 7311 24795
rect 7284 24775 7286 24792
rect 7380 24775 7382 24795
rect 7404 24775 7406 24795
rect 7476 24775 7478 24795
rect 7500 24775 7502 24795
rect 7572 24775 7574 24795
rect 7644 24775 7646 24795
rect 7668 24775 7670 24795
rect 7908 24775 7910 24795
rect 8124 24775 8126 24795
rect 8220 24775 8222 24795
rect 8652 24775 8654 24795
rect 8700 24775 8702 24795
rect 8748 24775 8750 24795
rect 8796 24775 8798 24795
rect 8844 24775 8846 24795
rect 8868 24775 8870 24795
rect 9516 24775 9518 24795
rect 9660 24775 9662 24795
rect 9684 24775 9686 24795
rect 9756 24775 9758 24795
rect 9780 24775 9782 24795
rect 9804 24775 9806 24795
rect 9852 24775 9854 24795
rect 9948 24775 9950 24795
rect 10044 24775 10046 24795
rect 10105 24790 10108 24795
rect 10116 24790 10118 24795
rect 10115 24776 10118 24790
rect 10081 24775 10115 24776
rect 10140 24775 10142 24795
rect 10188 24776 10190 24795
rect 10177 24775 10211 24776
rect 10236 24775 10238 24795
rect 10284 24775 10286 24795
rect 10332 24775 10334 24795
rect 10380 24775 10382 24795
rect 10428 24775 10430 24795
rect 10465 24790 10468 24795
rect 10476 24790 10478 24795
rect 10475 24776 10478 24790
rect 10524 24775 10526 24795
rect 10548 24775 10551 24792
rect 10620 24775 10622 24795
rect 10644 24775 10646 24795
rect 10716 24775 10718 24795
rect 10884 24775 10886 24795
rect 10956 24775 10958 24795
rect 11052 24775 11054 24795
rect 11100 24775 11102 24795
rect 11172 24775 11174 24795
rect 11220 24775 11222 24795
rect 11340 24775 11342 24795
rect 11436 24775 11438 24795
rect 11532 24775 11534 24795
rect 11628 24775 11630 24795
rect 11676 24775 11678 24795
rect 11724 24775 11726 24795
rect 11772 24775 11774 24795
rect 11796 24775 11798 24795
rect 11892 24776 11894 24795
rect 11881 24775 11915 24776
rect 11988 24775 11990 24795
rect 12060 24775 12062 24795
rect 12276 24775 12278 24795
rect 12324 24775 12326 24795
rect 12372 24775 12374 24795
rect 12420 24775 12422 24795
rect 12444 24775 12446 24795
rect 12468 24775 12470 24795
rect 12516 24776 12518 24795
rect 12505 24775 12539 24776
rect 12540 24775 12542 24795
rect 12564 24775 12566 24795
rect 12660 24775 12662 24795
rect 12756 24775 12758 24795
rect 12828 24775 12830 24795
rect 12876 24775 12878 24795
rect 12972 24775 12974 24795
rect 13044 24775 13046 24795
rect 13068 24775 13070 24795
rect 13284 24775 13286 24795
rect 13332 24775 13334 24795
rect 13500 24775 13502 24795
rect 13572 24775 13574 24795
rect 13668 24775 13670 24795
rect 13716 24775 13718 24795
rect 13764 24775 13766 24795
rect 13860 24775 13862 24795
rect 13956 24775 13958 24795
rect 14004 24775 14006 24795
rect 14100 24775 14102 24795
rect 14940 24775 14942 24795
rect 15036 24775 15038 24795
rect 15276 24775 15278 24795
rect 15420 24775 15422 24795
rect 15543 24792 15557 24795
rect 15564 24795 23147 24799
rect 15564 24792 15581 24795
rect 15564 24775 15566 24792
rect 15660 24775 15662 24795
rect 15708 24775 15710 24795
rect 15732 24775 15734 24795
rect 15756 24775 15758 24795
rect 15804 24775 15806 24795
rect 15828 24775 15830 24795
rect 15852 24775 15854 24795
rect 15948 24775 15950 24795
rect 15972 24775 15974 24795
rect 16044 24775 16046 24795
rect 16068 24775 16070 24795
rect 16164 24775 16166 24795
rect 16260 24775 16262 24795
rect 16332 24775 16334 24795
rect 16380 24775 16382 24795
rect 16476 24775 16478 24795
rect 16548 24775 16550 24795
rect 16572 24775 16574 24795
rect 16620 24775 16622 24795
rect 16668 24775 16670 24795
rect 16716 24775 16718 24795
rect 16764 24775 16766 24795
rect 16812 24775 16814 24795
rect 16884 24775 16886 24795
rect 16908 24775 16910 24795
rect 16980 24775 16982 24795
rect 17017 24790 17020 24795
rect 17148 24792 17150 24795
rect 17027 24776 17030 24790
rect 17028 24775 17030 24776
rect 17124 24775 17127 24792
rect 17148 24775 17151 24792
rect 17196 24775 17198 24795
rect 17220 24775 17222 24795
rect 17292 24775 17294 24795
rect 17316 24775 17318 24795
rect 17953 24775 18011 24776
rect 18132 24775 18134 24795
rect 18228 24775 18230 24795
rect 18492 24775 18494 24795
rect 18540 24775 18542 24795
rect 18636 24775 18638 24795
rect 18732 24775 18734 24795
rect 18828 24775 18830 24795
rect 18924 24775 18926 24795
rect 18972 24775 18974 24795
rect 19020 24775 19022 24795
rect 19068 24775 19070 24795
rect 19140 24775 19142 24795
rect 19164 24775 19166 24795
rect 19236 24775 19238 24795
rect 19260 24775 19262 24795
rect 19788 24775 19790 24795
rect 19836 24775 19838 24795
rect 19860 24775 19862 24795
rect 19884 24775 19886 24795
rect 19956 24775 19958 24795
rect 19980 24775 19982 24795
rect 20004 24775 20006 24795
rect 20052 24775 20054 24795
rect 20076 24775 20078 24795
rect 20100 24775 20102 24795
rect 20172 24775 20174 24795
rect 20196 24775 20198 24795
rect 20292 24775 20294 24795
rect 20388 24775 20390 24795
rect 20412 24775 20414 24795
rect 20508 24775 20510 24795
rect 20532 24775 20534 24795
rect 20604 24775 20606 24795
rect 20628 24775 20630 24795
rect 20892 24775 20894 24795
rect 20964 24775 20966 24795
rect 20988 24775 20990 24795
rect 21108 24775 21110 24795
rect 21204 24775 21206 24795
rect 21300 24775 21302 24795
rect 21324 24775 21326 24795
rect 21444 24775 21446 24795
rect 21468 24775 21470 24795
rect 21564 24775 21566 24795
rect 21588 24775 21590 24795
rect 21684 24775 21686 24795
rect 21708 24775 21710 24795
rect 21903 24792 21917 24795
rect 21924 24792 21927 24795
rect 22068 24775 22070 24795
rect 22188 24775 22190 24795
rect 22212 24775 22214 24795
rect 22884 24775 22886 24795
rect 22980 24775 22982 24795
rect 23076 24775 23078 24795
rect 23100 24776 23102 24795
rect 23113 24790 23116 24795
rect 23124 24790 23126 24795
rect 23123 24776 23126 24790
rect 23089 24775 23123 24776
rect -11303 24771 -2035 24775
rect -11196 24768 -11194 24771
rect -11196 24752 -11193 24768
rect -11207 24751 -11173 24752
rect -11100 24751 -11098 24771
rect -9900 24751 -9898 24771
rect -9732 24751 -9730 24771
rect -9636 24751 -9634 24771
rect -9540 24751 -9538 24771
rect -9444 24751 -9442 24771
rect -9348 24751 -9346 24771
rect -9228 24751 -9226 24771
rect -9108 24751 -9106 24771
rect -9012 24751 -9010 24771
rect -8916 24751 -8914 24771
rect -8628 24751 -8626 24771
rect -8532 24751 -8530 24771
rect -8436 24751 -8434 24771
rect -8375 24766 -8372 24771
rect -8364 24766 -8362 24771
rect -8365 24752 -8362 24766
rect -8340 24751 -8338 24771
rect -8268 24768 -8266 24771
rect -8268 24751 -8265 24768
rect -8124 24751 -8122 24771
rect -7764 24751 -7762 24771
rect -7524 24751 -7522 24771
rect -7356 24751 -7354 24771
rect -7308 24751 -7306 24771
rect -7140 24751 -7138 24771
rect -7044 24751 -7042 24771
rect -6948 24751 -6946 24771
rect -6852 24751 -6850 24771
rect -6732 24751 -6730 24771
rect -6516 24751 -6514 24771
rect -5892 24751 -5890 24771
rect -5436 24751 -5434 24771
rect -5340 24751 -5338 24771
rect -5196 24751 -5194 24771
rect -4716 24751 -4714 24771
rect -4500 24751 -4498 24771
rect -4404 24751 -4402 24771
rect -4308 24751 -4306 24771
rect -4164 24751 -4162 24771
rect -3876 24751 -3874 24771
rect -3540 24751 -3538 24771
rect -3468 24751 -3466 24771
rect -3324 24751 -3322 24771
rect -3108 24751 -3106 24771
rect -3012 24751 -3010 24771
rect -2964 24751 -2962 24771
rect -2916 24751 -2914 24771
rect -2868 24751 -2866 24771
rect -2820 24751 -2818 24771
rect -2772 24751 -2770 24771
rect -2676 24751 -2674 24771
rect -2364 24751 -2362 24771
rect -2316 24751 -2314 24771
rect -2076 24751 -2074 24771
rect -2049 24768 -2035 24771
rect -2025 24771 2141 24775
rect -2025 24768 -2011 24771
rect -1980 24751 -1978 24771
rect -1812 24751 -1810 24771
rect -1572 24751 -1570 24771
rect -1476 24751 -1474 24771
rect -1356 24751 -1354 24771
rect -1260 24751 -1258 24771
rect -1236 24751 -1234 24771
rect -1140 24751 -1138 24771
rect -876 24751 -874 24771
rect -660 24751 -658 24771
rect -492 24751 -490 24771
rect -396 24751 -394 24771
rect -372 24751 -370 24771
rect -276 24751 -274 24771
rect -12 24751 -10 24771
rect 84 24751 86 24771
rect 156 24751 158 24771
rect 252 24751 254 24771
rect 348 24751 350 24771
rect 468 24751 470 24771
rect 492 24751 494 24771
rect 564 24751 566 24771
rect 588 24751 590 24771
rect 636 24751 638 24771
rect 660 24751 662 24771
rect 732 24751 734 24771
rect 948 24751 950 24771
rect 1044 24751 1046 24771
rect 1092 24751 1094 24771
rect 1140 24751 1142 24771
rect 1308 24751 1310 24771
rect 1356 24751 1358 24771
rect 1428 24751 1430 24771
rect 1692 24751 1694 24771
rect 1860 24751 1862 24771
rect 2100 24768 2102 24771
rect 2127 24768 2141 24771
rect 2148 24771 3077 24775
rect 2148 24768 2165 24771
rect 2100 24751 2103 24768
rect 2148 24751 2150 24768
rect 2244 24751 2246 24771
rect 2460 24751 2462 24771
rect 2772 24751 2774 24771
rect 2868 24751 2870 24771
rect 2940 24751 2942 24771
rect 2988 24751 2990 24771
rect 3063 24768 3077 24771
rect 3087 24771 10541 24775
rect 3087 24768 3101 24771
rect 3108 24768 3111 24771
rect 3324 24751 3326 24771
rect 3396 24751 3398 24771
rect 3564 24751 3566 24771
rect 3660 24751 3662 24771
rect 3780 24751 3782 24771
rect 4092 24751 4094 24771
rect 4188 24751 4190 24771
rect 4308 24751 4310 24771
rect 4404 24751 4406 24771
rect 4500 24751 4502 24771
rect 4596 24751 4598 24771
rect 4692 24751 4694 24771
rect 4956 24751 4958 24771
rect 4980 24751 4982 24771
rect 5052 24751 5054 24771
rect 5124 24751 5126 24771
rect 5220 24751 5222 24771
rect 5388 24751 5390 24771
rect 5484 24751 5486 24771
rect 5508 24751 5510 24771
rect 5532 24751 5534 24771
rect 5628 24751 5630 24771
rect 5652 24751 5654 24771
rect 5748 24751 5750 24771
rect 5796 24751 5798 24771
rect 5844 24751 5846 24771
rect 5892 24751 5894 24771
rect 6276 24751 6278 24771
rect 6372 24751 6374 24771
rect 6420 24751 6422 24771
rect 6492 24751 6494 24771
rect 6516 24751 6518 24771
rect 6588 24751 6590 24771
rect 6612 24751 6614 24771
rect 6684 24751 6686 24771
rect 6708 24751 6710 24771
rect 6780 24751 6782 24771
rect 6804 24751 6806 24771
rect 6900 24751 6902 24771
rect 6924 24751 6926 24771
rect 7020 24751 7022 24771
rect 7164 24751 7166 24771
rect 7236 24751 7238 24771
rect 7284 24751 7286 24771
rect 7380 24751 7382 24771
rect 7404 24751 7406 24771
rect 7476 24751 7478 24771
rect 7500 24751 7502 24771
rect 7572 24751 7574 24771
rect 7644 24751 7646 24771
rect 7668 24751 7670 24771
rect 7908 24751 7910 24771
rect 8124 24751 8126 24771
rect 8220 24751 8222 24771
rect 8652 24751 8654 24771
rect 8700 24751 8702 24771
rect 8748 24751 8750 24771
rect 8796 24751 8798 24771
rect 8844 24751 8846 24771
rect 8868 24751 8870 24771
rect 9516 24751 9518 24771
rect 9660 24751 9662 24771
rect 9684 24751 9686 24771
rect 9756 24751 9758 24771
rect 9780 24751 9782 24771
rect 9804 24751 9806 24771
rect 9852 24751 9854 24771
rect 9948 24751 9950 24771
rect 10044 24751 10046 24771
rect 10140 24751 10142 24771
rect 10177 24766 10180 24771
rect 10188 24768 10190 24771
rect 10191 24768 10205 24771
rect 10188 24766 10191 24768
rect 10187 24752 10191 24766
rect 10236 24751 10238 24771
rect 10284 24768 10286 24771
rect 10284 24751 10287 24768
rect 10332 24751 10334 24771
rect 10380 24751 10382 24771
rect 10428 24751 10430 24771
rect 10524 24751 10526 24771
rect 10527 24768 10541 24771
rect 10548 24771 17117 24775
rect 10548 24768 10565 24771
rect 10548 24751 10550 24768
rect 10620 24751 10622 24771
rect 10644 24751 10646 24771
rect 10716 24751 10718 24771
rect 10884 24751 10886 24771
rect 10956 24751 10958 24771
rect 11052 24751 11054 24771
rect 11100 24751 11102 24771
rect 11172 24751 11174 24771
rect 11220 24751 11222 24771
rect 11340 24751 11342 24771
rect 11436 24751 11438 24771
rect 11532 24751 11534 24771
rect 11628 24751 11630 24771
rect 11676 24751 11678 24771
rect 11724 24751 11726 24771
rect 11772 24751 11774 24771
rect 11796 24751 11798 24771
rect 11881 24766 11884 24771
rect 11892 24766 11894 24771
rect 11891 24752 11894 24766
rect 11988 24768 11990 24771
rect 11988 24751 11991 24768
rect 12060 24751 12062 24771
rect 12276 24751 12278 24771
rect 12324 24751 12326 24771
rect 12372 24751 12374 24771
rect 12420 24751 12422 24771
rect 12444 24751 12446 24771
rect 12468 24751 12470 24771
rect 12505 24766 12508 24771
rect 12516 24766 12518 24771
rect 12515 24752 12518 24766
rect 12540 24751 12542 24771
rect 12564 24751 12566 24771
rect 12660 24751 12662 24771
rect 12756 24751 12758 24771
rect 12828 24751 12830 24771
rect 12876 24751 12878 24771
rect 12972 24751 12974 24771
rect 13044 24751 13046 24771
rect 13068 24751 13070 24771
rect 13284 24751 13286 24771
rect 13332 24751 13334 24771
rect 13500 24751 13502 24771
rect 13572 24751 13574 24771
rect 13668 24751 13670 24771
rect 13716 24751 13718 24771
rect 13764 24751 13766 24771
rect 13860 24751 13862 24771
rect 13956 24751 13958 24771
rect 14004 24751 14006 24771
rect 14100 24751 14102 24771
rect 14940 24751 14942 24771
rect 15036 24751 15038 24771
rect 15276 24751 15278 24771
rect 15420 24751 15422 24771
rect 15564 24751 15566 24771
rect 15660 24751 15662 24771
rect 15708 24751 15710 24771
rect 15732 24751 15734 24771
rect 15756 24751 15758 24771
rect 15804 24751 15806 24771
rect 15828 24751 15830 24771
rect 15852 24751 15854 24771
rect 15948 24751 15950 24771
rect 15972 24751 15974 24771
rect 16044 24751 16046 24771
rect 16068 24751 16070 24771
rect 16164 24751 16166 24771
rect 16260 24751 16262 24771
rect 16332 24751 16334 24771
rect 16380 24751 16382 24771
rect 16476 24751 16478 24771
rect 16548 24751 16550 24771
rect 16572 24751 16574 24771
rect 16620 24751 16622 24771
rect 16668 24751 16670 24771
rect 16716 24751 16718 24771
rect 16764 24751 16766 24771
rect 16812 24751 16814 24771
rect 16884 24751 16886 24771
rect 16908 24751 16910 24771
rect 16980 24751 16982 24771
rect 17028 24751 17030 24771
rect 17103 24768 17117 24771
rect 17124 24771 23123 24775
rect 17124 24768 17141 24771
rect 17148 24768 17151 24771
rect 17124 24751 17126 24768
rect 17196 24751 17198 24771
rect 17220 24751 17222 24771
rect 17292 24751 17294 24771
rect 17316 24751 17318 24771
rect 17953 24766 17956 24771
rect 17963 24752 17966 24766
rect 17964 24751 17966 24752
rect 18060 24751 18063 24768
rect 18132 24751 18134 24771
rect 18228 24751 18230 24771
rect 18492 24751 18494 24771
rect 18540 24751 18542 24771
rect 18636 24751 18638 24771
rect 18732 24751 18734 24771
rect 18828 24751 18830 24771
rect 18924 24751 18926 24771
rect 18972 24751 18974 24771
rect 19020 24751 19022 24771
rect 19068 24751 19070 24771
rect 19140 24751 19142 24771
rect 19164 24751 19166 24771
rect 19236 24751 19238 24771
rect 19260 24751 19262 24771
rect 19788 24751 19790 24771
rect 19836 24751 19838 24771
rect 19860 24751 19862 24771
rect 19884 24751 19886 24771
rect 19956 24751 19958 24771
rect 19980 24751 19982 24771
rect 20004 24751 20006 24771
rect 20052 24751 20054 24771
rect 20076 24751 20078 24771
rect 20100 24751 20102 24771
rect 20172 24751 20174 24771
rect 20196 24751 20198 24771
rect 20292 24751 20294 24771
rect 20388 24751 20390 24771
rect 20412 24751 20414 24771
rect 20508 24751 20510 24771
rect 20532 24751 20534 24771
rect 20604 24751 20606 24771
rect 20628 24751 20630 24771
rect 20892 24751 20894 24771
rect 20964 24751 20966 24771
rect 20988 24751 20990 24771
rect 21108 24751 21110 24771
rect 21204 24751 21206 24771
rect 21300 24751 21302 24771
rect 21324 24751 21326 24771
rect 21444 24751 21446 24771
rect 21468 24751 21470 24771
rect 21564 24751 21566 24771
rect 21588 24751 21590 24771
rect 21684 24751 21686 24771
rect 21708 24751 21710 24771
rect 22068 24751 22070 24771
rect 22188 24751 22190 24771
rect 22212 24751 22214 24771
rect 22884 24751 22886 24771
rect 22980 24751 22982 24771
rect 23076 24752 23078 24771
rect 23089 24766 23092 24771
rect 23100 24766 23102 24771
rect 23099 24752 23102 24766
rect 22993 24751 23051 24752
rect 23065 24751 23099 24752
rect -11207 24747 18053 24751
rect -11207 24744 -11203 24747
rect -11196 24744 -11193 24747
rect -11100 24744 -11098 24747
rect -11100 24728 -11097 24744
rect -11111 24727 -11077 24728
rect -9900 24727 -9898 24747
rect -9732 24727 -9730 24747
rect -9636 24727 -9634 24747
rect -9540 24727 -9538 24747
rect -9444 24727 -9442 24747
rect -9348 24727 -9346 24747
rect -9228 24727 -9226 24747
rect -9108 24727 -9106 24747
rect -9012 24727 -9010 24747
rect -8916 24727 -8914 24747
rect -8628 24727 -8626 24747
rect -8532 24727 -8530 24747
rect -8436 24727 -8434 24747
rect -8340 24727 -8338 24747
rect -8289 24744 -8275 24747
rect -8268 24744 -8265 24747
rect -8124 24727 -8122 24747
rect -7764 24727 -7762 24747
rect -7524 24727 -7522 24747
rect -7356 24727 -7354 24747
rect -7308 24727 -7306 24747
rect -7140 24727 -7138 24747
rect -7044 24727 -7042 24747
rect -6948 24727 -6946 24747
rect -6852 24727 -6850 24747
rect -6732 24727 -6730 24747
rect -6516 24727 -6514 24747
rect -5892 24727 -5890 24747
rect -5436 24727 -5434 24747
rect -5340 24727 -5338 24747
rect -5196 24727 -5194 24747
rect -4716 24727 -4714 24747
rect -4500 24727 -4498 24747
rect -4404 24727 -4402 24747
rect -4308 24727 -4306 24747
rect -4164 24727 -4162 24747
rect -3876 24727 -3874 24747
rect -3540 24727 -3538 24747
rect -3468 24727 -3466 24747
rect -3324 24727 -3322 24747
rect -3108 24727 -3106 24747
rect -3012 24727 -3010 24747
rect -2964 24727 -2962 24747
rect -2916 24727 -2914 24747
rect -2868 24727 -2866 24747
rect -2820 24727 -2818 24747
rect -2772 24727 -2770 24747
rect -2676 24727 -2674 24747
rect -2364 24727 -2362 24747
rect -2316 24727 -2314 24747
rect -2076 24727 -2074 24747
rect -1980 24727 -1978 24747
rect -1812 24727 -1810 24747
rect -1572 24727 -1570 24747
rect -1476 24727 -1474 24747
rect -1356 24727 -1354 24747
rect -1260 24727 -1258 24747
rect -1236 24727 -1234 24747
rect -1140 24727 -1138 24747
rect -876 24727 -874 24747
rect -660 24727 -658 24747
rect -492 24727 -490 24747
rect -396 24727 -394 24747
rect -372 24727 -370 24747
rect -276 24727 -274 24747
rect -12 24727 -10 24747
rect 84 24727 86 24747
rect 156 24727 158 24747
rect 252 24727 254 24747
rect 348 24727 350 24747
rect 468 24727 470 24747
rect 492 24727 494 24747
rect 564 24727 566 24747
rect 588 24727 590 24747
rect 636 24727 638 24747
rect 660 24727 662 24747
rect 732 24727 734 24747
rect 948 24727 950 24747
rect 1044 24727 1046 24747
rect 1092 24727 1094 24747
rect 1140 24727 1142 24747
rect 1308 24727 1310 24747
rect 1356 24727 1358 24747
rect 1428 24727 1430 24747
rect 1692 24727 1694 24747
rect 1860 24727 1862 24747
rect 2079 24744 2093 24747
rect 2100 24744 2103 24747
rect 2148 24727 2150 24747
rect 2244 24727 2246 24747
rect 2460 24727 2462 24747
rect 2772 24727 2774 24747
rect 2868 24727 2870 24747
rect 2940 24727 2942 24747
rect 2988 24727 2990 24747
rect 3324 24727 3326 24747
rect 3396 24727 3398 24747
rect 3564 24727 3566 24747
rect 3660 24727 3662 24747
rect 3780 24727 3782 24747
rect 4092 24727 4094 24747
rect 4188 24727 4190 24747
rect 4308 24727 4310 24747
rect 4404 24727 4406 24747
rect 4500 24727 4502 24747
rect 4596 24727 4598 24747
rect 4692 24727 4694 24747
rect 4956 24727 4958 24747
rect 4980 24727 4982 24747
rect 4983 24744 4997 24747
rect 5052 24727 5054 24747
rect 5124 24727 5126 24747
rect 5220 24727 5222 24747
rect 5388 24727 5390 24747
rect 5484 24727 5486 24747
rect 5508 24727 5510 24747
rect 5532 24727 5534 24747
rect 5628 24727 5630 24747
rect 5652 24727 5654 24747
rect 5748 24727 5750 24747
rect 5796 24727 5798 24747
rect 5844 24727 5846 24747
rect 5892 24727 5894 24747
rect 6276 24727 6278 24747
rect 6372 24727 6374 24747
rect 6420 24727 6422 24747
rect 6492 24727 6494 24747
rect 6516 24727 6518 24747
rect 6588 24727 6590 24747
rect 6612 24727 6614 24747
rect 6684 24727 6686 24747
rect 6708 24727 6710 24747
rect 6780 24727 6782 24747
rect 6804 24727 6806 24747
rect 6900 24727 6902 24747
rect 6924 24727 6926 24747
rect 7020 24727 7022 24747
rect 7164 24727 7166 24747
rect 7236 24727 7238 24747
rect 7284 24727 7286 24747
rect 7380 24727 7382 24747
rect 7404 24727 7406 24747
rect 7476 24727 7478 24747
rect 7500 24727 7502 24747
rect 7572 24727 7574 24747
rect 7644 24727 7646 24747
rect 7668 24727 7670 24747
rect 7908 24727 7910 24747
rect 8124 24727 8126 24747
rect 8220 24727 8222 24747
rect 8652 24727 8654 24747
rect 8700 24727 8702 24747
rect 8748 24727 8750 24747
rect 8796 24727 8798 24747
rect 8844 24727 8846 24747
rect 8868 24727 8870 24747
rect 9516 24727 9518 24747
rect 9660 24727 9662 24747
rect 9684 24727 9686 24747
rect 9756 24727 9758 24747
rect 9780 24727 9782 24747
rect 9804 24727 9806 24747
rect 9852 24727 9854 24747
rect 9948 24727 9950 24747
rect 10044 24727 10046 24747
rect 10140 24727 10142 24747
rect 10167 24744 10181 24747
rect 10236 24727 10238 24747
rect 10263 24744 10277 24747
rect 10284 24744 10287 24747
rect 10332 24727 10334 24747
rect 10380 24727 10382 24747
rect 10428 24727 10430 24747
rect 10524 24727 10526 24747
rect 10548 24727 10550 24747
rect 10620 24727 10622 24747
rect 10644 24727 10646 24747
rect 10716 24727 10718 24747
rect 10884 24727 10886 24747
rect 10956 24727 10958 24747
rect 11052 24727 11054 24747
rect 11100 24727 11102 24747
rect 11172 24727 11174 24747
rect 11220 24727 11222 24747
rect 11340 24727 11342 24747
rect 11436 24727 11438 24747
rect 11532 24727 11534 24747
rect 11628 24727 11630 24747
rect 11676 24727 11678 24747
rect 11724 24727 11726 24747
rect 11772 24727 11774 24747
rect 11796 24727 11798 24747
rect 11967 24744 11981 24747
rect 11988 24744 11991 24747
rect 12060 24727 12062 24747
rect 12276 24727 12278 24747
rect 12324 24727 12326 24747
rect 12372 24727 12374 24747
rect 12420 24727 12422 24747
rect 12444 24727 12446 24747
rect 12468 24727 12470 24747
rect 12540 24727 12542 24747
rect 12564 24727 12566 24747
rect 12591 24744 12605 24747
rect 12660 24727 12662 24747
rect 12756 24727 12758 24747
rect 12828 24727 12830 24747
rect 12876 24727 12878 24747
rect 12972 24727 12974 24747
rect 13044 24727 13046 24747
rect 13068 24727 13070 24747
rect 13284 24727 13286 24747
rect 13332 24727 13334 24747
rect 13500 24727 13502 24747
rect 13572 24727 13574 24747
rect 13668 24727 13670 24747
rect 13716 24727 13718 24747
rect 13764 24727 13766 24747
rect 13860 24727 13862 24747
rect 13956 24727 13958 24747
rect 14004 24727 14006 24747
rect 14100 24727 14102 24747
rect 14940 24727 14942 24747
rect 15036 24727 15038 24747
rect 15276 24727 15278 24747
rect 15420 24727 15422 24747
rect 15564 24727 15566 24747
rect 15660 24727 15662 24747
rect 15708 24727 15710 24747
rect 15732 24727 15734 24747
rect 15756 24727 15758 24747
rect 15804 24727 15806 24747
rect 15828 24727 15830 24747
rect 15852 24727 15854 24747
rect 15948 24727 15950 24747
rect 15972 24727 15974 24747
rect 16044 24727 16046 24747
rect 16068 24727 16070 24747
rect 16164 24727 16166 24747
rect 16260 24727 16262 24747
rect 16332 24727 16334 24747
rect 16380 24727 16382 24747
rect 16476 24727 16478 24747
rect 16548 24727 16550 24747
rect 16572 24727 16574 24747
rect 16620 24727 16622 24747
rect 16668 24727 16670 24747
rect 16716 24727 16718 24747
rect 16764 24727 16766 24747
rect 16812 24727 16814 24747
rect 16884 24727 16886 24747
rect 16908 24727 16910 24747
rect 16980 24727 16982 24747
rect 17028 24727 17030 24747
rect 17124 24727 17126 24747
rect 17196 24727 17198 24747
rect 17220 24727 17222 24747
rect 17292 24727 17294 24747
rect 17316 24727 17318 24747
rect 17964 24727 17966 24747
rect 18039 24744 18053 24747
rect 18060 24747 23099 24751
rect 18060 24744 18077 24747
rect 18060 24727 18062 24744
rect 18132 24727 18134 24747
rect 18228 24727 18230 24747
rect 18492 24727 18494 24747
rect 18540 24727 18542 24747
rect 18636 24727 18638 24747
rect 18732 24727 18734 24747
rect 18828 24727 18830 24747
rect 18924 24727 18926 24747
rect 18972 24727 18974 24747
rect 19020 24727 19022 24747
rect 19068 24727 19070 24747
rect 19140 24727 19142 24747
rect 19164 24727 19166 24747
rect 19236 24727 19238 24747
rect 19260 24727 19262 24747
rect 19788 24727 19790 24747
rect 19836 24727 19838 24747
rect 19860 24727 19862 24747
rect 19884 24727 19886 24747
rect 19956 24727 19958 24747
rect 19980 24727 19982 24747
rect 20004 24727 20006 24747
rect 20052 24727 20054 24747
rect 20076 24727 20078 24747
rect 20100 24727 20102 24747
rect 20172 24727 20174 24747
rect 20196 24727 20198 24747
rect 20292 24727 20294 24747
rect 20388 24727 20390 24747
rect 20412 24727 20414 24747
rect 20508 24727 20510 24747
rect 20532 24727 20534 24747
rect 20604 24727 20606 24747
rect 20628 24727 20630 24747
rect 20892 24727 20894 24747
rect 20964 24727 20966 24747
rect 20988 24727 20990 24747
rect 21108 24727 21110 24747
rect 21204 24727 21206 24747
rect 21300 24727 21302 24747
rect 21324 24727 21326 24747
rect 21444 24727 21446 24747
rect 21468 24727 21470 24747
rect 21564 24727 21566 24747
rect 21588 24727 21590 24747
rect 21684 24727 21686 24747
rect 21708 24727 21710 24747
rect 22068 24727 22070 24747
rect 22188 24727 22190 24747
rect 22212 24727 22214 24747
rect 22884 24727 22886 24747
rect 22980 24728 22982 24747
rect 23065 24742 23068 24747
rect 23076 24742 23078 24747
rect 23075 24728 23078 24742
rect 23089 24734 23093 24742
rect 23079 24728 23089 24734
rect 22969 24727 23003 24728
rect -11111 24723 23003 24727
rect -11111 24720 -11107 24723
rect -11100 24720 -11097 24723
rect -10871 24703 -10837 24704
rect -9900 24703 -9898 24723
rect -9732 24703 -9730 24723
rect -9636 24703 -9634 24723
rect -9540 24703 -9538 24723
rect -9444 24703 -9442 24723
rect -9348 24703 -9346 24723
rect -9228 24703 -9226 24723
rect -9108 24703 -9106 24723
rect -9012 24703 -9010 24723
rect -8916 24703 -8914 24723
rect -8628 24703 -8626 24723
rect -8532 24703 -8530 24723
rect -8436 24703 -8434 24723
rect -8340 24703 -8338 24723
rect -8124 24703 -8122 24723
rect -7764 24703 -7762 24723
rect -7524 24703 -7522 24723
rect -7356 24703 -7354 24723
rect -7308 24703 -7306 24723
rect -7140 24703 -7138 24723
rect -7044 24703 -7042 24723
rect -6948 24703 -6946 24723
rect -6852 24703 -6850 24723
rect -6732 24703 -6730 24723
rect -6516 24703 -6514 24723
rect -5892 24703 -5890 24723
rect -5436 24703 -5434 24723
rect -5340 24703 -5338 24723
rect -5196 24703 -5194 24723
rect -4716 24703 -4714 24723
rect -4500 24703 -4498 24723
rect -4404 24703 -4402 24723
rect -4308 24703 -4306 24723
rect -4164 24703 -4162 24723
rect -3876 24703 -3874 24723
rect -3540 24703 -3538 24723
rect -3468 24703 -3466 24723
rect -3324 24703 -3322 24723
rect -3108 24703 -3106 24723
rect -3012 24703 -3010 24723
rect -2964 24703 -2962 24723
rect -2916 24703 -2914 24723
rect -2868 24703 -2866 24723
rect -2820 24703 -2818 24723
rect -2772 24703 -2770 24723
rect -2676 24703 -2674 24723
rect -2364 24703 -2362 24723
rect -2316 24703 -2314 24723
rect -2076 24703 -2074 24723
rect -1980 24703 -1978 24723
rect -1812 24703 -1810 24723
rect -1572 24703 -1570 24723
rect -1476 24703 -1474 24723
rect -1356 24703 -1354 24723
rect -1260 24703 -1258 24723
rect -1236 24703 -1234 24723
rect -1140 24703 -1138 24723
rect -876 24703 -874 24723
rect -660 24703 -658 24723
rect -492 24703 -490 24723
rect -396 24703 -394 24723
rect -372 24703 -370 24723
rect -276 24703 -274 24723
rect -12 24703 -10 24723
rect 84 24703 86 24723
rect 156 24703 158 24723
rect 252 24703 254 24723
rect 348 24703 350 24723
rect 468 24703 470 24723
rect 492 24703 494 24723
rect 564 24703 566 24723
rect 588 24703 590 24723
rect 636 24703 638 24723
rect 660 24703 662 24723
rect 732 24703 734 24723
rect 948 24703 950 24723
rect 1044 24703 1046 24723
rect 1092 24703 1094 24723
rect 1140 24703 1142 24723
rect 1308 24703 1310 24723
rect 1356 24703 1358 24723
rect 1428 24703 1430 24723
rect 1692 24703 1694 24723
rect 1860 24703 1862 24723
rect 2148 24703 2150 24723
rect 2244 24703 2246 24723
rect 2460 24703 2462 24723
rect 2772 24703 2774 24723
rect 2868 24703 2870 24723
rect 2940 24703 2942 24723
rect 2988 24703 2990 24723
rect 3324 24703 3326 24723
rect 3396 24703 3398 24723
rect 3564 24703 3566 24723
rect 3660 24703 3662 24723
rect 3780 24703 3782 24723
rect 4092 24703 4094 24723
rect 4188 24703 4190 24723
rect 4308 24703 4310 24723
rect 4404 24703 4406 24723
rect 4500 24703 4502 24723
rect 4596 24703 4598 24723
rect 4692 24703 4694 24723
rect 4956 24703 4958 24723
rect 4980 24703 4982 24723
rect 5052 24703 5054 24723
rect 5124 24703 5126 24723
rect 5220 24703 5222 24723
rect 5388 24703 5390 24723
rect 5484 24703 5486 24723
rect 5508 24703 5510 24723
rect 5532 24703 5534 24723
rect 5628 24703 5630 24723
rect 5652 24703 5654 24723
rect 5748 24703 5750 24723
rect 5796 24703 5798 24723
rect 5844 24703 5846 24723
rect 5892 24703 5894 24723
rect 6276 24703 6278 24723
rect 6372 24703 6374 24723
rect 6420 24703 6422 24723
rect 6492 24703 6494 24723
rect 6516 24703 6518 24723
rect 6529 24703 6587 24704
rect 6588 24703 6590 24723
rect 6612 24703 6614 24723
rect 6684 24703 6686 24723
rect 6708 24703 6710 24723
rect 6780 24703 6782 24723
rect 6804 24703 6806 24723
rect 6900 24703 6902 24723
rect 6924 24703 6926 24723
rect 7020 24703 7022 24723
rect 7164 24703 7166 24723
rect 7236 24703 7238 24723
rect 7284 24703 7286 24723
rect 7380 24703 7382 24723
rect 7404 24703 7406 24723
rect 7476 24703 7478 24723
rect 7500 24703 7502 24723
rect 7572 24703 7574 24723
rect 7644 24703 7646 24723
rect 7668 24703 7670 24723
rect 7908 24703 7910 24723
rect 8124 24703 8126 24723
rect 8220 24703 8222 24723
rect 8652 24703 8654 24723
rect 8700 24703 8702 24723
rect 8748 24703 8750 24723
rect 8796 24703 8798 24723
rect 8844 24703 8846 24723
rect 8868 24703 8870 24723
rect 9516 24703 9518 24723
rect 9660 24703 9662 24723
rect 9684 24703 9686 24723
rect 9756 24703 9758 24723
rect 9780 24703 9782 24723
rect 9804 24703 9806 24723
rect 9852 24703 9854 24723
rect 9948 24703 9950 24723
rect 10044 24703 10046 24723
rect 10140 24703 10142 24723
rect 10236 24703 10238 24723
rect 10332 24703 10334 24723
rect 10380 24703 10382 24723
rect 10428 24703 10430 24723
rect 10524 24703 10526 24723
rect 10548 24703 10550 24723
rect 10620 24703 10622 24723
rect 10644 24703 10646 24723
rect 10716 24703 10718 24723
rect 10884 24703 10886 24723
rect 10956 24703 10958 24723
rect 11052 24703 11054 24723
rect 11100 24703 11102 24723
rect 11172 24703 11174 24723
rect 11220 24703 11222 24723
rect 11340 24703 11342 24723
rect 11436 24703 11438 24723
rect 11532 24704 11534 24723
rect 11497 24703 11555 24704
rect 11628 24703 11630 24723
rect 11676 24703 11678 24723
rect 11724 24703 11726 24723
rect 11772 24703 11774 24723
rect 11796 24703 11798 24723
rect 12060 24703 12062 24723
rect 12276 24703 12278 24723
rect 12324 24703 12326 24723
rect 12372 24703 12374 24723
rect 12420 24703 12422 24723
rect 12444 24703 12446 24723
rect 12468 24703 12470 24723
rect 12540 24703 12542 24723
rect 12564 24703 12566 24723
rect 12660 24703 12662 24723
rect 12756 24703 12758 24723
rect 12828 24703 12830 24723
rect 12876 24703 12878 24723
rect 12972 24703 12974 24723
rect 13044 24703 13046 24723
rect 13068 24703 13070 24723
rect 13284 24703 13286 24723
rect 13332 24703 13334 24723
rect 13500 24703 13502 24723
rect 13572 24703 13574 24723
rect 13668 24703 13670 24723
rect 13716 24703 13718 24723
rect 13764 24703 13766 24723
rect 13860 24703 13862 24723
rect 13956 24703 13958 24723
rect 14004 24703 14006 24723
rect 14100 24703 14102 24723
rect 14940 24703 14942 24723
rect 15036 24703 15038 24723
rect 15276 24703 15278 24723
rect 15420 24703 15422 24723
rect 15564 24703 15566 24723
rect 15660 24703 15662 24723
rect 15708 24703 15710 24723
rect 15732 24703 15734 24723
rect 15756 24703 15758 24723
rect 15804 24703 15806 24723
rect 15828 24703 15830 24723
rect 15852 24703 15854 24723
rect 15948 24703 15950 24723
rect 15972 24703 15974 24723
rect 16044 24703 16046 24723
rect 16068 24703 16070 24723
rect 16164 24703 16166 24723
rect 16260 24703 16262 24723
rect 16332 24703 16334 24723
rect 16380 24703 16382 24723
rect 16476 24703 16478 24723
rect 16548 24703 16550 24723
rect 16572 24703 16574 24723
rect 16620 24704 16622 24723
rect 16585 24703 16643 24704
rect 16668 24703 16670 24723
rect 16716 24703 16718 24723
rect 16764 24703 16766 24723
rect 16812 24703 16814 24723
rect 16884 24703 16886 24723
rect 16908 24703 16910 24723
rect 16980 24703 16982 24723
rect 17028 24703 17030 24723
rect 17124 24703 17126 24723
rect 17196 24703 17198 24723
rect 17220 24703 17222 24723
rect 17292 24703 17294 24723
rect 17316 24703 17318 24723
rect 17964 24703 17966 24723
rect 18060 24703 18062 24723
rect 18132 24703 18134 24723
rect 18228 24703 18230 24723
rect 18492 24703 18494 24723
rect 18540 24703 18542 24723
rect 18636 24703 18638 24723
rect 18732 24703 18734 24723
rect 18828 24703 18830 24723
rect 18924 24703 18926 24723
rect 18972 24703 18974 24723
rect 19020 24703 19022 24723
rect 19068 24703 19070 24723
rect 19140 24703 19142 24723
rect 19164 24703 19166 24723
rect 19236 24703 19238 24723
rect 19260 24703 19262 24723
rect 19788 24703 19790 24723
rect 19836 24703 19838 24723
rect 19860 24703 19862 24723
rect 19884 24703 19886 24723
rect 19956 24703 19958 24723
rect 19980 24703 19982 24723
rect 20004 24703 20006 24723
rect 20052 24703 20054 24723
rect 20076 24703 20078 24723
rect 20100 24703 20102 24723
rect 20172 24703 20174 24723
rect 20196 24703 20198 24723
rect 20292 24703 20294 24723
rect 20388 24703 20390 24723
rect 20412 24703 20414 24723
rect 20508 24703 20510 24723
rect 20532 24703 20534 24723
rect 20604 24703 20606 24723
rect 20628 24703 20630 24723
rect 20892 24703 20894 24723
rect 20964 24703 20966 24723
rect 20988 24703 20990 24723
rect 21108 24703 21110 24723
rect 21204 24703 21206 24723
rect 21300 24703 21302 24723
rect 21324 24703 21326 24723
rect 21444 24703 21446 24723
rect 21468 24703 21470 24723
rect 21564 24703 21566 24723
rect 21588 24703 21590 24723
rect 21684 24703 21686 24723
rect 21708 24703 21710 24723
rect 22068 24703 22070 24723
rect 22188 24703 22190 24723
rect 22212 24703 22214 24723
rect 22884 24704 22886 24723
rect 22969 24718 22972 24723
rect 22980 24718 22982 24723
rect 22979 24704 22982 24718
rect 22777 24703 22811 24704
rect -10871 24699 22811 24703
rect 22873 24703 22907 24704
rect 22945 24703 22979 24704
rect 22873 24699 22979 24703
rect -10751 24679 -10717 24680
rect -9900 24679 -9898 24699
rect -9732 24679 -9730 24699
rect -9636 24679 -9634 24699
rect -9540 24679 -9538 24699
rect -9444 24679 -9442 24699
rect -9348 24679 -9346 24699
rect -9228 24679 -9226 24699
rect -9108 24679 -9106 24699
rect -9012 24679 -9010 24699
rect -8916 24679 -8914 24699
rect -8628 24679 -8626 24699
rect -8532 24679 -8530 24699
rect -8436 24679 -8434 24699
rect -8340 24679 -8338 24699
rect -8124 24679 -8122 24699
rect -7764 24679 -7762 24699
rect -7524 24679 -7522 24699
rect -7356 24679 -7354 24699
rect -7308 24679 -7306 24699
rect -7140 24679 -7138 24699
rect -7044 24679 -7042 24699
rect -6948 24679 -6946 24699
rect -6852 24679 -6850 24699
rect -6732 24679 -6730 24699
rect -6516 24679 -6514 24699
rect -5892 24679 -5890 24699
rect -5436 24679 -5434 24699
rect -5340 24679 -5338 24699
rect -5196 24679 -5194 24699
rect -4716 24679 -4714 24699
rect -4500 24679 -4498 24699
rect -4404 24679 -4402 24699
rect -4308 24679 -4306 24699
rect -4164 24679 -4162 24699
rect -3876 24679 -3874 24699
rect -3540 24679 -3538 24699
rect -3468 24679 -3466 24699
rect -3324 24679 -3322 24699
rect -3108 24679 -3106 24699
rect -3012 24679 -3010 24699
rect -2964 24679 -2962 24699
rect -2916 24679 -2914 24699
rect -2868 24679 -2866 24699
rect -2820 24679 -2818 24699
rect -2772 24679 -2770 24699
rect -2676 24679 -2674 24699
rect -2364 24679 -2362 24699
rect -2351 24679 -2317 24680
rect -2316 24679 -2314 24699
rect -2183 24679 -2149 24680
rect -2076 24679 -2074 24699
rect -1980 24679 -1978 24699
rect -1812 24679 -1810 24699
rect -1572 24679 -1570 24699
rect -1476 24679 -1474 24699
rect -1356 24679 -1354 24699
rect -1260 24679 -1258 24699
rect -1236 24679 -1234 24699
rect -1140 24679 -1138 24699
rect -876 24679 -874 24699
rect -660 24679 -658 24699
rect -492 24679 -490 24699
rect -396 24679 -394 24699
rect -372 24679 -370 24699
rect -276 24679 -274 24699
rect -12 24679 -10 24699
rect 84 24679 86 24699
rect 156 24679 158 24699
rect 252 24679 254 24699
rect 348 24679 350 24699
rect 468 24679 470 24699
rect 492 24679 494 24699
rect 564 24679 566 24699
rect 588 24679 590 24699
rect 636 24679 638 24699
rect 660 24679 662 24699
rect 732 24679 734 24699
rect 948 24679 950 24699
rect 1044 24679 1046 24699
rect 1092 24679 1094 24699
rect 1140 24679 1142 24699
rect 1308 24679 1310 24699
rect 1356 24679 1358 24699
rect 1428 24679 1430 24699
rect 1692 24679 1694 24699
rect 1860 24679 1862 24699
rect 2148 24679 2150 24699
rect 2244 24679 2246 24699
rect 2460 24679 2462 24699
rect 2772 24679 2774 24699
rect 2868 24679 2870 24699
rect 2940 24679 2942 24699
rect 2988 24679 2990 24699
rect 3324 24679 3326 24699
rect 3396 24679 3398 24699
rect 3564 24679 3566 24699
rect 3660 24679 3662 24699
rect 3780 24679 3782 24699
rect 4092 24679 4094 24699
rect 4188 24679 4190 24699
rect 4308 24679 4310 24699
rect 4404 24679 4406 24699
rect 4500 24679 4502 24699
rect 4596 24679 4598 24699
rect 4692 24679 4694 24699
rect 4956 24679 4958 24699
rect 4980 24679 4982 24699
rect 5052 24679 5054 24699
rect 5124 24679 5126 24699
rect 5220 24679 5222 24699
rect 5388 24679 5390 24699
rect 5484 24679 5486 24699
rect 5508 24679 5510 24699
rect 5532 24679 5534 24699
rect 5628 24679 5630 24699
rect 5652 24679 5654 24699
rect 5748 24679 5750 24699
rect 5796 24679 5798 24699
rect 5844 24679 5846 24699
rect 5892 24679 5894 24699
rect 6276 24679 6278 24699
rect 6372 24679 6374 24699
rect 6420 24679 6422 24699
rect 6492 24679 6494 24699
rect 6516 24679 6518 24699
rect 6588 24679 6590 24699
rect 6612 24679 6614 24699
rect 6636 24679 6639 24696
rect 6684 24679 6686 24699
rect 6708 24679 6710 24699
rect 6780 24679 6782 24699
rect 6804 24679 6806 24699
rect 6900 24679 6902 24699
rect 6924 24679 6926 24699
rect 7020 24679 7022 24699
rect 7164 24679 7166 24699
rect 7236 24679 7238 24699
rect 7284 24679 7286 24699
rect 7380 24679 7382 24699
rect 7404 24679 7406 24699
rect 7476 24679 7478 24699
rect 7500 24679 7502 24699
rect 7572 24679 7574 24699
rect 7644 24679 7646 24699
rect 7668 24679 7670 24699
rect 7908 24679 7910 24699
rect 8124 24679 8126 24699
rect 8220 24679 8222 24699
rect 8652 24679 8654 24699
rect 8700 24679 8702 24699
rect 8748 24679 8750 24699
rect 8796 24679 8798 24699
rect 8844 24679 8846 24699
rect 8868 24679 8870 24699
rect 9516 24679 9518 24699
rect 9660 24679 9662 24699
rect 9684 24679 9686 24699
rect 9756 24679 9758 24699
rect 9780 24679 9782 24699
rect 9804 24679 9806 24699
rect 9852 24679 9854 24699
rect 9948 24679 9950 24699
rect 10044 24679 10046 24699
rect 10140 24679 10142 24699
rect 10236 24679 10238 24699
rect 10332 24679 10334 24699
rect 10380 24679 10382 24699
rect 10428 24679 10430 24699
rect 10524 24679 10526 24699
rect 10548 24679 10550 24699
rect 10620 24679 10622 24699
rect 10644 24679 10646 24699
rect 10716 24679 10718 24699
rect 10884 24679 10886 24699
rect 10956 24679 10958 24699
rect 11052 24679 11054 24699
rect 11100 24679 11102 24699
rect 11172 24679 11174 24699
rect 11220 24679 11222 24699
rect 11340 24679 11342 24699
rect 11436 24679 11438 24699
rect 11521 24694 11524 24699
rect 11532 24694 11534 24699
rect 11531 24680 11534 24694
rect 11628 24696 11630 24699
rect 11628 24679 11631 24696
rect 11676 24679 11678 24699
rect 11724 24679 11726 24699
rect 11772 24679 11774 24699
rect 11796 24679 11798 24699
rect 12060 24679 12062 24699
rect 12276 24679 12278 24699
rect 12324 24679 12326 24699
rect 12372 24679 12374 24699
rect 12420 24679 12422 24699
rect 12444 24679 12446 24699
rect 12468 24679 12470 24699
rect 12540 24679 12542 24699
rect 12564 24679 12566 24699
rect 12660 24679 12662 24699
rect 12756 24679 12758 24699
rect 12828 24679 12830 24699
rect 12876 24679 12878 24699
rect 12972 24679 12974 24699
rect 13044 24679 13046 24699
rect 13068 24679 13070 24699
rect 13284 24679 13286 24699
rect 13332 24679 13334 24699
rect 13500 24679 13502 24699
rect 13572 24679 13574 24699
rect 13668 24679 13670 24699
rect 13716 24679 13718 24699
rect 13764 24679 13766 24699
rect 13860 24679 13862 24699
rect 13956 24679 13958 24699
rect 14004 24679 14006 24699
rect 14100 24679 14102 24699
rect 14940 24679 14942 24699
rect 15036 24679 15038 24699
rect 15276 24679 15278 24699
rect 15420 24679 15422 24699
rect 15564 24679 15566 24699
rect 15660 24679 15662 24699
rect 15708 24679 15710 24699
rect 15732 24679 15734 24699
rect 15756 24679 15758 24699
rect 15804 24679 15806 24699
rect 15828 24679 15830 24699
rect 15852 24679 15854 24699
rect 15948 24679 15950 24699
rect 15972 24679 15974 24699
rect 16044 24679 16046 24699
rect 16068 24679 16070 24699
rect 16164 24679 16166 24699
rect 16260 24679 16262 24699
rect 16332 24679 16334 24699
rect 16380 24679 16382 24699
rect 16476 24679 16478 24699
rect 16548 24679 16550 24699
rect 16572 24679 16574 24699
rect 16609 24694 16612 24699
rect 16620 24694 16622 24699
rect 16619 24680 16622 24694
rect 16668 24679 16670 24699
rect 16716 24696 16718 24699
rect 16716 24679 16719 24696
rect 16764 24679 16766 24699
rect 16812 24679 16814 24699
rect 16884 24679 16886 24699
rect 16908 24679 16910 24699
rect 16980 24679 16982 24699
rect 17028 24679 17030 24699
rect 17124 24679 17126 24699
rect 17196 24679 17198 24699
rect 17220 24679 17222 24699
rect 17292 24679 17294 24699
rect 17316 24679 17318 24699
rect 17964 24679 17966 24699
rect 18060 24679 18062 24699
rect 18132 24679 18134 24699
rect 18228 24679 18230 24699
rect 18492 24679 18494 24699
rect 18540 24679 18542 24699
rect 18636 24679 18638 24699
rect 18732 24679 18734 24699
rect 18828 24679 18830 24699
rect 18924 24679 18926 24699
rect 18972 24679 18974 24699
rect 19020 24679 19022 24699
rect 19068 24679 19070 24699
rect 19140 24679 19142 24699
rect 19164 24679 19166 24699
rect 19236 24679 19238 24699
rect 19260 24679 19262 24699
rect 19788 24679 19790 24699
rect 19836 24679 19838 24699
rect 19860 24679 19862 24699
rect 19884 24679 19886 24699
rect 19956 24679 19958 24699
rect 19980 24679 19982 24699
rect 20004 24679 20006 24699
rect 20052 24679 20054 24699
rect 20076 24679 20078 24699
rect 20100 24679 20102 24699
rect 20172 24679 20174 24699
rect 20196 24679 20198 24699
rect 20292 24679 20294 24699
rect 20388 24679 20390 24699
rect 20412 24679 20414 24699
rect 20508 24679 20510 24699
rect 20532 24679 20534 24699
rect 20604 24679 20606 24699
rect 20628 24679 20630 24699
rect 20892 24679 20894 24699
rect 20964 24679 20966 24699
rect 20988 24679 20990 24699
rect 21108 24679 21110 24699
rect 21204 24679 21206 24699
rect 21300 24679 21302 24699
rect 21324 24679 21326 24699
rect 21444 24679 21446 24699
rect 21468 24679 21470 24699
rect 21564 24679 21566 24699
rect 21588 24679 21590 24699
rect 21684 24679 21686 24699
rect 21708 24679 21710 24699
rect 22068 24679 22070 24699
rect 22188 24679 22190 24699
rect 22212 24679 22214 24699
rect 22873 24694 22876 24699
rect 22884 24696 22886 24699
rect 22884 24694 22887 24696
rect 22883 24680 22887 24694
rect 22969 24686 22973 24694
rect 22959 24680 22969 24686
rect 22369 24679 22403 24680
rect -10751 24675 6629 24679
rect -10535 24655 -10501 24656
rect -9900 24655 -9898 24675
rect -9732 24655 -9730 24675
rect -9636 24655 -9634 24675
rect -9540 24655 -9538 24675
rect -9444 24655 -9442 24675
rect -9348 24655 -9346 24675
rect -9228 24655 -9226 24675
rect -9108 24655 -9106 24675
rect -9012 24655 -9010 24675
rect -8916 24655 -8914 24675
rect -8628 24655 -8626 24675
rect -8532 24655 -8530 24675
rect -8436 24655 -8434 24675
rect -8340 24655 -8338 24675
rect -8124 24655 -8122 24675
rect -7943 24655 -7909 24656
rect -7764 24655 -7762 24675
rect -7524 24655 -7522 24675
rect -7356 24655 -7354 24675
rect -7308 24655 -7306 24675
rect -7140 24655 -7138 24675
rect -7044 24656 -7042 24675
rect -7055 24655 -7021 24656
rect -6948 24655 -6946 24675
rect -6852 24655 -6850 24675
rect -6791 24655 -6757 24656
rect -6732 24655 -6730 24675
rect -6516 24655 -6514 24675
rect -5892 24655 -5890 24675
rect -5436 24655 -5434 24675
rect -5340 24655 -5338 24675
rect -5196 24655 -5194 24675
rect -4716 24655 -4714 24675
rect -4500 24655 -4498 24675
rect -4404 24655 -4402 24675
rect -4308 24655 -4306 24675
rect -4164 24655 -4162 24675
rect -3876 24655 -3874 24675
rect -3540 24655 -3538 24675
rect -3468 24655 -3466 24675
rect -3324 24655 -3322 24675
rect -3108 24655 -3106 24675
rect -3012 24655 -3010 24675
rect -2964 24655 -2962 24675
rect -2916 24655 -2914 24675
rect -2868 24655 -2866 24675
rect -2820 24655 -2818 24675
rect -2772 24655 -2770 24675
rect -2676 24655 -2674 24675
rect -2364 24655 -2362 24675
rect -2316 24655 -2314 24675
rect -2076 24672 -2074 24675
rect -2076 24655 -2073 24672
rect -1980 24655 -1978 24675
rect -1812 24655 -1810 24675
rect -1572 24655 -1570 24675
rect -1476 24655 -1474 24675
rect -1356 24655 -1354 24675
rect -1260 24655 -1258 24675
rect -1236 24655 -1234 24675
rect -1140 24655 -1138 24675
rect -876 24655 -874 24675
rect -660 24655 -658 24675
rect -492 24655 -490 24675
rect -396 24655 -394 24675
rect -372 24656 -370 24675
rect -383 24655 -349 24656
rect -276 24655 -274 24675
rect -12 24655 -10 24675
rect 84 24655 86 24675
rect 156 24655 158 24675
rect 252 24655 254 24675
rect 348 24655 350 24675
rect 468 24655 470 24675
rect 492 24655 494 24675
rect 564 24655 566 24675
rect 588 24655 590 24675
rect 636 24655 638 24675
rect 660 24655 662 24675
rect 732 24655 734 24675
rect 948 24655 950 24675
rect 1044 24655 1046 24675
rect 1092 24655 1094 24675
rect 1140 24655 1142 24675
rect 1308 24655 1310 24675
rect 1356 24655 1358 24675
rect 1428 24655 1430 24675
rect 1692 24655 1694 24675
rect 1860 24655 1862 24675
rect 2148 24655 2150 24675
rect 2244 24655 2246 24675
rect 2460 24655 2462 24675
rect 2772 24655 2774 24675
rect 2868 24655 2870 24675
rect 2940 24655 2942 24675
rect 2988 24655 2990 24675
rect 3324 24655 3326 24675
rect 3396 24655 3398 24675
rect 3564 24655 3566 24675
rect 3660 24655 3662 24675
rect 3780 24655 3782 24675
rect 4092 24655 4094 24675
rect 4188 24655 4190 24675
rect 4308 24655 4310 24675
rect 4404 24655 4406 24675
rect 4500 24655 4502 24675
rect 4596 24655 4598 24675
rect 4692 24655 4694 24675
rect 4956 24656 4958 24675
rect 4921 24655 4979 24656
rect 4980 24655 4982 24675
rect 5052 24655 5054 24675
rect 5124 24655 5126 24675
rect 5220 24655 5222 24675
rect 5388 24655 5390 24675
rect 5484 24655 5486 24675
rect 5508 24655 5510 24675
rect 5532 24655 5534 24675
rect 5628 24655 5630 24675
rect 5652 24655 5654 24675
rect 5748 24655 5750 24675
rect 5796 24655 5798 24675
rect 5844 24655 5846 24675
rect 5892 24655 5894 24675
rect 6276 24655 6278 24675
rect 6372 24655 6374 24675
rect 6420 24655 6422 24675
rect 6492 24655 6494 24675
rect 6516 24655 6518 24675
rect 6588 24655 6590 24675
rect 6612 24655 6614 24675
rect 6615 24672 6629 24675
rect 6636 24675 11597 24679
rect 6636 24672 6653 24675
rect 6636 24655 6638 24672
rect 6684 24655 6686 24675
rect 6708 24655 6710 24675
rect 6780 24655 6782 24675
rect 6804 24655 6806 24675
rect 6900 24655 6902 24675
rect 6924 24655 6926 24675
rect 7020 24655 7022 24675
rect 7164 24655 7166 24675
rect 7236 24655 7238 24675
rect 7284 24655 7286 24675
rect 7380 24655 7382 24675
rect 7404 24655 7406 24675
rect 7476 24655 7478 24675
rect 7500 24655 7502 24675
rect 7572 24655 7574 24675
rect 7644 24655 7646 24675
rect 7668 24655 7670 24675
rect 7908 24655 7910 24675
rect 8124 24655 8126 24675
rect 8220 24655 8222 24675
rect 8652 24655 8654 24675
rect 8700 24655 8702 24675
rect 8748 24655 8750 24675
rect 8796 24655 8798 24675
rect 8844 24655 8846 24675
rect 8868 24655 8870 24675
rect 9516 24655 9518 24675
rect 9660 24655 9662 24675
rect 9684 24655 9686 24675
rect 9756 24655 9758 24675
rect 9780 24655 9782 24675
rect 9804 24655 9806 24675
rect 9852 24655 9854 24675
rect 9948 24655 9950 24675
rect 10044 24655 10046 24675
rect 10140 24655 10142 24675
rect 10236 24655 10238 24675
rect 10332 24655 10334 24675
rect 10380 24655 10382 24675
rect 10428 24655 10430 24675
rect 10524 24655 10526 24675
rect 10548 24655 10550 24675
rect 10620 24655 10622 24675
rect 10644 24655 10646 24675
rect 10716 24655 10718 24675
rect 10884 24655 10886 24675
rect 10956 24655 10958 24675
rect 11052 24655 11054 24675
rect 11100 24655 11102 24675
rect 11172 24655 11174 24675
rect 11220 24655 11222 24675
rect 11340 24655 11342 24675
rect 11436 24655 11438 24675
rect 11583 24672 11597 24675
rect 11607 24675 16685 24679
rect 11607 24672 11621 24675
rect 11628 24672 11631 24675
rect 11676 24655 11678 24675
rect 11724 24655 11726 24675
rect 11772 24655 11774 24675
rect 11796 24655 11798 24675
rect 12060 24655 12062 24675
rect 12276 24655 12278 24675
rect 12324 24655 12326 24675
rect 12372 24655 12374 24675
rect 12420 24655 12422 24675
rect 12444 24655 12446 24675
rect 12468 24655 12470 24675
rect 12540 24655 12542 24675
rect 12564 24655 12566 24675
rect 12660 24655 12662 24675
rect 12756 24655 12758 24675
rect 12828 24655 12830 24675
rect 12876 24655 12878 24675
rect 12972 24655 12974 24675
rect 13044 24655 13046 24675
rect 13068 24655 13070 24675
rect 13284 24655 13286 24675
rect 13332 24655 13334 24675
rect 13500 24655 13502 24675
rect 13572 24655 13574 24675
rect 13668 24655 13670 24675
rect 13716 24655 13718 24675
rect 13764 24655 13766 24675
rect 13860 24655 13862 24675
rect 13956 24655 13958 24675
rect 14004 24655 14006 24675
rect 14100 24655 14102 24675
rect 14940 24655 14942 24675
rect 15036 24655 15038 24675
rect 15276 24655 15278 24675
rect 15420 24655 15422 24675
rect 15564 24655 15566 24675
rect 15660 24655 15662 24675
rect 15708 24655 15710 24675
rect 15732 24655 15734 24675
rect 15756 24655 15758 24675
rect 15804 24655 15806 24675
rect 15828 24655 15830 24675
rect 15852 24655 15854 24675
rect 15948 24655 15950 24675
rect 15972 24655 15974 24675
rect 16044 24655 16046 24675
rect 16068 24655 16070 24675
rect 16164 24655 16166 24675
rect 16260 24655 16262 24675
rect 16332 24655 16334 24675
rect 16380 24655 16382 24675
rect 16476 24655 16478 24675
rect 16548 24655 16550 24675
rect 16572 24655 16574 24675
rect 16668 24655 16670 24675
rect 16671 24672 16685 24675
rect 16695 24675 22403 24679
rect 16695 24672 16709 24675
rect 16716 24672 16719 24675
rect 16764 24655 16766 24675
rect 16812 24655 16814 24675
rect 16884 24655 16886 24675
rect 16908 24655 16910 24675
rect 16980 24655 16982 24675
rect 17028 24655 17030 24675
rect 17124 24655 17126 24675
rect 17196 24655 17198 24675
rect 17220 24655 17222 24675
rect 17292 24655 17294 24675
rect 17316 24655 17318 24675
rect 17964 24655 17966 24675
rect 18060 24655 18062 24675
rect 18132 24655 18134 24675
rect 18228 24655 18230 24675
rect 18492 24655 18494 24675
rect 18540 24655 18542 24675
rect 18636 24655 18638 24675
rect 18732 24655 18734 24675
rect 18828 24655 18830 24675
rect 18924 24655 18926 24675
rect 18972 24655 18974 24675
rect 19020 24655 19022 24675
rect 19068 24655 19070 24675
rect 19140 24655 19142 24675
rect 19164 24655 19166 24675
rect 19236 24655 19238 24675
rect 19260 24655 19262 24675
rect 19788 24655 19790 24675
rect 19836 24655 19838 24675
rect 19860 24655 19862 24675
rect 19884 24655 19886 24675
rect 19956 24655 19958 24675
rect 19980 24655 19982 24675
rect 20004 24655 20006 24675
rect 20052 24655 20054 24675
rect 20076 24655 20078 24675
rect 20100 24655 20102 24675
rect 20172 24655 20174 24675
rect 20196 24655 20198 24675
rect 20292 24655 20294 24675
rect 20388 24655 20390 24675
rect 20412 24655 20414 24675
rect 20508 24655 20510 24675
rect 20532 24655 20534 24675
rect 20604 24655 20606 24675
rect 20628 24655 20630 24675
rect 20892 24655 20894 24675
rect 20964 24655 20966 24675
rect 20988 24655 20990 24675
rect 21108 24655 21110 24675
rect 21204 24655 21206 24675
rect 21300 24655 21302 24675
rect 21324 24655 21326 24675
rect 21444 24655 21446 24675
rect 21468 24655 21470 24675
rect 21564 24655 21566 24675
rect 21588 24655 21590 24675
rect 21684 24655 21686 24675
rect 21708 24655 21710 24675
rect 22068 24655 22070 24675
rect 22188 24655 22190 24675
rect 22212 24655 22214 24675
rect 22225 24655 22259 24656
rect -10535 24651 22259 24655
rect -9900 24631 -9898 24651
rect -9732 24631 -9730 24651
rect -9636 24631 -9634 24651
rect -9540 24631 -9538 24651
rect -9444 24631 -9442 24651
rect -9348 24631 -9346 24651
rect -9228 24631 -9226 24651
rect -9108 24631 -9106 24651
rect -9012 24631 -9010 24651
rect -8916 24631 -8914 24651
rect -8628 24631 -8626 24651
rect -8532 24631 -8530 24651
rect -8436 24631 -8434 24651
rect -8340 24631 -8338 24651
rect -8124 24631 -8122 24651
rect -7764 24631 -7762 24651
rect -7524 24631 -7522 24651
rect -7356 24631 -7354 24651
rect -7308 24631 -7306 24651
rect -7140 24631 -7138 24651
rect -7055 24646 -7052 24651
rect -7044 24646 -7042 24651
rect -7045 24632 -7042 24646
rect -6948 24648 -6946 24651
rect -6948 24631 -6945 24648
rect -6852 24631 -6850 24651
rect -6732 24631 -6730 24651
rect -6516 24631 -6514 24651
rect -5892 24631 -5890 24651
rect -5436 24631 -5434 24651
rect -5340 24631 -5338 24651
rect -5196 24631 -5194 24651
rect -4716 24631 -4714 24651
rect -4500 24631 -4498 24651
rect -4404 24631 -4402 24651
rect -4308 24631 -4306 24651
rect -4164 24631 -4162 24651
rect -3876 24631 -3874 24651
rect -3540 24631 -3538 24651
rect -3468 24631 -3466 24651
rect -3324 24631 -3322 24651
rect -3108 24631 -3106 24651
rect -3012 24631 -3010 24651
rect -2964 24631 -2962 24651
rect -2916 24631 -2914 24651
rect -2868 24631 -2866 24651
rect -2820 24631 -2818 24651
rect -2772 24631 -2770 24651
rect -2676 24631 -2674 24651
rect -2364 24631 -2362 24651
rect -2316 24631 -2314 24651
rect -2265 24648 -2251 24651
rect -2097 24648 -2083 24651
rect -2076 24648 -2073 24651
rect -1980 24631 -1978 24651
rect -1812 24631 -1810 24651
rect -1572 24631 -1570 24651
rect -1476 24631 -1474 24651
rect -1356 24631 -1354 24651
rect -1260 24631 -1258 24651
rect -1236 24631 -1234 24651
rect -1140 24631 -1138 24651
rect -876 24631 -874 24651
rect -660 24631 -658 24651
rect -492 24631 -490 24651
rect -396 24631 -394 24651
rect -383 24646 -380 24651
rect -372 24646 -370 24651
rect -373 24632 -370 24646
rect -276 24648 -274 24651
rect -276 24631 -273 24648
rect -12 24631 -10 24651
rect 84 24631 86 24651
rect 156 24631 158 24651
rect 252 24631 254 24651
rect 348 24631 350 24651
rect 468 24631 470 24651
rect 492 24631 494 24651
rect 564 24631 566 24651
rect 588 24631 590 24651
rect 636 24631 638 24651
rect 660 24631 662 24651
rect 732 24631 734 24651
rect 948 24631 950 24651
rect 1044 24631 1046 24651
rect 1092 24631 1094 24651
rect 1140 24631 1142 24651
rect 1308 24631 1310 24651
rect 1356 24631 1358 24651
rect 1428 24631 1430 24651
rect 1692 24631 1694 24651
rect 1860 24631 1862 24651
rect 2148 24631 2150 24651
rect 2244 24631 2246 24651
rect 2460 24631 2462 24651
rect 2772 24631 2774 24651
rect 2868 24631 2870 24651
rect 2940 24631 2942 24651
rect 2988 24631 2990 24651
rect 3324 24631 3326 24651
rect 3396 24631 3398 24651
rect 3564 24631 3566 24651
rect 3660 24631 3662 24651
rect 3780 24631 3782 24651
rect 4092 24631 4094 24651
rect 4188 24631 4190 24651
rect 4308 24631 4310 24651
rect 4404 24631 4406 24651
rect 4500 24631 4502 24651
rect 4596 24631 4598 24651
rect 4692 24631 4694 24651
rect 4921 24646 4924 24651
rect 4945 24646 4948 24651
rect 4956 24646 4958 24651
rect 4931 24632 4934 24646
rect 4955 24632 4958 24646
rect 4932 24631 4934 24632
rect 4980 24631 4982 24651
rect 5052 24648 5054 24651
rect 5028 24631 5031 24648
rect 5052 24631 5055 24648
rect 5124 24631 5126 24651
rect 5220 24631 5222 24651
rect 5388 24631 5390 24651
rect 5484 24632 5486 24651
rect 5449 24631 5507 24632
rect 5508 24631 5510 24651
rect 5532 24631 5534 24651
rect 5628 24631 5630 24651
rect 5652 24631 5654 24651
rect 5748 24631 5750 24651
rect 5796 24631 5798 24651
rect 5844 24631 5846 24651
rect 5892 24631 5894 24651
rect 6276 24631 6278 24651
rect 6372 24631 6374 24651
rect 6420 24631 6422 24651
rect 6492 24631 6494 24651
rect 6516 24631 6518 24651
rect 6588 24631 6590 24651
rect 6612 24631 6614 24651
rect 6636 24631 6638 24651
rect 6684 24631 6686 24651
rect 6708 24631 6710 24651
rect 6780 24631 6782 24651
rect 6804 24631 6806 24651
rect 6900 24631 6902 24651
rect 6924 24631 6926 24651
rect 7020 24631 7022 24651
rect 7164 24631 7166 24651
rect 7236 24631 7238 24651
rect 7284 24631 7286 24651
rect 7380 24631 7382 24651
rect 7404 24631 7406 24651
rect 7476 24631 7478 24651
rect 7500 24631 7502 24651
rect 7572 24631 7574 24651
rect 7644 24631 7646 24651
rect 7668 24631 7670 24651
rect 7908 24631 7910 24651
rect 8124 24631 8126 24651
rect 8220 24631 8222 24651
rect 8652 24631 8654 24651
rect 8700 24631 8702 24651
rect 8748 24631 8750 24651
rect 8796 24631 8798 24651
rect 8844 24631 8846 24651
rect 8868 24631 8870 24651
rect 9516 24631 9518 24651
rect 9660 24631 9662 24651
rect 9684 24631 9686 24651
rect 9756 24631 9758 24651
rect 9780 24631 9782 24651
rect 9804 24631 9806 24651
rect 9852 24631 9854 24651
rect 9948 24631 9950 24651
rect 10044 24631 10046 24651
rect 10140 24631 10142 24651
rect 10236 24631 10238 24651
rect 10332 24631 10334 24651
rect 10380 24631 10382 24651
rect 10428 24631 10430 24651
rect 10524 24631 10526 24651
rect 10548 24631 10550 24651
rect 10620 24631 10622 24651
rect 10644 24631 10646 24651
rect 10716 24631 10718 24651
rect 10884 24631 10886 24651
rect 10956 24631 10958 24651
rect 11052 24631 11054 24651
rect 11100 24631 11102 24651
rect 11172 24631 11174 24651
rect 11220 24631 11222 24651
rect 11340 24631 11342 24651
rect 11436 24631 11438 24651
rect 11676 24631 11678 24651
rect 11724 24631 11726 24651
rect 11772 24631 11774 24651
rect 11796 24631 11798 24651
rect 12060 24631 12062 24651
rect 12276 24631 12278 24651
rect 12324 24631 12326 24651
rect 12372 24631 12374 24651
rect 12420 24631 12422 24651
rect 12444 24631 12446 24651
rect 12468 24631 12470 24651
rect 12540 24631 12542 24651
rect 12564 24631 12566 24651
rect 12660 24631 12662 24651
rect 12673 24631 12731 24632
rect 12756 24631 12758 24651
rect 12828 24631 12830 24651
rect 12876 24631 12878 24651
rect 12972 24631 12974 24651
rect 13044 24631 13046 24651
rect 13068 24631 13070 24651
rect 13284 24631 13286 24651
rect 13332 24631 13334 24651
rect 13500 24631 13502 24651
rect 13572 24631 13574 24651
rect 13668 24631 13670 24651
rect 13716 24631 13718 24651
rect 13764 24631 13766 24651
rect 13860 24631 13862 24651
rect 13956 24631 13958 24651
rect 14004 24631 14006 24651
rect 14100 24631 14102 24651
rect 14940 24631 14942 24651
rect 15036 24631 15038 24651
rect 15276 24631 15278 24651
rect 15420 24631 15422 24651
rect 15564 24631 15566 24651
rect 15660 24631 15662 24651
rect 15708 24631 15710 24651
rect 15732 24631 15734 24651
rect 15756 24631 15758 24651
rect 15804 24631 15806 24651
rect 15828 24631 15830 24651
rect 15852 24631 15854 24651
rect 15948 24631 15950 24651
rect 15972 24631 15974 24651
rect 16044 24631 16046 24651
rect 16068 24631 16070 24651
rect 16164 24631 16166 24651
rect 16260 24631 16262 24651
rect 16332 24631 16334 24651
rect 16380 24631 16382 24651
rect 16476 24631 16478 24651
rect 16548 24631 16550 24651
rect 16572 24631 16574 24651
rect 16668 24631 16670 24651
rect 16764 24631 16766 24651
rect 16812 24631 16814 24651
rect 16884 24631 16886 24651
rect 16908 24631 16910 24651
rect 16980 24631 16982 24651
rect 17028 24631 17030 24651
rect 17124 24631 17126 24651
rect 17196 24631 17198 24651
rect 17220 24631 17222 24651
rect 17292 24631 17294 24651
rect 17316 24631 17318 24651
rect 17964 24631 17966 24651
rect 18060 24631 18062 24651
rect 18132 24631 18134 24651
rect 18228 24631 18230 24651
rect 18492 24631 18494 24651
rect 18540 24631 18542 24651
rect 18636 24631 18638 24651
rect 18732 24631 18734 24651
rect 18828 24631 18830 24651
rect 18924 24631 18926 24651
rect 18972 24631 18974 24651
rect 19020 24631 19022 24651
rect 19068 24631 19070 24651
rect 19140 24631 19142 24651
rect 19164 24631 19166 24651
rect 19236 24631 19238 24651
rect 19260 24631 19262 24651
rect 19788 24631 19790 24651
rect 19836 24631 19838 24651
rect 19860 24631 19862 24651
rect 19884 24631 19886 24651
rect 19956 24631 19958 24651
rect 19980 24631 19982 24651
rect 20004 24631 20006 24651
rect 20052 24631 20054 24651
rect 20076 24631 20078 24651
rect 20100 24631 20102 24651
rect 20172 24631 20174 24651
rect 20196 24631 20198 24651
rect 20292 24631 20294 24651
rect 20388 24631 20390 24651
rect 20412 24631 20414 24651
rect 20508 24631 20510 24651
rect 20532 24631 20534 24651
rect 20604 24631 20606 24651
rect 20628 24631 20630 24651
rect 20892 24631 20894 24651
rect 20964 24631 20966 24651
rect 20988 24631 20990 24651
rect 21108 24631 21110 24651
rect 21204 24631 21206 24651
rect 21300 24631 21302 24651
rect 21324 24631 21326 24651
rect 21444 24631 21446 24651
rect 21468 24631 21470 24651
rect 21564 24631 21566 24651
rect 21588 24631 21590 24651
rect 21684 24631 21686 24651
rect 21708 24631 21710 24651
rect 22068 24631 22070 24651
rect 22188 24631 22190 24651
rect 22212 24632 22214 24651
rect 22201 24631 22235 24632
rect -10449 24627 5021 24631
rect -10449 24624 -10435 24627
rect -10007 24607 -9973 24608
rect -9900 24607 -9898 24627
rect -9732 24608 -9730 24627
rect -9743 24607 -9709 24608
rect -9636 24607 -9634 24627
rect -9540 24607 -9538 24627
rect -9444 24607 -9442 24627
rect -9348 24607 -9346 24627
rect -9228 24607 -9226 24627
rect -9108 24607 -9106 24627
rect -9012 24607 -9010 24627
rect -8916 24607 -8914 24627
rect -8628 24607 -8626 24627
rect -8532 24607 -8530 24627
rect -8436 24607 -8434 24627
rect -8340 24607 -8338 24627
rect -8124 24607 -8122 24627
rect -7857 24624 -7843 24627
rect -7764 24607 -7762 24627
rect -7524 24607 -7522 24627
rect -7356 24607 -7354 24627
rect -7308 24607 -7306 24627
rect -7140 24607 -7138 24627
rect -6969 24624 -6955 24627
rect -6948 24624 -6945 24627
rect -6852 24607 -6850 24627
rect -6732 24607 -6730 24627
rect -6705 24624 -6691 24627
rect -6516 24607 -6514 24627
rect -6359 24607 -6301 24608
rect -5892 24607 -5890 24627
rect -5436 24607 -5434 24627
rect -5340 24607 -5338 24627
rect -5196 24607 -5194 24627
rect -4716 24607 -4714 24627
rect -4500 24607 -4498 24627
rect -4404 24607 -4402 24627
rect -4308 24607 -4306 24627
rect -4164 24607 -4162 24627
rect -3876 24607 -3874 24627
rect -3540 24607 -3538 24627
rect -3468 24607 -3466 24627
rect -3324 24607 -3322 24627
rect -3108 24607 -3106 24627
rect -3012 24607 -3010 24627
rect -2964 24607 -2962 24627
rect -2916 24607 -2914 24627
rect -2868 24607 -2866 24627
rect -2820 24607 -2818 24627
rect -2772 24607 -2770 24627
rect -2676 24607 -2674 24627
rect -2364 24607 -2362 24627
rect -2316 24607 -2314 24627
rect -1980 24607 -1978 24627
rect -1812 24607 -1810 24627
rect -1572 24607 -1570 24627
rect -1476 24607 -1474 24627
rect -1356 24607 -1354 24627
rect -1260 24607 -1258 24627
rect -1236 24607 -1234 24627
rect -1140 24607 -1138 24627
rect -876 24607 -874 24627
rect -660 24607 -658 24627
rect -492 24607 -490 24627
rect -396 24607 -394 24627
rect -297 24624 -283 24627
rect -276 24624 -273 24627
rect -12 24607 -10 24627
rect 84 24607 86 24627
rect 156 24607 158 24627
rect 252 24607 254 24627
rect 348 24607 350 24627
rect 468 24607 470 24627
rect 492 24607 494 24627
rect 564 24607 566 24627
rect 588 24607 590 24627
rect 636 24607 638 24627
rect 660 24607 662 24627
rect 732 24607 734 24627
rect 948 24607 950 24627
rect 1044 24607 1046 24627
rect 1092 24607 1094 24627
rect 1140 24607 1142 24627
rect 1308 24607 1310 24627
rect 1356 24607 1358 24627
rect 1428 24607 1430 24627
rect 1692 24607 1694 24627
rect 1860 24607 1862 24627
rect 2148 24607 2150 24627
rect 2244 24607 2246 24627
rect 2460 24607 2462 24627
rect 2772 24607 2774 24627
rect 2868 24607 2870 24627
rect 2940 24607 2942 24627
rect 2988 24607 2990 24627
rect 3324 24607 3326 24627
rect 3396 24607 3398 24627
rect 3564 24607 3566 24627
rect 3660 24607 3662 24627
rect 3780 24607 3782 24627
rect 4092 24607 4094 24627
rect 4188 24607 4190 24627
rect 4308 24607 4310 24627
rect 4404 24607 4406 24627
rect 4500 24607 4502 24627
rect 4596 24607 4598 24627
rect 4692 24607 4694 24627
rect 4932 24607 4934 24627
rect 4980 24607 4982 24627
rect 5007 24624 5021 24627
rect 5028 24627 22235 24631
rect 5028 24624 5045 24627
rect 5052 24624 5055 24627
rect 5028 24607 5030 24624
rect 5124 24607 5126 24627
rect 5220 24607 5222 24627
rect 5388 24607 5390 24627
rect 5473 24622 5476 24627
rect 5484 24622 5486 24627
rect 5483 24608 5486 24622
rect 5508 24607 5510 24627
rect 5532 24607 5534 24627
rect 5556 24607 5559 24624
rect 5628 24607 5630 24627
rect 5652 24607 5654 24627
rect 5748 24607 5750 24627
rect 5796 24607 5798 24627
rect 5844 24607 5846 24627
rect 5892 24607 5894 24627
rect 6276 24607 6278 24627
rect 6372 24607 6374 24627
rect 6420 24607 6422 24627
rect 6492 24607 6494 24627
rect 6516 24607 6518 24627
rect 6588 24607 6590 24627
rect 6612 24607 6614 24627
rect 6636 24607 6638 24627
rect 6684 24607 6686 24627
rect 6708 24607 6710 24627
rect 6780 24607 6782 24627
rect 6804 24607 6806 24627
rect 6900 24607 6902 24627
rect 6924 24607 6926 24627
rect 7020 24607 7022 24627
rect 7164 24607 7166 24627
rect 7236 24607 7238 24627
rect 7284 24607 7286 24627
rect 7380 24607 7382 24627
rect 7404 24607 7406 24627
rect 7476 24607 7478 24627
rect 7500 24607 7502 24627
rect 7572 24607 7574 24627
rect 7644 24607 7646 24627
rect 7668 24607 7670 24627
rect 7908 24607 7910 24627
rect 8124 24607 8126 24627
rect 8220 24607 8222 24627
rect 8652 24607 8654 24627
rect 8700 24607 8702 24627
rect 8748 24607 8750 24627
rect 8796 24607 8798 24627
rect 8844 24607 8846 24627
rect 8868 24607 8870 24627
rect 9516 24607 9518 24627
rect 9660 24607 9662 24627
rect 9684 24607 9686 24627
rect 9756 24607 9758 24627
rect 9780 24607 9782 24627
rect 9804 24607 9806 24627
rect 9852 24607 9854 24627
rect 9948 24607 9950 24627
rect 10044 24607 10046 24627
rect 10140 24607 10142 24627
rect 10236 24607 10238 24627
rect 10332 24607 10334 24627
rect 10380 24607 10382 24627
rect 10428 24607 10430 24627
rect 10524 24607 10526 24627
rect 10548 24607 10550 24627
rect 10620 24607 10622 24627
rect 10644 24607 10646 24627
rect 10716 24607 10718 24627
rect 10884 24607 10886 24627
rect 10956 24607 10958 24627
rect 11052 24607 11054 24627
rect 11100 24607 11102 24627
rect 11172 24607 11174 24627
rect 11220 24607 11222 24627
rect 11340 24607 11342 24627
rect 11436 24607 11438 24627
rect 11676 24607 11678 24627
rect 11724 24607 11726 24627
rect 11772 24607 11774 24627
rect 11796 24607 11798 24627
rect 12060 24607 12062 24627
rect 12276 24607 12278 24627
rect 12324 24607 12326 24627
rect 12372 24607 12374 24627
rect 12420 24607 12422 24627
rect 12444 24607 12446 24627
rect 12468 24607 12470 24627
rect 12540 24607 12542 24627
rect 12564 24607 12566 24627
rect 12660 24607 12662 24627
rect 12756 24607 12758 24627
rect 12780 24607 12783 24624
rect 12828 24607 12830 24627
rect 12876 24607 12878 24627
rect 12972 24607 12974 24627
rect 13044 24607 13046 24627
rect 13068 24607 13070 24627
rect 13284 24607 13286 24627
rect 13332 24607 13334 24627
rect 13500 24607 13502 24627
rect 13572 24607 13574 24627
rect 13668 24607 13670 24627
rect 13716 24607 13718 24627
rect 13764 24607 13766 24627
rect 13860 24607 13862 24627
rect 13956 24607 13958 24627
rect 14004 24607 14006 24627
rect 14100 24607 14102 24627
rect 14940 24607 14942 24627
rect 15036 24607 15038 24627
rect 15276 24607 15278 24627
rect 15420 24607 15422 24627
rect 15564 24607 15566 24627
rect 15660 24607 15662 24627
rect 15708 24607 15710 24627
rect 15732 24607 15734 24627
rect 15756 24607 15758 24627
rect 15804 24607 15806 24627
rect 15828 24607 15830 24627
rect 15852 24607 15854 24627
rect 15948 24607 15950 24627
rect 15972 24607 15974 24627
rect 16044 24607 16046 24627
rect 16068 24607 16070 24627
rect 16164 24607 16166 24627
rect 16260 24607 16262 24627
rect 16332 24607 16334 24627
rect 16380 24607 16382 24627
rect 16476 24607 16478 24627
rect 16548 24607 16550 24627
rect 16572 24607 16574 24627
rect 16668 24607 16670 24627
rect 16764 24607 16766 24627
rect 16812 24607 16814 24627
rect 16884 24607 16886 24627
rect 16908 24607 16910 24627
rect 16980 24607 16982 24627
rect 17028 24607 17030 24627
rect 17124 24607 17126 24627
rect 17196 24607 17198 24627
rect 17220 24607 17222 24627
rect 17292 24607 17294 24627
rect 17316 24607 17318 24627
rect 17964 24607 17966 24627
rect 18060 24607 18062 24627
rect 18132 24607 18134 24627
rect 18228 24607 18230 24627
rect 18492 24607 18494 24627
rect 18540 24607 18542 24627
rect 18636 24607 18638 24627
rect 18732 24607 18734 24627
rect 18828 24607 18830 24627
rect 18924 24607 18926 24627
rect 18972 24607 18974 24627
rect 19020 24607 19022 24627
rect 19068 24607 19070 24627
rect 19140 24607 19142 24627
rect 19164 24607 19166 24627
rect 19236 24607 19238 24627
rect 19260 24607 19262 24627
rect 19788 24607 19790 24627
rect 19836 24607 19838 24627
rect 19860 24607 19862 24627
rect 19884 24607 19886 24627
rect 19956 24607 19958 24627
rect 19980 24607 19982 24627
rect 20004 24607 20006 24627
rect 20052 24607 20054 24627
rect 20076 24607 20078 24627
rect 20100 24607 20102 24627
rect 20172 24607 20174 24627
rect 20196 24607 20198 24627
rect 20292 24607 20294 24627
rect 20388 24607 20390 24627
rect 20412 24607 20414 24627
rect 20508 24607 20510 24627
rect 20532 24607 20534 24627
rect 20604 24607 20606 24627
rect 20628 24607 20630 24627
rect 20892 24607 20894 24627
rect 20964 24607 20966 24627
rect 20988 24607 20990 24627
rect 21108 24607 21110 24627
rect 21204 24607 21206 24627
rect 21300 24607 21302 24627
rect 21324 24607 21326 24627
rect 21444 24607 21446 24627
rect 21468 24607 21470 24627
rect 21564 24607 21566 24627
rect 21588 24607 21590 24627
rect 21684 24607 21686 24627
rect 21708 24607 21710 24627
rect 22068 24607 22070 24627
rect 22188 24608 22190 24627
rect 22201 24622 22204 24627
rect 22212 24622 22214 24627
rect 22211 24608 22214 24622
rect 22177 24607 22211 24608
rect -10007 24603 5549 24607
rect -9900 24600 -9898 24603
rect -9900 24584 -9897 24600
rect -9743 24598 -9740 24603
rect -9732 24598 -9730 24603
rect -9733 24584 -9730 24598
rect -9636 24600 -9634 24603
rect -9911 24583 -9877 24584
rect -9636 24583 -9633 24600
rect -9540 24583 -9538 24603
rect -9444 24583 -9442 24603
rect -9348 24583 -9346 24603
rect -9228 24583 -9226 24603
rect -9108 24583 -9106 24603
rect -9012 24583 -9010 24603
rect -8916 24583 -8914 24603
rect -8628 24583 -8626 24603
rect -8532 24583 -8530 24603
rect -8436 24583 -8434 24603
rect -8340 24583 -8338 24603
rect -8124 24583 -8122 24603
rect -7764 24583 -7762 24603
rect -7655 24583 -7597 24584
rect -7524 24583 -7522 24603
rect -7356 24583 -7354 24603
rect -7308 24583 -7306 24603
rect -7140 24583 -7138 24603
rect -6852 24583 -6850 24603
rect -6732 24583 -6730 24603
rect -6516 24583 -6514 24603
rect -6359 24598 -6356 24603
rect -6349 24584 -6346 24598
rect -6348 24583 -6346 24584
rect -6252 24583 -6249 24600
rect -5892 24583 -5890 24603
rect -5436 24583 -5434 24603
rect -5340 24583 -5338 24603
rect -5196 24583 -5194 24603
rect -4716 24583 -4714 24603
rect -4500 24583 -4498 24603
rect -4404 24584 -4402 24603
rect -4415 24583 -4381 24584
rect -4308 24583 -4306 24603
rect -4164 24583 -4162 24603
rect -3876 24583 -3874 24603
rect -3540 24583 -3538 24603
rect -3468 24583 -3466 24603
rect -3324 24583 -3322 24603
rect -3108 24583 -3106 24603
rect -3012 24583 -3010 24603
rect -2964 24583 -2962 24603
rect -2916 24583 -2914 24603
rect -2868 24583 -2866 24603
rect -2820 24583 -2818 24603
rect -2772 24583 -2770 24603
rect -2676 24583 -2674 24603
rect -2447 24583 -2389 24584
rect -2364 24583 -2362 24603
rect -2316 24583 -2314 24603
rect -1980 24583 -1978 24603
rect -1812 24583 -1810 24603
rect -1572 24583 -1570 24603
rect -1476 24583 -1474 24603
rect -1356 24583 -1354 24603
rect -1260 24583 -1258 24603
rect -1236 24583 -1234 24603
rect -1140 24583 -1138 24603
rect -876 24583 -874 24603
rect -660 24583 -658 24603
rect -492 24583 -490 24603
rect -396 24583 -394 24603
rect -12 24583 -10 24603
rect 84 24583 86 24603
rect 156 24583 158 24603
rect 252 24583 254 24603
rect 348 24583 350 24603
rect 468 24583 470 24603
rect 492 24583 494 24603
rect 564 24583 566 24603
rect 588 24583 590 24603
rect 636 24583 638 24603
rect 660 24583 662 24603
rect 732 24583 734 24603
rect 948 24583 950 24603
rect 1044 24583 1046 24603
rect 1092 24583 1094 24603
rect 1140 24583 1142 24603
rect 1308 24583 1310 24603
rect 1356 24583 1358 24603
rect 1428 24583 1430 24603
rect 1692 24583 1694 24603
rect 1860 24583 1862 24603
rect 1945 24583 2003 24584
rect 2148 24583 2150 24603
rect 2244 24583 2246 24603
rect 2460 24583 2462 24603
rect 2772 24583 2774 24603
rect 2868 24583 2870 24603
rect 2940 24583 2942 24603
rect 2988 24583 2990 24603
rect 3324 24583 3326 24603
rect 3396 24583 3398 24603
rect 3564 24583 3566 24603
rect 3660 24583 3662 24603
rect 3780 24583 3782 24603
rect 4092 24583 4094 24603
rect 4188 24583 4190 24603
rect 4308 24583 4310 24603
rect 4404 24583 4406 24603
rect 4500 24583 4502 24603
rect 4596 24583 4598 24603
rect 4692 24583 4694 24603
rect 4932 24583 4934 24603
rect 4980 24583 4982 24603
rect 5028 24583 5030 24603
rect 5124 24583 5126 24603
rect 5220 24583 5222 24603
rect 5388 24583 5390 24603
rect 5508 24583 5510 24603
rect 5532 24583 5534 24603
rect 5535 24600 5549 24603
rect 5556 24603 12773 24607
rect 5556 24600 5573 24603
rect 5556 24583 5558 24600
rect 5628 24583 5630 24603
rect 5652 24583 5654 24603
rect 5748 24583 5750 24603
rect 5796 24583 5798 24603
rect 5844 24583 5846 24603
rect 5892 24583 5894 24603
rect 6276 24583 6278 24603
rect 6372 24583 6374 24603
rect 6420 24583 6422 24603
rect 6492 24583 6494 24603
rect 6516 24583 6518 24603
rect 6588 24583 6590 24603
rect 6612 24583 6614 24603
rect 6636 24583 6638 24603
rect 6684 24583 6686 24603
rect 6708 24583 6710 24603
rect 6780 24583 6782 24603
rect 6804 24583 6806 24603
rect 6900 24583 6902 24603
rect 6924 24583 6926 24603
rect 7020 24583 7022 24603
rect 7164 24583 7166 24603
rect 7236 24583 7238 24603
rect 7284 24583 7286 24603
rect 7380 24583 7382 24603
rect 7404 24583 7406 24603
rect 7476 24583 7478 24603
rect 7500 24583 7502 24603
rect 7572 24583 7574 24603
rect 7644 24583 7646 24603
rect 7668 24583 7670 24603
rect 7908 24583 7910 24603
rect 8124 24583 8126 24603
rect 8220 24583 8222 24603
rect 8652 24583 8654 24603
rect 8700 24583 8702 24603
rect 8748 24583 8750 24603
rect 8796 24583 8798 24603
rect 8844 24583 8846 24603
rect 8868 24583 8870 24603
rect 9516 24583 9518 24603
rect 9660 24583 9662 24603
rect 9684 24583 9686 24603
rect 9756 24583 9758 24603
rect 9780 24583 9782 24603
rect 9804 24583 9806 24603
rect 9852 24584 9854 24603
rect 9817 24583 9875 24584
rect 9948 24583 9950 24603
rect 10044 24583 10046 24603
rect 10140 24583 10142 24603
rect 10236 24583 10238 24603
rect 10332 24583 10334 24603
rect 10380 24583 10382 24603
rect 10428 24583 10430 24603
rect 10524 24583 10526 24603
rect 10548 24583 10550 24603
rect 10620 24583 10622 24603
rect 10644 24583 10646 24603
rect 10716 24583 10718 24603
rect 10884 24583 10886 24603
rect 10956 24583 10958 24603
rect 11052 24583 11054 24603
rect 11100 24583 11102 24603
rect 11172 24583 11174 24603
rect 11220 24583 11222 24603
rect 11340 24583 11342 24603
rect 11436 24583 11438 24603
rect 11676 24583 11678 24603
rect 11724 24583 11726 24603
rect 11772 24583 11774 24603
rect 11796 24583 11798 24603
rect 12060 24583 12062 24603
rect 12276 24583 12278 24603
rect 12324 24583 12326 24603
rect 12372 24583 12374 24603
rect 12420 24583 12422 24603
rect 12444 24583 12446 24603
rect 12468 24583 12470 24603
rect 12540 24583 12542 24603
rect 12564 24583 12566 24603
rect 12660 24583 12662 24603
rect 12756 24583 12758 24603
rect 12759 24600 12773 24603
rect 12780 24603 22211 24607
rect 12780 24600 12797 24603
rect 12780 24583 12782 24600
rect 12828 24583 12830 24603
rect 12876 24583 12878 24603
rect 12972 24583 12974 24603
rect 13044 24583 13046 24603
rect 13068 24583 13070 24603
rect 13284 24583 13286 24603
rect 13332 24583 13334 24603
rect 13500 24583 13502 24603
rect 13572 24583 13574 24603
rect 13668 24583 13670 24603
rect 13716 24583 13718 24603
rect 13764 24583 13766 24603
rect 13860 24583 13862 24603
rect 13956 24583 13958 24603
rect 14004 24583 14006 24603
rect 14100 24583 14102 24603
rect 14940 24583 14942 24603
rect 15036 24583 15038 24603
rect 15276 24583 15278 24603
rect 15420 24583 15422 24603
rect 15564 24583 15566 24603
rect 15660 24583 15662 24603
rect 15708 24583 15710 24603
rect 15732 24583 15734 24603
rect 15756 24583 15758 24603
rect 15804 24583 15806 24603
rect 15828 24583 15830 24603
rect 15852 24583 15854 24603
rect 15948 24583 15950 24603
rect 15972 24583 15974 24603
rect 16044 24583 16046 24603
rect 16068 24583 16070 24603
rect 16164 24583 16166 24603
rect 16260 24583 16262 24603
rect 16332 24583 16334 24603
rect 16380 24583 16382 24603
rect 16476 24583 16478 24603
rect 16548 24583 16550 24603
rect 16572 24583 16574 24603
rect 16668 24583 16670 24603
rect 16764 24583 16766 24603
rect 16812 24583 16814 24603
rect 16884 24583 16886 24603
rect 16908 24583 16910 24603
rect 16980 24583 16982 24603
rect 17028 24583 17030 24603
rect 17124 24583 17126 24603
rect 17196 24583 17198 24603
rect 17220 24583 17222 24603
rect 17292 24583 17294 24603
rect 17316 24583 17318 24603
rect 17964 24583 17966 24603
rect 18060 24583 18062 24603
rect 18132 24583 18134 24603
rect 18228 24583 18230 24603
rect 18492 24583 18494 24603
rect 18540 24583 18542 24603
rect 18636 24583 18638 24603
rect 18732 24583 18734 24603
rect 18828 24583 18830 24603
rect 18924 24583 18926 24603
rect 18972 24583 18974 24603
rect 19020 24583 19022 24603
rect 19068 24583 19070 24603
rect 19140 24583 19142 24603
rect 19164 24583 19166 24603
rect 19236 24583 19238 24603
rect 19260 24583 19262 24603
rect 19788 24583 19790 24603
rect 19836 24583 19838 24603
rect 19860 24583 19862 24603
rect 19884 24583 19886 24603
rect 19956 24583 19958 24603
rect 19980 24583 19982 24603
rect 20004 24583 20006 24603
rect 20052 24583 20054 24603
rect 20076 24583 20078 24603
rect 20100 24583 20102 24603
rect 20172 24583 20174 24603
rect 20196 24583 20198 24603
rect 20292 24583 20294 24603
rect 20388 24583 20390 24603
rect 20412 24583 20414 24603
rect 20508 24583 20510 24603
rect 20532 24583 20534 24603
rect 20604 24583 20606 24603
rect 20628 24583 20630 24603
rect 20892 24583 20894 24603
rect 20964 24583 20966 24603
rect 20988 24583 20990 24603
rect 21108 24583 21110 24603
rect 21204 24583 21206 24603
rect 21300 24583 21302 24603
rect 21324 24583 21326 24603
rect 21444 24583 21446 24603
rect 21468 24583 21470 24603
rect 21564 24583 21566 24603
rect 21588 24583 21590 24603
rect 21684 24583 21686 24603
rect 21708 24583 21710 24603
rect 22068 24583 22070 24603
rect 22177 24598 22180 24603
rect 22188 24598 22190 24603
rect 22187 24584 22190 24598
rect 22105 24583 22139 24584
rect -9911 24579 -6259 24583
rect -9911 24576 -9907 24579
rect -9900 24576 -9897 24579
rect -9657 24576 -9643 24579
rect -9636 24576 -9633 24579
rect -9825 24559 -9805 24560
rect -9540 24559 -9538 24579
rect -9444 24559 -9442 24579
rect -9348 24559 -9346 24579
rect -9228 24559 -9226 24579
rect -9108 24559 -9106 24579
rect -9012 24559 -9010 24579
rect -8916 24559 -8914 24579
rect -8628 24559 -8626 24579
rect -8532 24559 -8530 24579
rect -8436 24559 -8434 24579
rect -8340 24559 -8338 24579
rect -8124 24559 -8122 24579
rect -7764 24559 -7762 24579
rect -7524 24576 -7522 24579
rect -7524 24559 -7521 24576
rect -7356 24559 -7354 24579
rect -7308 24559 -7306 24579
rect -7140 24559 -7138 24579
rect -6852 24559 -6850 24579
rect -6732 24559 -6730 24579
rect -6516 24559 -6514 24579
rect -6348 24559 -6346 24579
rect -6273 24576 -6259 24579
rect -6252 24579 22139 24583
rect -6252 24576 -6235 24579
rect -6252 24559 -6250 24576
rect -5892 24559 -5890 24579
rect -5436 24559 -5434 24579
rect -5340 24559 -5338 24579
rect -5196 24559 -5194 24579
rect -4716 24559 -4714 24579
rect -4500 24559 -4498 24579
rect -4415 24574 -4412 24579
rect -4404 24574 -4402 24579
rect -4405 24560 -4402 24574
rect -4308 24576 -4306 24579
rect -4308 24559 -4305 24576
rect -4295 24559 -4237 24560
rect -4164 24559 -4162 24579
rect -3876 24559 -3874 24579
rect -3540 24559 -3538 24579
rect -3468 24559 -3466 24579
rect -3324 24559 -3322 24579
rect -3108 24559 -3106 24579
rect -3012 24559 -3010 24579
rect -2964 24559 -2962 24579
rect -2916 24559 -2914 24579
rect -2868 24559 -2866 24579
rect -2820 24559 -2818 24579
rect -2772 24559 -2770 24579
rect -2676 24559 -2674 24579
rect -2364 24559 -2362 24579
rect -2316 24576 -2314 24579
rect -2316 24559 -2313 24576
rect -1980 24559 -1978 24579
rect -1812 24559 -1810 24579
rect -1572 24559 -1570 24579
rect -1476 24559 -1474 24579
rect -1356 24559 -1354 24579
rect -1260 24559 -1258 24579
rect -1236 24559 -1234 24579
rect -1140 24559 -1138 24579
rect -876 24559 -874 24579
rect -660 24559 -658 24579
rect -492 24560 -490 24579
rect -503 24559 -469 24560
rect -396 24559 -394 24579
rect -287 24559 -253 24560
rect -12 24559 -10 24579
rect 84 24559 86 24579
rect 156 24559 158 24579
rect 252 24559 254 24579
rect 348 24559 350 24579
rect 468 24559 470 24579
rect 492 24559 494 24579
rect 564 24559 566 24579
rect 588 24559 590 24579
rect 636 24559 638 24579
rect 660 24559 662 24579
rect 732 24559 734 24579
rect 948 24559 950 24579
rect 1044 24559 1046 24579
rect 1092 24559 1094 24579
rect 1140 24559 1142 24579
rect 1308 24559 1310 24579
rect 1356 24559 1358 24579
rect 1428 24559 1430 24579
rect 1692 24559 1694 24579
rect 1860 24559 1862 24579
rect 1945 24574 1948 24579
rect 1955 24560 1958 24574
rect 1956 24559 1958 24560
rect 2052 24559 2055 24576
rect 2148 24559 2150 24579
rect 2244 24559 2246 24579
rect 2460 24559 2462 24579
rect 2772 24559 2774 24579
rect 2868 24559 2870 24579
rect 2940 24559 2942 24579
rect 2988 24559 2990 24579
rect 3324 24559 3326 24579
rect 3396 24559 3398 24579
rect 3564 24559 3566 24579
rect 3660 24559 3662 24579
rect 3780 24559 3782 24579
rect 4092 24559 4094 24579
rect 4188 24559 4190 24579
rect 4308 24559 4310 24579
rect 4404 24559 4406 24579
rect 4500 24559 4502 24579
rect 4596 24559 4598 24579
rect 4692 24559 4694 24579
rect 4932 24559 4934 24579
rect 4980 24559 4982 24579
rect 5028 24559 5030 24579
rect 5124 24559 5126 24579
rect 5220 24559 5222 24579
rect 5388 24559 5390 24579
rect 5508 24559 5510 24579
rect 5532 24559 5534 24579
rect 5556 24559 5558 24579
rect 5628 24559 5630 24579
rect 5652 24559 5654 24579
rect 5748 24559 5750 24579
rect 5796 24559 5798 24579
rect 5844 24559 5846 24579
rect 5892 24559 5894 24579
rect 6276 24559 6278 24579
rect 6372 24559 6374 24579
rect 6420 24559 6422 24579
rect 6492 24559 6494 24579
rect 6516 24559 6518 24579
rect 6588 24559 6590 24579
rect 6612 24559 6614 24579
rect 6636 24559 6638 24579
rect 6684 24559 6686 24579
rect 6708 24559 6710 24579
rect 6780 24559 6782 24579
rect 6804 24559 6806 24579
rect 6900 24559 6902 24579
rect 6924 24559 6926 24579
rect 7020 24559 7022 24579
rect 7164 24559 7166 24579
rect 7236 24559 7238 24579
rect 7284 24559 7286 24579
rect 7380 24559 7382 24579
rect 7404 24559 7406 24579
rect 7476 24559 7478 24579
rect 7500 24559 7502 24579
rect 7572 24559 7574 24579
rect 7644 24559 7646 24579
rect 7668 24559 7670 24579
rect 7908 24559 7910 24579
rect 8124 24559 8126 24579
rect 8220 24559 8222 24579
rect 8652 24559 8654 24579
rect 8700 24559 8702 24579
rect 8748 24559 8750 24579
rect 8796 24559 8798 24579
rect 8844 24559 8846 24579
rect 8868 24559 8870 24579
rect 9516 24559 9518 24579
rect 9660 24559 9662 24579
rect 9684 24559 9686 24579
rect 9756 24559 9758 24579
rect 9780 24559 9782 24579
rect 9804 24559 9806 24579
rect 9841 24574 9844 24579
rect 9852 24574 9854 24579
rect 9851 24560 9854 24574
rect 9948 24576 9950 24579
rect 9948 24559 9951 24576
rect 10044 24559 10046 24579
rect 10140 24559 10142 24579
rect 10236 24559 10238 24579
rect 10332 24559 10334 24579
rect 10380 24559 10382 24579
rect 10428 24559 10430 24579
rect 10524 24559 10526 24579
rect 10548 24559 10550 24579
rect 10620 24559 10622 24579
rect 10644 24559 10646 24579
rect 10716 24559 10718 24579
rect 10884 24559 10886 24579
rect 10956 24559 10958 24579
rect 11052 24559 11054 24579
rect 11100 24559 11102 24579
rect 11172 24559 11174 24579
rect 11220 24559 11222 24579
rect 11340 24559 11342 24579
rect 11436 24559 11438 24579
rect 11676 24559 11678 24579
rect 11724 24559 11726 24579
rect 11772 24559 11774 24579
rect 11796 24559 11798 24579
rect 12060 24559 12062 24579
rect 12276 24559 12278 24579
rect 12324 24559 12326 24579
rect 12372 24559 12374 24579
rect 12420 24559 12422 24579
rect 12444 24560 12446 24579
rect 12433 24559 12467 24560
rect 12468 24559 12470 24579
rect 12540 24559 12542 24579
rect 12564 24559 12566 24579
rect 12660 24559 12662 24579
rect 12756 24559 12758 24579
rect 12780 24559 12782 24579
rect 12828 24559 12830 24579
rect 12876 24559 12878 24579
rect 12972 24559 12974 24579
rect 13044 24559 13046 24579
rect 13068 24559 13070 24579
rect 13284 24559 13286 24579
rect 13332 24559 13334 24579
rect 13500 24559 13502 24579
rect 13572 24559 13574 24579
rect 13668 24559 13670 24579
rect 13716 24559 13718 24579
rect 13764 24560 13766 24579
rect 13729 24559 13787 24560
rect 13860 24559 13862 24579
rect 13956 24559 13958 24579
rect 14004 24559 14006 24579
rect 14100 24559 14102 24579
rect 14940 24559 14942 24579
rect 15036 24559 15038 24579
rect 15276 24559 15278 24579
rect 15420 24559 15422 24579
rect 15564 24559 15566 24579
rect 15660 24559 15662 24579
rect 15708 24559 15710 24579
rect 15732 24559 15734 24579
rect 15756 24559 15758 24579
rect 15804 24559 15806 24579
rect 15828 24559 15830 24579
rect 15852 24559 15854 24579
rect 15948 24559 15950 24579
rect 15972 24559 15974 24579
rect 16044 24559 16046 24579
rect 16068 24559 16070 24579
rect 16164 24559 16166 24579
rect 16260 24559 16262 24579
rect 16332 24559 16334 24579
rect 16380 24559 16382 24579
rect 16476 24559 16478 24579
rect 16548 24559 16550 24579
rect 16572 24559 16574 24579
rect 16668 24559 16670 24579
rect 16764 24559 16766 24579
rect 16812 24559 16814 24579
rect 16884 24559 16886 24579
rect 16908 24559 16910 24579
rect 16980 24559 16982 24579
rect 17028 24559 17030 24579
rect 17124 24559 17126 24579
rect 17196 24559 17198 24579
rect 17220 24559 17222 24579
rect 17292 24559 17294 24579
rect 17316 24559 17318 24579
rect 17964 24559 17966 24579
rect 18060 24559 18062 24579
rect 18132 24559 18134 24579
rect 18228 24559 18230 24579
rect 18492 24559 18494 24579
rect 18540 24559 18542 24579
rect 18636 24559 18638 24579
rect 18732 24559 18734 24579
rect 18828 24559 18830 24579
rect 18924 24559 18926 24579
rect 18972 24559 18974 24579
rect 19020 24559 19022 24579
rect 19068 24559 19070 24579
rect 19140 24559 19142 24579
rect 19164 24559 19166 24579
rect 19236 24559 19238 24579
rect 19260 24559 19262 24579
rect 19788 24559 19790 24579
rect 19836 24559 19838 24579
rect 19860 24559 19862 24579
rect 19884 24559 19886 24579
rect 19956 24559 19958 24579
rect 19980 24559 19982 24579
rect 20004 24559 20006 24579
rect 20052 24559 20054 24579
rect 20076 24559 20078 24579
rect 20100 24559 20102 24579
rect 20172 24559 20174 24579
rect 20196 24559 20198 24579
rect 20292 24559 20294 24579
rect 20388 24559 20390 24579
rect 20412 24559 20414 24579
rect 20508 24559 20510 24579
rect 20532 24559 20534 24579
rect 20604 24559 20606 24579
rect 20628 24559 20630 24579
rect 20892 24559 20894 24579
rect 20964 24559 20966 24579
rect 20988 24559 20990 24579
rect 21108 24559 21110 24579
rect 21204 24559 21206 24579
rect 21300 24559 21302 24579
rect 21324 24559 21326 24579
rect 21444 24559 21446 24579
rect 21468 24559 21470 24579
rect 21564 24559 21566 24579
rect 21588 24559 21590 24579
rect 21684 24559 21686 24579
rect 21708 24559 21710 24579
rect 22068 24559 22070 24579
rect 22081 24559 22115 24560
rect -9825 24555 -7555 24559
rect -9825 24552 -9811 24555
rect -9540 24535 -9538 24555
rect -9444 24535 -9442 24555
rect -9348 24535 -9346 24555
rect -9228 24535 -9226 24555
rect -9108 24535 -9106 24555
rect -9012 24535 -9010 24555
rect -8916 24535 -8914 24555
rect -8628 24535 -8626 24555
rect -8532 24535 -8530 24555
rect -8436 24535 -8434 24555
rect -8340 24535 -8338 24555
rect -8124 24535 -8122 24555
rect -7764 24535 -7762 24555
rect -7569 24552 -7555 24555
rect -7545 24555 -2347 24559
rect -7545 24552 -7531 24555
rect -7524 24552 -7521 24555
rect -7356 24535 -7354 24555
rect -7308 24535 -7306 24555
rect -7140 24535 -7138 24555
rect -6852 24535 -6850 24555
rect -6732 24535 -6730 24555
rect -6516 24535 -6514 24555
rect -6348 24535 -6346 24555
rect -6252 24535 -6250 24555
rect -5892 24535 -5890 24555
rect -5759 24535 -5725 24536
rect -5436 24535 -5434 24555
rect -5340 24535 -5338 24555
rect -5303 24535 -5269 24536
rect -5196 24535 -5194 24555
rect -4716 24535 -4714 24555
rect -4500 24535 -4498 24555
rect -4329 24552 -4315 24555
rect -4308 24552 -4305 24555
rect -4295 24550 -4292 24555
rect -4164 24552 -4162 24555
rect -4285 24536 -4282 24550
rect -4284 24535 -4282 24536
rect -4164 24535 -4161 24552
rect -3876 24535 -3874 24555
rect -3540 24535 -3538 24555
rect -3468 24535 -3466 24555
rect -3324 24535 -3322 24555
rect -3108 24535 -3106 24555
rect -3012 24535 -3010 24555
rect -2964 24535 -2962 24555
rect -2916 24535 -2914 24555
rect -2868 24535 -2866 24555
rect -2820 24535 -2818 24555
rect -2772 24535 -2770 24555
rect -2676 24535 -2674 24555
rect -2364 24535 -2362 24555
rect -2361 24552 -2347 24555
rect -2337 24555 2045 24559
rect -2337 24552 -2323 24555
rect -2316 24552 -2313 24555
rect -1980 24535 -1978 24555
rect -1812 24535 -1810 24555
rect -1572 24535 -1570 24555
rect -1476 24535 -1474 24555
rect -1356 24535 -1354 24555
rect -1260 24535 -1258 24555
rect -1236 24535 -1234 24555
rect -1140 24535 -1138 24555
rect -876 24535 -874 24555
rect -660 24535 -658 24555
rect -503 24550 -500 24555
rect -492 24550 -490 24555
rect -493 24536 -490 24550
rect -396 24552 -394 24555
rect -396 24535 -393 24552
rect -12 24535 -10 24555
rect 84 24535 86 24555
rect 156 24535 158 24555
rect 252 24535 254 24555
rect 348 24535 350 24555
rect 468 24535 470 24555
rect 492 24535 494 24555
rect 564 24535 566 24555
rect 588 24535 590 24555
rect 636 24535 638 24555
rect 660 24535 662 24555
rect 732 24535 734 24555
rect 948 24535 950 24555
rect 1044 24535 1046 24555
rect 1092 24535 1094 24555
rect 1140 24535 1142 24555
rect 1308 24535 1310 24555
rect 1356 24535 1358 24555
rect 1428 24535 1430 24555
rect 1561 24535 1619 24536
rect 1692 24535 1694 24555
rect 1860 24535 1862 24555
rect 1956 24535 1958 24555
rect 2031 24552 2045 24555
rect 2052 24555 9917 24559
rect 2052 24552 2069 24555
rect 2052 24535 2054 24552
rect 2148 24535 2150 24555
rect 2244 24535 2246 24555
rect 2460 24535 2462 24555
rect 2772 24535 2774 24555
rect 2868 24535 2870 24555
rect 2940 24535 2942 24555
rect 2988 24535 2990 24555
rect 3324 24535 3326 24555
rect 3396 24535 3398 24555
rect 3564 24535 3566 24555
rect 3660 24535 3662 24555
rect 3780 24535 3782 24555
rect 4092 24535 4094 24555
rect 4188 24535 4190 24555
rect 4308 24535 4310 24555
rect 4404 24535 4406 24555
rect 4500 24535 4502 24555
rect 4596 24535 4598 24555
rect 4692 24535 4694 24555
rect 4932 24535 4934 24555
rect 4980 24535 4982 24555
rect 5028 24535 5030 24555
rect 5124 24535 5126 24555
rect 5220 24535 5222 24555
rect 5388 24535 5390 24555
rect 5508 24535 5510 24555
rect 5532 24535 5534 24555
rect 5556 24535 5558 24555
rect 5628 24535 5630 24555
rect 5652 24535 5654 24555
rect 5748 24535 5750 24555
rect 5796 24535 5798 24555
rect 5844 24535 5846 24555
rect 5892 24535 5894 24555
rect 6276 24535 6278 24555
rect 6372 24535 6374 24555
rect 6420 24535 6422 24555
rect 6492 24535 6494 24555
rect 6516 24535 6518 24555
rect 6588 24535 6590 24555
rect 6612 24535 6614 24555
rect 6636 24535 6638 24555
rect 6684 24535 6686 24555
rect 6708 24535 6710 24555
rect 6780 24535 6782 24555
rect 6804 24535 6806 24555
rect 6900 24535 6902 24555
rect 6924 24536 6926 24555
rect 6913 24535 6947 24536
rect 7020 24535 7022 24555
rect 7164 24535 7166 24555
rect 7236 24535 7238 24555
rect 7284 24535 7286 24555
rect 7380 24535 7382 24555
rect 7404 24535 7406 24555
rect 7476 24535 7478 24555
rect 7500 24535 7502 24555
rect 7572 24535 7574 24555
rect 7644 24535 7646 24555
rect 7668 24535 7670 24555
rect 7908 24535 7910 24555
rect 8124 24535 8126 24555
rect 8220 24535 8222 24555
rect 8652 24535 8654 24555
rect 8700 24535 8702 24555
rect 8748 24535 8750 24555
rect 8796 24535 8798 24555
rect 8844 24535 8846 24555
rect 8868 24535 8870 24555
rect 9516 24535 9518 24555
rect 9660 24535 9662 24555
rect 9684 24535 9686 24555
rect 9756 24536 9758 24555
rect 9721 24535 9779 24536
rect 9780 24535 9782 24555
rect 9804 24535 9806 24555
rect 9903 24552 9917 24555
rect 9927 24555 22115 24559
rect 9927 24552 9941 24555
rect 9948 24552 9951 24555
rect 10044 24535 10046 24555
rect 10140 24535 10142 24555
rect 10236 24535 10238 24555
rect 10332 24535 10334 24555
rect 10380 24535 10382 24555
rect 10428 24535 10430 24555
rect 10524 24535 10526 24555
rect 10548 24535 10550 24555
rect 10620 24535 10622 24555
rect 10644 24535 10646 24555
rect 10716 24535 10718 24555
rect 10884 24535 10886 24555
rect 10956 24535 10958 24555
rect 11052 24535 11054 24555
rect 11100 24535 11102 24555
rect 11172 24535 11174 24555
rect 11220 24535 11222 24555
rect 11340 24535 11342 24555
rect 11436 24535 11438 24555
rect 11676 24535 11678 24555
rect 11724 24535 11726 24555
rect 11772 24535 11774 24555
rect 11796 24535 11798 24555
rect 12060 24535 12062 24555
rect 12276 24535 12278 24555
rect 12324 24535 12326 24555
rect 12372 24535 12374 24555
rect 12420 24535 12422 24555
rect 12433 24550 12436 24555
rect 12444 24550 12446 24555
rect 12443 24536 12446 24550
rect 12468 24535 12470 24555
rect 12540 24552 12542 24555
rect 12540 24535 12543 24552
rect 12564 24535 12566 24555
rect 12660 24535 12662 24555
rect 12756 24535 12758 24555
rect 12780 24535 12782 24555
rect 12828 24535 12830 24555
rect 12876 24535 12878 24555
rect 12972 24535 12974 24555
rect 13044 24535 13046 24555
rect 13068 24535 13070 24555
rect 13284 24535 13286 24555
rect 13332 24535 13334 24555
rect 13500 24535 13502 24555
rect 13572 24535 13574 24555
rect 13668 24535 13670 24555
rect 13716 24535 13718 24555
rect 13753 24550 13756 24555
rect 13764 24550 13766 24555
rect 13763 24536 13766 24550
rect 13860 24552 13862 24555
rect 13860 24535 13863 24552
rect 13956 24535 13958 24555
rect 14004 24535 14006 24555
rect 14100 24535 14102 24555
rect 14940 24535 14942 24555
rect 15036 24535 15038 24555
rect 15276 24535 15278 24555
rect 15361 24535 15419 24536
rect 15420 24535 15422 24555
rect 15564 24535 15566 24555
rect 15660 24535 15662 24555
rect 15708 24535 15710 24555
rect 15732 24535 15734 24555
rect 15756 24535 15758 24555
rect 15804 24535 15806 24555
rect 15828 24535 15830 24555
rect 15852 24535 15854 24555
rect 15948 24535 15950 24555
rect 15972 24535 15974 24555
rect 16044 24535 16046 24555
rect 16068 24535 16070 24555
rect 16164 24535 16166 24555
rect 16260 24535 16262 24555
rect 16332 24535 16334 24555
rect 16380 24535 16382 24555
rect 16476 24535 16478 24555
rect 16548 24535 16550 24555
rect 16572 24535 16574 24555
rect 16668 24535 16670 24555
rect 16764 24535 16766 24555
rect 16812 24535 16814 24555
rect 16884 24535 16886 24555
rect 16908 24535 16910 24555
rect 16980 24535 16982 24555
rect 17028 24535 17030 24555
rect 17124 24535 17126 24555
rect 17196 24535 17198 24555
rect 17220 24535 17222 24555
rect 17292 24535 17294 24555
rect 17316 24535 17318 24555
rect 17964 24535 17966 24555
rect 18060 24535 18062 24555
rect 18132 24535 18134 24555
rect 18228 24535 18230 24555
rect 18492 24535 18494 24555
rect 18540 24535 18542 24555
rect 18636 24535 18638 24555
rect 18732 24535 18734 24555
rect 18828 24535 18830 24555
rect 18924 24535 18926 24555
rect 18972 24535 18974 24555
rect 19020 24535 19022 24555
rect 19068 24535 19070 24555
rect 19140 24535 19142 24555
rect 19164 24535 19166 24555
rect 19236 24535 19238 24555
rect 19260 24535 19262 24555
rect 19788 24535 19790 24555
rect 19836 24535 19838 24555
rect 19860 24535 19862 24555
rect 19884 24535 19886 24555
rect 19956 24535 19958 24555
rect 19980 24535 19982 24555
rect 20004 24535 20006 24555
rect 20052 24535 20054 24555
rect 20076 24535 20078 24555
rect 20100 24535 20102 24555
rect 20172 24535 20174 24555
rect 20196 24535 20198 24555
rect 20292 24535 20294 24555
rect 20388 24535 20390 24555
rect 20412 24535 20414 24555
rect 20508 24535 20510 24555
rect 20532 24535 20534 24555
rect 20604 24535 20606 24555
rect 20628 24535 20630 24555
rect 20892 24535 20894 24555
rect 20964 24535 20966 24555
rect 20988 24535 20990 24555
rect 21108 24535 21110 24555
rect 21204 24535 21206 24555
rect 21300 24535 21302 24555
rect 21324 24535 21326 24555
rect 21444 24535 21446 24555
rect 21468 24535 21470 24555
rect 21564 24535 21566 24555
rect 21588 24535 21590 24555
rect 21684 24535 21686 24555
rect 21708 24535 21710 24555
rect 22068 24536 22070 24555
rect 22057 24535 22091 24536
rect -9753 24531 -4195 24535
rect -9753 24528 -9739 24531
rect -9647 24511 -9613 24512
rect -9540 24511 -9538 24531
rect -9444 24512 -9442 24531
rect -9348 24512 -9346 24531
rect -9479 24511 -9421 24512
rect -9359 24511 -9301 24512
rect -9228 24511 -9226 24531
rect -9108 24511 -9106 24531
rect -9012 24511 -9010 24531
rect -8916 24511 -8914 24531
rect -8628 24511 -8626 24531
rect -8532 24511 -8530 24531
rect -8436 24511 -8434 24531
rect -8340 24511 -8338 24531
rect -8124 24511 -8122 24531
rect -7764 24511 -7762 24531
rect -7356 24511 -7354 24531
rect -7308 24511 -7306 24531
rect -7140 24511 -7138 24531
rect -6852 24511 -6850 24531
rect -6732 24511 -6730 24531
rect -6516 24512 -6514 24531
rect -6551 24511 -6493 24512
rect -6348 24511 -6346 24531
rect -6252 24511 -6250 24531
rect -5892 24511 -5890 24531
rect -5436 24511 -5434 24531
rect -5340 24511 -5338 24531
rect -5196 24528 -5194 24531
rect -5196 24511 -5193 24528
rect -4751 24511 -4717 24512
rect -4716 24511 -4714 24531
rect -4500 24511 -4498 24531
rect -4284 24511 -4282 24531
rect -4209 24528 -4195 24531
rect -4185 24531 13829 24535
rect -4185 24528 -4171 24531
rect -4164 24528 -4161 24531
rect -3876 24511 -3874 24531
rect -3540 24511 -3538 24531
rect -3468 24511 -3466 24531
rect -3324 24511 -3322 24531
rect -3108 24511 -3106 24531
rect -3012 24511 -3010 24531
rect -2964 24511 -2962 24531
rect -2916 24511 -2914 24531
rect -2868 24511 -2866 24531
rect -2820 24511 -2818 24531
rect -2772 24511 -2770 24531
rect -2676 24511 -2674 24531
rect -2364 24511 -2362 24531
rect -1980 24511 -1978 24531
rect -1812 24512 -1810 24531
rect -1572 24512 -1570 24531
rect -1823 24511 -1789 24512
rect -1583 24511 -1501 24512
rect -1476 24511 -1474 24531
rect -1356 24511 -1354 24531
rect -1260 24511 -1258 24531
rect -1236 24511 -1234 24531
rect -1140 24511 -1138 24531
rect -876 24511 -874 24531
rect -660 24511 -658 24531
rect -417 24528 -403 24531
rect -396 24528 -393 24531
rect -201 24528 -187 24531
rect -12 24511 -10 24531
rect 49 24511 83 24512
rect 84 24511 86 24531
rect 156 24511 158 24531
rect 252 24511 254 24531
rect 348 24511 350 24531
rect 468 24511 470 24531
rect 492 24511 494 24531
rect 564 24511 566 24531
rect 588 24511 590 24531
rect 636 24511 638 24531
rect 660 24511 662 24531
rect 732 24511 734 24531
rect 948 24511 950 24531
rect 1044 24511 1046 24531
rect 1092 24511 1094 24531
rect 1140 24511 1142 24531
rect 1308 24511 1310 24531
rect 1356 24511 1358 24531
rect 1428 24511 1430 24531
rect 1561 24526 1564 24531
rect 1692 24528 1694 24531
rect 1571 24512 1574 24526
rect 1537 24511 1571 24512
rect 1572 24511 1574 24512
rect 1692 24511 1695 24528
rect 1860 24511 1862 24531
rect 1921 24511 1955 24512
rect 1956 24511 1958 24531
rect 2052 24511 2054 24531
rect 2148 24511 2150 24531
rect 2244 24511 2246 24531
rect 2460 24511 2462 24531
rect 2497 24511 2531 24512
rect 2772 24511 2774 24531
rect 2868 24511 2870 24531
rect 2940 24511 2942 24531
rect 2988 24511 2990 24531
rect 3324 24511 3326 24531
rect 3396 24512 3398 24531
rect 3385 24511 3419 24512
rect 3433 24511 3491 24512
rect 3564 24511 3566 24531
rect 3660 24511 3662 24531
rect 3780 24511 3782 24531
rect 4092 24511 4094 24531
rect 4188 24511 4190 24531
rect 4308 24511 4310 24531
rect 4404 24511 4406 24531
rect 4500 24511 4502 24531
rect 4596 24511 4598 24531
rect 4692 24511 4694 24531
rect 4932 24511 4934 24531
rect 4980 24511 4982 24531
rect 5028 24511 5030 24531
rect 5124 24511 5126 24531
rect 5220 24511 5222 24531
rect 5388 24511 5390 24531
rect 5508 24511 5510 24531
rect 5532 24511 5534 24531
rect 5556 24511 5558 24531
rect 5628 24511 5630 24531
rect 5652 24511 5654 24531
rect 5748 24511 5750 24531
rect 5796 24511 5798 24531
rect 5844 24511 5846 24531
rect 5892 24511 5894 24531
rect 6276 24511 6278 24531
rect 6372 24511 6374 24531
rect 6420 24511 6422 24531
rect 6492 24511 6494 24531
rect 6516 24511 6518 24531
rect 6588 24511 6590 24531
rect 6612 24511 6614 24531
rect 6636 24511 6638 24531
rect 6684 24511 6686 24531
rect 6708 24511 6710 24531
rect 6780 24511 6782 24531
rect 6804 24511 6806 24531
rect 6900 24511 6902 24531
rect 6913 24526 6916 24531
rect 6924 24526 6926 24531
rect 6923 24512 6926 24526
rect 7020 24528 7022 24531
rect 7020 24511 7023 24528
rect 7164 24511 7166 24531
rect 7236 24511 7238 24531
rect 7284 24511 7286 24531
rect 7380 24511 7382 24531
rect 7404 24511 7406 24531
rect 7476 24511 7478 24531
rect 7500 24511 7502 24531
rect 7572 24511 7574 24531
rect 7644 24511 7646 24531
rect 7668 24511 7670 24531
rect 7908 24511 7910 24531
rect 8124 24511 8126 24531
rect 8220 24511 8222 24531
rect 8652 24511 8654 24531
rect 8700 24511 8702 24531
rect 8748 24511 8750 24531
rect 8796 24511 8798 24531
rect 8844 24511 8846 24531
rect 8868 24511 8870 24531
rect 9516 24511 9518 24531
rect 9660 24511 9662 24531
rect 9684 24511 9686 24531
rect 9745 24526 9748 24531
rect 9756 24526 9758 24531
rect 9755 24512 9758 24526
rect 9780 24511 9782 24531
rect 9804 24511 9806 24531
rect 9828 24511 9831 24528
rect 10044 24511 10046 24531
rect 10140 24511 10142 24531
rect 10236 24511 10238 24531
rect 10332 24511 10334 24531
rect 10380 24511 10382 24531
rect 10428 24511 10430 24531
rect 10524 24511 10526 24531
rect 10548 24511 10550 24531
rect 10620 24511 10622 24531
rect 10644 24511 10646 24531
rect 10716 24511 10718 24531
rect 10884 24511 10886 24531
rect 10956 24511 10958 24531
rect 11052 24511 11054 24531
rect 11100 24511 11102 24531
rect 11172 24511 11174 24531
rect 11220 24511 11222 24531
rect 11340 24511 11342 24531
rect 11436 24511 11438 24531
rect 11676 24511 11678 24531
rect 11724 24511 11726 24531
rect 11772 24511 11774 24531
rect 11796 24511 11798 24531
rect 12060 24511 12062 24531
rect 12276 24511 12278 24531
rect 12324 24511 12326 24531
rect 12372 24511 12374 24531
rect 12420 24511 12422 24531
rect 12468 24511 12470 24531
rect 12519 24528 12533 24531
rect 12540 24528 12543 24531
rect 12564 24511 12566 24531
rect 12660 24512 12662 24531
rect 12649 24511 12683 24512
rect 12756 24511 12758 24531
rect 12780 24511 12782 24531
rect 12828 24511 12830 24531
rect 12876 24511 12878 24531
rect 12972 24511 12974 24531
rect 13044 24511 13046 24531
rect 13068 24511 13070 24531
rect 13284 24511 13286 24531
rect 13332 24511 13334 24531
rect 13500 24511 13502 24531
rect 13572 24511 13574 24531
rect 13668 24511 13670 24531
rect 13716 24511 13718 24531
rect 13815 24528 13829 24531
rect 13839 24531 22091 24535
rect 13839 24528 13853 24531
rect 13860 24528 13863 24531
rect 13956 24511 13958 24531
rect 14004 24511 14006 24531
rect 14100 24511 14102 24531
rect 14940 24511 14942 24531
rect 15036 24511 15038 24531
rect 15276 24511 15278 24531
rect 15361 24526 15364 24531
rect 15371 24512 15374 24526
rect 15372 24511 15374 24512
rect 15420 24511 15422 24531
rect 15468 24511 15471 24528
rect 15564 24511 15566 24531
rect 15660 24511 15662 24531
rect 15708 24511 15710 24531
rect 15732 24511 15734 24531
rect 15756 24511 15758 24531
rect 15804 24511 15806 24531
rect 15828 24511 15830 24531
rect 15852 24511 15854 24531
rect 15948 24511 15950 24531
rect 15972 24511 15974 24531
rect 16044 24511 16046 24531
rect 16068 24511 16070 24531
rect 16164 24511 16166 24531
rect 16260 24511 16262 24531
rect 16332 24511 16334 24531
rect 16380 24511 16382 24531
rect 16476 24511 16478 24531
rect 16548 24511 16550 24531
rect 16572 24511 16574 24531
rect 16668 24511 16670 24531
rect 16764 24511 16766 24531
rect 16812 24511 16814 24531
rect 16884 24511 16886 24531
rect 16908 24511 16910 24531
rect 16980 24512 16982 24531
rect 16969 24511 17003 24512
rect 17028 24511 17030 24531
rect 17124 24511 17126 24531
rect 17196 24511 17198 24531
rect 17220 24511 17222 24531
rect 17292 24511 17294 24531
rect 17316 24511 17318 24531
rect 17964 24511 17966 24531
rect 18060 24511 18062 24531
rect 18132 24511 18134 24531
rect 18228 24511 18230 24531
rect 18492 24511 18494 24531
rect 18540 24511 18542 24531
rect 18636 24511 18638 24531
rect 18732 24511 18734 24531
rect 18828 24511 18830 24531
rect 18924 24511 18926 24531
rect 18972 24511 18974 24531
rect 19020 24511 19022 24531
rect 19068 24511 19070 24531
rect 19140 24511 19142 24531
rect 19164 24511 19166 24531
rect 19236 24511 19238 24531
rect 19260 24511 19262 24531
rect 19788 24511 19790 24531
rect 19836 24511 19838 24531
rect 19860 24511 19862 24531
rect 19884 24511 19886 24531
rect 19956 24511 19958 24531
rect 19980 24511 19982 24531
rect 20004 24511 20006 24531
rect 20052 24511 20054 24531
rect 20076 24511 20078 24531
rect 20100 24511 20102 24531
rect 20172 24511 20174 24531
rect 20196 24511 20198 24531
rect 20292 24511 20294 24531
rect 20388 24511 20390 24531
rect 20412 24511 20414 24531
rect 20508 24511 20510 24531
rect 20532 24511 20534 24531
rect 20604 24511 20606 24531
rect 20628 24511 20630 24531
rect 20892 24511 20894 24531
rect 20964 24511 20966 24531
rect 20988 24511 20990 24531
rect 21108 24511 21110 24531
rect 21204 24511 21206 24531
rect 21300 24511 21302 24531
rect 21324 24511 21326 24531
rect 21444 24511 21446 24531
rect 21468 24511 21470 24531
rect 21564 24511 21566 24531
rect 21588 24511 21590 24531
rect 21684 24511 21686 24531
rect 21708 24511 21710 24531
rect 22057 24526 22060 24531
rect 22068 24526 22070 24531
rect 22067 24512 22070 24526
rect 22033 24511 22067 24512
rect -9647 24507 1661 24511
rect -9540 24504 -9538 24507
rect -9540 24488 -9537 24504
rect -9455 24502 -9452 24507
rect -9444 24502 -9442 24507
rect -9359 24502 -9356 24507
rect -9348 24504 -9346 24507
rect -9228 24504 -9226 24507
rect -9348 24502 -9345 24504
rect -9445 24488 -9442 24502
rect -9349 24488 -9345 24502
rect -9228 24488 -9225 24504
rect -9551 24487 -9517 24488
rect -9503 24487 -9469 24488
rect -9551 24483 -9469 24487
rect -9287 24483 -9259 24488
rect -9239 24487 -9181 24488
rect -9108 24487 -9106 24507
rect -9012 24487 -9010 24507
rect -8916 24487 -8914 24507
rect -8628 24487 -8626 24507
rect -8532 24487 -8530 24507
rect -8436 24487 -8434 24507
rect -8340 24487 -8338 24507
rect -8124 24487 -8122 24507
rect -7764 24487 -7762 24507
rect -7356 24487 -7354 24507
rect -7308 24487 -7306 24507
rect -7140 24487 -7138 24507
rect -6852 24487 -6850 24507
rect -6732 24487 -6730 24507
rect -6527 24502 -6524 24507
rect -6516 24502 -6514 24507
rect -6517 24488 -6514 24502
rect -6444 24487 -6441 24504
rect -6348 24487 -6346 24507
rect -6252 24487 -6250 24507
rect -5892 24487 -5890 24507
rect -5673 24504 -5659 24507
rect -5436 24487 -5434 24507
rect -5340 24487 -5338 24507
rect -5217 24504 -5203 24507
rect -5196 24504 -5193 24507
rect -4716 24487 -4714 24507
rect -4500 24487 -4498 24507
rect -4284 24487 -4282 24507
rect -3876 24487 -3874 24507
rect -3540 24487 -3538 24507
rect -3468 24487 -3466 24507
rect -3324 24487 -3322 24507
rect -3108 24487 -3106 24507
rect -3012 24487 -3010 24507
rect -2964 24487 -2962 24507
rect -2916 24487 -2914 24507
rect -2868 24487 -2866 24507
rect -2820 24487 -2818 24507
rect -2772 24487 -2770 24507
rect -2676 24487 -2674 24507
rect -2364 24487 -2362 24507
rect -1980 24487 -1978 24507
rect -1823 24502 -1820 24507
rect -1812 24502 -1810 24507
rect -1583 24502 -1580 24507
rect -1572 24502 -1570 24507
rect -1813 24488 -1810 24502
rect -1573 24488 -1570 24502
rect -1476 24504 -1474 24507
rect -1476 24487 -1473 24504
rect -1452 24487 -1449 24504
rect -1356 24487 -1354 24507
rect -1260 24487 -1258 24507
rect -1236 24487 -1234 24507
rect -1140 24487 -1138 24507
rect -876 24487 -874 24507
rect -791 24487 -733 24488
rect -660 24487 -658 24507
rect -575 24487 -517 24488
rect -12 24487 -10 24507
rect 84 24487 86 24507
rect 156 24504 158 24507
rect 156 24487 159 24504
rect 252 24487 254 24507
rect 348 24487 350 24507
rect 468 24487 470 24507
rect 492 24487 494 24507
rect 564 24487 566 24507
rect 588 24487 590 24507
rect 636 24487 638 24507
rect 660 24487 662 24507
rect 732 24487 734 24507
rect 913 24487 947 24488
rect 948 24487 950 24507
rect 1044 24487 1046 24507
rect 1092 24487 1094 24507
rect 1140 24487 1142 24507
rect 1308 24487 1310 24507
rect 1356 24487 1358 24507
rect 1428 24487 1430 24507
rect 1572 24487 1574 24507
rect 1647 24504 1661 24507
rect 1671 24507 9821 24511
rect 1671 24504 1685 24507
rect 1692 24504 1695 24507
rect 1860 24487 1862 24507
rect 1956 24487 1958 24507
rect 2052 24487 2054 24507
rect 2148 24487 2150 24507
rect 2244 24487 2246 24507
rect 2460 24487 2462 24507
rect 2772 24487 2774 24507
rect 2868 24487 2870 24507
rect 2940 24487 2942 24507
rect 2988 24487 2990 24507
rect 3324 24487 3326 24507
rect 3385 24502 3388 24507
rect 3396 24502 3398 24507
rect 3564 24504 3566 24507
rect 3395 24488 3398 24502
rect 3481 24494 3485 24502
rect 3471 24488 3481 24494
rect 3540 24487 3543 24504
rect 3564 24487 3567 24504
rect 3660 24487 3662 24507
rect 3780 24487 3782 24507
rect 4092 24487 4094 24507
rect 4188 24487 4190 24507
rect 4308 24487 4310 24507
rect 4404 24487 4406 24507
rect 4500 24487 4502 24507
rect 4596 24487 4598 24507
rect 4692 24487 4694 24507
rect 4932 24487 4934 24507
rect 4980 24487 4982 24507
rect 5028 24487 5030 24507
rect 5124 24487 5126 24507
rect 5220 24487 5222 24507
rect 5388 24487 5390 24507
rect 5425 24487 5459 24488
rect 5508 24487 5510 24507
rect 5532 24488 5534 24507
rect 5521 24487 5555 24488
rect 5556 24487 5558 24507
rect 5628 24487 5630 24507
rect 5652 24487 5654 24507
rect 5748 24487 5750 24507
rect 5796 24487 5798 24507
rect 5844 24487 5846 24507
rect 5892 24487 5894 24507
rect 6276 24487 6278 24507
rect 6372 24487 6374 24507
rect 6420 24487 6422 24507
rect 6492 24487 6494 24507
rect 6516 24487 6518 24507
rect 6588 24487 6590 24507
rect 6612 24487 6614 24507
rect 6636 24487 6638 24507
rect 6684 24487 6686 24507
rect 6708 24487 6710 24507
rect 6780 24487 6782 24507
rect 6804 24487 6806 24507
rect 6900 24487 6902 24507
rect 6999 24504 7013 24507
rect 7020 24504 7023 24507
rect 7164 24487 7166 24507
rect 7236 24487 7238 24507
rect 7284 24487 7286 24507
rect 7380 24487 7382 24507
rect 7404 24487 7406 24507
rect 7476 24487 7478 24507
rect 7500 24487 7502 24507
rect 7572 24487 7574 24507
rect 7644 24487 7646 24507
rect 7668 24487 7670 24507
rect 7908 24487 7910 24507
rect 8124 24487 8126 24507
rect 8220 24487 8222 24507
rect 8652 24487 8654 24507
rect 8700 24487 8702 24507
rect 8748 24487 8750 24507
rect 8796 24487 8798 24507
rect 8844 24487 8846 24507
rect 8868 24487 8870 24507
rect 9516 24487 9518 24507
rect 9660 24487 9662 24507
rect 9684 24487 9686 24507
rect 9780 24487 9782 24507
rect 9804 24487 9806 24507
rect 9807 24504 9821 24507
rect 9828 24507 15461 24511
rect 9828 24504 9845 24507
rect 9828 24487 9830 24504
rect 10044 24487 10046 24507
rect 10140 24487 10142 24507
rect 10236 24487 10238 24507
rect 10332 24487 10334 24507
rect 10380 24487 10382 24507
rect 10428 24487 10430 24507
rect 10524 24487 10526 24507
rect 10548 24487 10550 24507
rect 10620 24487 10622 24507
rect 10644 24487 10646 24507
rect 10716 24487 10718 24507
rect 10884 24487 10886 24507
rect 10956 24487 10958 24507
rect 11052 24487 11054 24507
rect 11100 24487 11102 24507
rect 11172 24487 11174 24507
rect 11220 24487 11222 24507
rect 11340 24487 11342 24507
rect 11436 24487 11438 24507
rect 11676 24487 11678 24507
rect 11724 24487 11726 24507
rect 11772 24487 11774 24507
rect 11796 24487 11798 24507
rect 12060 24487 12062 24507
rect 12276 24487 12278 24507
rect 12324 24487 12326 24507
rect 12372 24487 12374 24507
rect 12420 24487 12422 24507
rect 12468 24487 12470 24507
rect 12564 24487 12566 24507
rect 12649 24502 12652 24507
rect 12660 24502 12662 24507
rect 12659 24488 12662 24502
rect 12756 24504 12758 24507
rect 12756 24487 12759 24504
rect 12780 24487 12782 24507
rect 12828 24487 12830 24507
rect 12876 24487 12878 24507
rect 12972 24487 12974 24507
rect 13044 24487 13046 24507
rect 13068 24487 13070 24507
rect 13284 24487 13286 24507
rect 13332 24487 13334 24507
rect 13500 24487 13502 24507
rect 13572 24487 13574 24507
rect 13668 24487 13670 24507
rect 13716 24487 13718 24507
rect 13956 24487 13958 24507
rect 14004 24487 14006 24507
rect 14100 24487 14102 24507
rect 14940 24487 14942 24507
rect 15036 24487 15038 24507
rect 15276 24487 15278 24507
rect 15372 24487 15374 24507
rect 15420 24487 15422 24507
rect 15447 24504 15461 24507
rect 15468 24507 22067 24511
rect 15468 24504 15485 24507
rect 15468 24487 15470 24504
rect 15564 24487 15566 24507
rect 15660 24487 15662 24507
rect 15708 24487 15710 24507
rect 15732 24487 15734 24507
rect 15756 24487 15758 24507
rect 15804 24487 15806 24507
rect 15828 24487 15830 24507
rect 15852 24487 15854 24507
rect 15948 24487 15950 24507
rect 15972 24487 15974 24507
rect 16044 24487 16046 24507
rect 16068 24487 16070 24507
rect 16164 24487 16166 24507
rect 16260 24487 16262 24507
rect 16332 24487 16334 24507
rect 16380 24487 16382 24507
rect 16476 24487 16478 24507
rect 16548 24487 16550 24507
rect 16572 24487 16574 24507
rect 16668 24487 16670 24507
rect 16764 24487 16766 24507
rect 16812 24487 16814 24507
rect 16884 24487 16886 24507
rect 16908 24487 16910 24507
rect 16969 24502 16972 24507
rect 16980 24502 16982 24507
rect 16979 24488 16982 24502
rect 17028 24487 17030 24507
rect 17124 24487 17126 24507
rect 17196 24487 17198 24507
rect 17220 24487 17222 24507
rect 17292 24487 17294 24507
rect 17316 24487 17318 24507
rect 17964 24487 17966 24507
rect 18060 24487 18062 24507
rect 18132 24487 18134 24507
rect 18228 24487 18230 24507
rect 18492 24487 18494 24507
rect 18540 24487 18542 24507
rect 18636 24487 18638 24507
rect 18732 24487 18734 24507
rect 18828 24487 18830 24507
rect 18924 24487 18926 24507
rect 18972 24487 18974 24507
rect 19020 24487 19022 24507
rect 19068 24487 19070 24507
rect 19140 24487 19142 24507
rect 19164 24487 19166 24507
rect 19236 24487 19238 24507
rect 19260 24487 19262 24507
rect 19788 24487 19790 24507
rect 19836 24487 19838 24507
rect 19860 24487 19862 24507
rect 19884 24487 19886 24507
rect 19956 24487 19958 24507
rect 19980 24487 19982 24507
rect 20004 24487 20006 24507
rect 20052 24487 20054 24507
rect 20076 24487 20078 24507
rect 20100 24487 20102 24507
rect 20172 24487 20174 24507
rect 20196 24487 20198 24507
rect 20292 24487 20294 24507
rect 20388 24487 20390 24507
rect 20412 24487 20414 24507
rect 20508 24487 20510 24507
rect 20532 24487 20534 24507
rect 20604 24487 20606 24507
rect 20628 24487 20630 24507
rect 20892 24487 20894 24507
rect 20964 24487 20966 24507
rect 20988 24487 20990 24507
rect 21108 24487 21110 24507
rect 21204 24487 21206 24507
rect 21300 24487 21302 24507
rect 21324 24487 21326 24507
rect 21444 24487 21446 24507
rect 21468 24487 21470 24507
rect 21564 24487 21566 24507
rect 21588 24487 21590 24507
rect 21684 24487 21686 24507
rect 21708 24487 21710 24507
rect 21961 24487 21995 24488
rect -9551 24480 -9547 24483
rect -9540 24480 -9537 24483
rect -9273 24480 -9259 24483
rect -9249 24483 -6451 24487
rect -9249 24480 -9235 24483
rect -9228 24480 -9225 24483
rect -9108 24480 -9106 24483
rect -9191 24470 -9187 24478
rect -9201 24464 -9191 24470
rect -9108 24464 -9105 24480
rect -9012 24464 -9010 24483
rect -8916 24464 -8914 24483
rect -9119 24463 -9085 24464
rect -9047 24463 -8989 24464
rect -8927 24463 -8893 24464
rect -9119 24459 -8893 24463
rect -8879 24463 -8845 24464
rect -8628 24463 -8626 24483
rect -8532 24463 -8530 24483
rect -8436 24463 -8434 24483
rect -8340 24463 -8338 24483
rect -8124 24463 -8122 24483
rect -7764 24463 -7762 24483
rect -7356 24463 -7354 24483
rect -7308 24463 -7306 24483
rect -7140 24463 -7138 24483
rect -6852 24463 -6850 24483
rect -6732 24463 -6730 24483
rect -6465 24480 -6451 24483
rect -6444 24483 -1459 24487
rect -6444 24480 -6427 24483
rect -6444 24463 -6442 24480
rect -6348 24463 -6346 24483
rect -6252 24463 -6250 24483
rect -5892 24463 -5890 24483
rect -5436 24463 -5434 24483
rect -5340 24463 -5338 24483
rect -4716 24463 -4714 24483
rect -4665 24480 -4651 24483
rect -4500 24463 -4498 24483
rect -4284 24463 -4282 24483
rect -3876 24463 -3874 24483
rect -3540 24463 -3538 24483
rect -3468 24463 -3466 24483
rect -3324 24463 -3322 24483
rect -3108 24463 -3106 24483
rect -3012 24463 -3010 24483
rect -2964 24463 -2962 24483
rect -2916 24463 -2914 24483
rect -2868 24463 -2866 24483
rect -2820 24463 -2818 24483
rect -2772 24463 -2770 24483
rect -2676 24463 -2674 24483
rect -2364 24463 -2362 24483
rect -1980 24464 -1978 24483
rect -1737 24480 -1723 24483
rect -1497 24480 -1483 24483
rect -1476 24480 -1459 24483
rect -1452 24483 3533 24487
rect -1452 24480 -1435 24483
rect -2015 24463 -1957 24464
rect -1452 24463 -1450 24480
rect -1356 24463 -1354 24483
rect -1260 24463 -1258 24483
rect -1236 24463 -1234 24483
rect -1140 24463 -1138 24483
rect -876 24463 -874 24483
rect -791 24478 -788 24483
rect -660 24480 -658 24483
rect -781 24464 -778 24478
rect -780 24463 -778 24464
rect -660 24463 -657 24480
rect -575 24478 -572 24483
rect -565 24464 -562 24478
rect -564 24463 -562 24464
rect -468 24463 -465 24480
rect -12 24463 -10 24483
rect 84 24463 86 24483
rect 135 24480 149 24483
rect 156 24480 159 24483
rect 252 24463 254 24483
rect 348 24463 350 24483
rect 468 24463 470 24483
rect 492 24463 494 24483
rect 564 24463 566 24483
rect 588 24463 590 24483
rect 636 24463 638 24483
rect 660 24463 662 24483
rect 732 24463 734 24483
rect 948 24463 950 24483
rect 1044 24463 1046 24483
rect 1092 24463 1094 24483
rect 1140 24463 1142 24483
rect 1308 24463 1310 24483
rect 1356 24463 1358 24483
rect 1428 24463 1430 24483
rect 1572 24463 1574 24483
rect 1623 24480 1637 24483
rect 1860 24463 1862 24483
rect 1956 24463 1958 24483
rect 2007 24480 2021 24483
rect 2052 24463 2054 24483
rect 2148 24463 2150 24483
rect 2244 24463 2246 24483
rect 2460 24463 2462 24483
rect 2583 24480 2597 24483
rect 2772 24463 2774 24483
rect 2868 24463 2870 24483
rect 2940 24463 2942 24483
rect 2988 24463 2990 24483
rect 3324 24463 3326 24483
rect 3471 24480 3485 24483
rect 3519 24480 3533 24483
rect 3540 24483 21995 24487
rect 3540 24480 3557 24483
rect 3564 24480 3567 24483
rect 3540 24463 3542 24480
rect 3660 24463 3662 24483
rect 3780 24463 3782 24483
rect 4092 24463 4094 24483
rect 4188 24463 4190 24483
rect 4308 24463 4310 24483
rect 4404 24463 4406 24483
rect 4500 24463 4502 24483
rect 4596 24463 4598 24483
rect 4692 24463 4694 24483
rect 4932 24463 4934 24483
rect 4980 24463 4982 24483
rect 5028 24463 5030 24483
rect 5124 24463 5126 24483
rect 5220 24463 5222 24483
rect 5388 24463 5390 24483
rect 5508 24463 5510 24483
rect 5521 24478 5524 24483
rect 5532 24480 5534 24483
rect 5532 24478 5535 24480
rect 5531 24464 5535 24478
rect 5556 24463 5558 24483
rect 5628 24480 5630 24483
rect 5628 24463 5631 24480
rect 5652 24463 5654 24483
rect 5748 24463 5750 24483
rect 5796 24463 5798 24483
rect 5844 24463 5846 24483
rect 5892 24463 5894 24483
rect 6276 24463 6278 24483
rect 6372 24463 6374 24483
rect 6420 24463 6422 24483
rect 6492 24463 6494 24483
rect 6516 24463 6518 24483
rect 6588 24463 6590 24483
rect 6612 24463 6614 24483
rect 6636 24463 6638 24483
rect 6684 24463 6686 24483
rect 6708 24463 6710 24483
rect 6780 24464 6782 24483
rect 6745 24463 6803 24464
rect 6804 24463 6806 24483
rect 6900 24463 6902 24483
rect 7164 24463 7166 24483
rect 7236 24463 7238 24483
rect 7284 24463 7286 24483
rect 7380 24463 7382 24483
rect 7404 24463 7406 24483
rect 7476 24463 7478 24483
rect 7500 24463 7502 24483
rect 7572 24463 7574 24483
rect 7644 24463 7646 24483
rect 7668 24463 7670 24483
rect 7908 24463 7910 24483
rect 8124 24463 8126 24483
rect 8220 24463 8222 24483
rect 8652 24463 8654 24483
rect 8700 24463 8702 24483
rect 8748 24463 8750 24483
rect 8796 24463 8798 24483
rect 8844 24463 8846 24483
rect 8868 24463 8870 24483
rect 9516 24463 9518 24483
rect 9660 24463 9662 24483
rect 9684 24463 9686 24483
rect 9780 24463 9782 24483
rect 9804 24463 9806 24483
rect 9828 24463 9830 24483
rect 10044 24463 10046 24483
rect 10140 24463 10142 24483
rect 10236 24463 10238 24483
rect 10332 24463 10334 24483
rect 10380 24463 10382 24483
rect 10428 24463 10430 24483
rect 10524 24463 10526 24483
rect 10548 24463 10550 24483
rect 10620 24463 10622 24483
rect 10644 24463 10646 24483
rect 10716 24463 10718 24483
rect 10884 24463 10886 24483
rect 10956 24463 10958 24483
rect 11052 24463 11054 24483
rect 11100 24463 11102 24483
rect 11172 24463 11174 24483
rect 11220 24463 11222 24483
rect 11340 24463 11342 24483
rect 11436 24463 11438 24483
rect 11676 24463 11678 24483
rect 11724 24463 11726 24483
rect 11772 24463 11774 24483
rect 11796 24463 11798 24483
rect 12060 24463 12062 24483
rect 12276 24463 12278 24483
rect 12324 24463 12326 24483
rect 12372 24463 12374 24483
rect 12420 24463 12422 24483
rect 12468 24463 12470 24483
rect 12564 24463 12566 24483
rect 12735 24480 12749 24483
rect 12756 24480 12759 24483
rect 12780 24463 12782 24483
rect 12828 24463 12830 24483
rect 12876 24463 12878 24483
rect 12972 24463 12974 24483
rect 13044 24463 13046 24483
rect 13068 24463 13070 24483
rect 13284 24463 13286 24483
rect 13332 24463 13334 24483
rect 13500 24463 13502 24483
rect 13572 24463 13574 24483
rect 13668 24463 13670 24483
rect 13716 24463 13718 24483
rect 13825 24463 13883 24464
rect 13956 24463 13958 24483
rect 14004 24463 14006 24483
rect 14100 24463 14102 24483
rect 14940 24463 14942 24483
rect 15036 24463 15038 24483
rect 15276 24463 15278 24483
rect 15372 24463 15374 24483
rect 15420 24463 15422 24483
rect 15468 24463 15470 24483
rect 15564 24463 15566 24483
rect 15660 24463 15662 24483
rect 15708 24463 15710 24483
rect 15732 24463 15734 24483
rect 15756 24463 15758 24483
rect 15804 24463 15806 24483
rect 15828 24463 15830 24483
rect 15852 24463 15854 24483
rect 15948 24463 15950 24483
rect 15972 24463 15974 24483
rect 16044 24463 16046 24483
rect 16068 24463 16070 24483
rect 16164 24463 16166 24483
rect 16260 24463 16262 24483
rect 16332 24463 16334 24483
rect 16380 24463 16382 24483
rect 16476 24463 16478 24483
rect 16548 24463 16550 24483
rect 16572 24463 16574 24483
rect 16668 24463 16670 24483
rect 16764 24463 16766 24483
rect 16812 24463 16814 24483
rect 16884 24463 16886 24483
rect 16908 24463 16910 24483
rect 17028 24463 17030 24483
rect 17055 24480 17069 24483
rect 17124 24463 17126 24483
rect 17196 24463 17198 24483
rect 17220 24463 17222 24483
rect 17292 24463 17294 24483
rect 17316 24463 17318 24483
rect 17964 24463 17966 24483
rect 18060 24463 18062 24483
rect 18132 24463 18134 24483
rect 18228 24463 18230 24483
rect 18492 24463 18494 24483
rect 18540 24463 18542 24483
rect 18636 24463 18638 24483
rect 18732 24463 18734 24483
rect 18828 24463 18830 24483
rect 18924 24463 18926 24483
rect 18972 24463 18974 24483
rect 19020 24463 19022 24483
rect 19068 24463 19070 24483
rect 19140 24463 19142 24483
rect 19164 24463 19166 24483
rect 19236 24463 19238 24483
rect 19260 24463 19262 24483
rect 19788 24463 19790 24483
rect 19836 24463 19838 24483
rect 19860 24463 19862 24483
rect 19884 24463 19886 24483
rect 19956 24463 19958 24483
rect 19980 24463 19982 24483
rect 20004 24463 20006 24483
rect 20052 24463 20054 24483
rect 20076 24463 20078 24483
rect 20100 24463 20102 24483
rect 20172 24463 20174 24483
rect 20196 24463 20198 24483
rect 20292 24463 20294 24483
rect 20388 24463 20390 24483
rect 20412 24463 20414 24483
rect 20508 24463 20510 24483
rect 20532 24463 20534 24483
rect 20604 24463 20606 24483
rect 20628 24463 20630 24483
rect 20892 24463 20894 24483
rect 20964 24463 20966 24483
rect 20988 24463 20990 24483
rect 21108 24463 21110 24483
rect 21204 24463 21206 24483
rect 21300 24463 21302 24483
rect 21324 24463 21326 24483
rect 21444 24463 21446 24483
rect 21468 24463 21470 24483
rect 21564 24463 21566 24483
rect 21588 24463 21590 24483
rect 21684 24463 21686 24483
rect 21708 24463 21710 24483
rect 21913 24463 21947 24464
rect -8879 24459 -691 24463
rect -9119 24456 -9115 24459
rect -9108 24456 -9105 24459
rect -9023 24454 -9020 24459
rect -9012 24456 -9010 24459
rect -9012 24454 -9009 24456
rect -8927 24454 -8924 24459
rect -8916 24456 -8914 24459
rect -8916 24454 -8913 24456
rect -9023 24446 -9019 24454
rect -9033 24440 -9023 24446
rect -9013 24440 -9009 24454
rect -8917 24440 -8913 24454
rect -8735 24439 -8701 24440
rect -8628 24439 -8626 24459
rect -8532 24439 -8530 24459
rect -8436 24439 -8434 24459
rect -8340 24439 -8338 24459
rect -8124 24439 -8122 24459
rect -7764 24439 -7762 24459
rect -7356 24439 -7354 24459
rect -7308 24439 -7306 24459
rect -7140 24439 -7138 24459
rect -6959 24439 -6877 24440
rect -6852 24439 -6850 24459
rect -6732 24439 -6730 24459
rect -6444 24439 -6442 24459
rect -6348 24439 -6346 24459
rect -6252 24439 -6250 24459
rect -5892 24439 -5890 24459
rect -5567 24439 -5509 24440
rect -5436 24439 -5434 24459
rect -5340 24439 -5338 24459
rect -4716 24439 -4714 24459
rect -4500 24439 -4498 24459
rect -4284 24439 -4282 24459
rect -3876 24439 -3874 24459
rect -3540 24439 -3538 24459
rect -3468 24439 -3466 24459
rect -3324 24439 -3322 24459
rect -3108 24439 -3106 24459
rect -3012 24439 -3010 24459
rect -2964 24439 -2962 24459
rect -2916 24439 -2914 24459
rect -2868 24439 -2866 24459
rect -2820 24440 -2818 24459
rect -2831 24439 -2797 24440
rect -2772 24439 -2770 24459
rect -2676 24440 -2674 24459
rect -2687 24439 -2653 24440
rect -2364 24439 -2362 24459
rect -1991 24454 -1988 24459
rect -1980 24454 -1978 24459
rect -1981 24440 -1978 24454
rect -1908 24439 -1905 24456
rect -1452 24439 -1450 24459
rect -1356 24439 -1354 24459
rect -1260 24439 -1258 24459
rect -1236 24439 -1234 24459
rect -1140 24439 -1138 24459
rect -876 24439 -874 24459
rect -780 24439 -778 24459
rect -705 24456 -691 24459
rect -681 24459 -475 24463
rect -681 24456 -667 24459
rect -660 24456 -657 24459
rect -564 24439 -562 24459
rect -489 24456 -475 24459
rect -468 24459 21947 24463
rect -468 24456 -451 24459
rect -468 24439 -466 24456
rect -12 24439 -10 24459
rect 84 24439 86 24459
rect 121 24439 155 24440
rect 252 24439 254 24459
rect 348 24439 350 24459
rect 468 24439 470 24459
rect 492 24439 494 24459
rect 564 24439 566 24459
rect 588 24439 590 24459
rect 636 24439 638 24459
rect 660 24439 662 24459
rect 732 24439 734 24459
rect 948 24439 950 24459
rect 999 24456 1013 24459
rect 1044 24439 1046 24459
rect 1092 24439 1094 24459
rect 1140 24439 1142 24459
rect 1308 24439 1310 24459
rect 1356 24439 1358 24459
rect 1428 24439 1430 24459
rect 1572 24439 1574 24459
rect 1860 24439 1862 24459
rect 1956 24439 1958 24459
rect 2052 24439 2054 24459
rect 2148 24439 2150 24459
rect 2244 24439 2246 24459
rect 2460 24439 2462 24459
rect 2772 24439 2774 24459
rect 2868 24439 2870 24459
rect 2940 24439 2942 24459
rect 2988 24439 2990 24459
rect 3324 24439 3326 24459
rect 3540 24439 3542 24459
rect 3660 24439 3662 24459
rect 3780 24439 3782 24459
rect 4092 24439 4094 24459
rect 4188 24439 4190 24459
rect 4308 24439 4310 24459
rect 4404 24439 4406 24459
rect 4500 24439 4502 24459
rect 4596 24439 4598 24459
rect 4692 24439 4694 24459
rect 4932 24439 4934 24459
rect 4980 24439 4982 24459
rect 5028 24439 5030 24459
rect 5124 24439 5126 24459
rect 5220 24439 5222 24459
rect 5388 24439 5390 24459
rect 5508 24439 5510 24459
rect 5511 24456 5525 24459
rect 5556 24439 5558 24459
rect 5607 24456 5621 24459
rect 5628 24456 5631 24459
rect 5652 24439 5654 24459
rect 5748 24439 5750 24459
rect 5796 24439 5798 24459
rect 5844 24439 5846 24459
rect 5892 24439 5894 24459
rect 6276 24439 6278 24459
rect 6372 24439 6374 24459
rect 6420 24439 6422 24459
rect 6492 24439 6494 24459
rect 6516 24439 6518 24459
rect 6588 24439 6590 24459
rect 6612 24439 6614 24459
rect 6636 24439 6638 24459
rect 6684 24439 6686 24459
rect 6708 24439 6710 24459
rect 6769 24454 6772 24459
rect 6780 24454 6782 24459
rect 6779 24440 6782 24454
rect 6804 24439 6806 24459
rect 6900 24439 6902 24459
rect 7164 24439 7166 24459
rect 7236 24439 7238 24459
rect 7284 24439 7286 24459
rect 7380 24439 7382 24459
rect 7404 24439 7406 24459
rect 7476 24439 7478 24459
rect 7500 24439 7502 24459
rect 7537 24439 7571 24440
rect 7572 24439 7574 24459
rect 7644 24439 7646 24459
rect 7668 24439 7670 24459
rect 7908 24439 7910 24459
rect 8124 24439 8126 24459
rect 8220 24439 8222 24459
rect 8652 24439 8654 24459
rect 8700 24439 8702 24459
rect 8748 24439 8750 24459
rect 8796 24439 8798 24459
rect 8844 24439 8846 24459
rect 8868 24439 8870 24459
rect 9516 24439 9518 24459
rect 9660 24439 9662 24459
rect 9684 24439 9686 24459
rect 9780 24439 9782 24459
rect 9804 24439 9806 24459
rect 9828 24439 9830 24459
rect 10044 24439 10046 24459
rect 10140 24439 10142 24459
rect 10236 24439 10238 24459
rect 10332 24439 10334 24459
rect 10380 24439 10382 24459
rect 10428 24439 10430 24459
rect 10524 24439 10526 24459
rect 10548 24439 10550 24459
rect 10620 24439 10622 24459
rect 10644 24439 10646 24459
rect 10716 24439 10718 24459
rect 10884 24439 10886 24459
rect 10956 24439 10958 24459
rect 11052 24439 11054 24459
rect 11100 24439 11102 24459
rect 11172 24439 11174 24459
rect 11220 24439 11222 24459
rect 11340 24439 11342 24459
rect 11436 24439 11438 24459
rect 11676 24439 11678 24459
rect 11724 24439 11726 24459
rect 11772 24439 11774 24459
rect 11796 24439 11798 24459
rect 12060 24439 12062 24459
rect 12276 24439 12278 24459
rect 12324 24439 12326 24459
rect 12372 24439 12374 24459
rect 12420 24439 12422 24459
rect 12468 24439 12470 24459
rect 12564 24439 12566 24459
rect 12780 24439 12782 24459
rect 12828 24439 12830 24459
rect 12876 24439 12878 24459
rect 12972 24439 12974 24459
rect 13044 24439 13046 24459
rect 13068 24439 13070 24459
rect 13284 24439 13286 24459
rect 13332 24439 13334 24459
rect 13500 24439 13502 24459
rect 13572 24439 13574 24459
rect 13668 24439 13670 24459
rect 13716 24439 13718 24459
rect 13825 24454 13828 24459
rect 13956 24456 13958 24459
rect 13835 24440 13838 24454
rect 13836 24439 13838 24440
rect 13956 24439 13959 24456
rect 14004 24439 14006 24459
rect 14100 24439 14102 24459
rect 14940 24439 14942 24459
rect 15036 24439 15038 24459
rect 15276 24439 15278 24459
rect 15372 24439 15374 24459
rect 15420 24439 15422 24459
rect 15468 24439 15470 24459
rect 15564 24439 15566 24459
rect 15577 24439 15635 24440
rect 15660 24439 15662 24459
rect 15708 24439 15710 24459
rect 15732 24439 15734 24459
rect 15756 24439 15758 24459
rect 15804 24439 15806 24459
rect 15828 24439 15830 24459
rect 15852 24439 15854 24459
rect 15948 24439 15950 24459
rect 15972 24439 15974 24459
rect 16044 24439 16046 24459
rect 16068 24439 16070 24459
rect 16164 24439 16166 24459
rect 16260 24439 16262 24459
rect 16332 24439 16334 24459
rect 16380 24439 16382 24459
rect 16476 24439 16478 24459
rect 16548 24439 16550 24459
rect 16572 24439 16574 24459
rect 16668 24439 16670 24459
rect 16764 24439 16766 24459
rect 16812 24439 16814 24459
rect 16884 24439 16886 24459
rect 16908 24439 16910 24459
rect 17028 24439 17030 24459
rect 17124 24439 17126 24459
rect 17196 24439 17198 24459
rect 17220 24439 17222 24459
rect 17292 24439 17294 24459
rect 17316 24439 17318 24459
rect 17964 24439 17966 24459
rect 18060 24439 18062 24459
rect 18132 24439 18134 24459
rect 18228 24439 18230 24459
rect 18492 24439 18494 24459
rect 18540 24439 18542 24459
rect 18636 24439 18638 24459
rect 18732 24439 18734 24459
rect 18828 24439 18830 24459
rect 18924 24439 18926 24459
rect 18972 24439 18974 24459
rect 19020 24439 19022 24459
rect 19068 24439 19070 24459
rect 19140 24439 19142 24459
rect 19164 24439 19166 24459
rect 19236 24439 19238 24459
rect 19260 24439 19262 24459
rect 19788 24439 19790 24459
rect 19836 24439 19838 24459
rect 19860 24439 19862 24459
rect 19884 24439 19886 24459
rect 19956 24439 19958 24459
rect 19980 24439 19982 24459
rect 20004 24439 20006 24459
rect 20052 24439 20054 24459
rect 20076 24439 20078 24459
rect 20100 24439 20102 24459
rect 20172 24439 20174 24459
rect 20196 24439 20198 24459
rect 20292 24439 20294 24459
rect 20388 24439 20390 24459
rect 20412 24439 20414 24459
rect 20508 24439 20510 24459
rect 20532 24439 20534 24459
rect 20604 24439 20606 24459
rect 20628 24439 20630 24459
rect 20892 24439 20894 24459
rect 20964 24439 20966 24459
rect 20988 24439 20990 24459
rect 21108 24439 21110 24459
rect 21204 24439 21206 24459
rect 21300 24439 21302 24459
rect 21324 24439 21326 24459
rect 21444 24439 21446 24459
rect 21468 24439 21470 24459
rect 21564 24439 21566 24459
rect 21588 24439 21590 24459
rect 21684 24439 21686 24459
rect 21708 24439 21710 24459
rect 21841 24439 21875 24440
rect -8735 24435 -1915 24439
rect -8628 24432 -8626 24435
rect -8628 24416 -8625 24432
rect -8639 24415 -8605 24416
rect -8532 24415 -8530 24435
rect -8436 24415 -8434 24435
rect -8340 24415 -8338 24435
rect -8124 24415 -8122 24435
rect -7764 24415 -7762 24435
rect -7356 24415 -7354 24435
rect -7308 24415 -7306 24435
rect -7140 24415 -7138 24435
rect -6852 24432 -6850 24435
rect -6852 24415 -6849 24432
rect -6828 24415 -6825 24432
rect -6732 24415 -6730 24435
rect -6444 24415 -6442 24435
rect -6348 24415 -6346 24435
rect -6252 24415 -6250 24435
rect -5892 24415 -5890 24435
rect -5436 24432 -5434 24435
rect -5436 24415 -5433 24432
rect -5340 24415 -5338 24435
rect -4716 24415 -4714 24435
rect -4500 24415 -4498 24435
rect -4284 24415 -4282 24435
rect -3876 24415 -3874 24435
rect -3540 24415 -3538 24435
rect -3468 24415 -3466 24435
rect -3324 24415 -3322 24435
rect -3108 24415 -3106 24435
rect -3012 24415 -3010 24435
rect -2964 24415 -2962 24435
rect -2916 24415 -2914 24435
rect -2868 24415 -2866 24435
rect -2831 24430 -2828 24435
rect -2820 24430 -2818 24435
rect -2821 24416 -2818 24430
rect -2772 24415 -2770 24435
rect -2687 24430 -2684 24435
rect -2676 24430 -2674 24435
rect -2677 24416 -2674 24430
rect -2364 24415 -2362 24435
rect -1929 24432 -1915 24435
rect -1908 24435 6845 24439
rect -1908 24432 -1891 24435
rect -1908 24415 -1906 24432
rect -1452 24415 -1450 24435
rect -1356 24415 -1354 24435
rect -1260 24415 -1258 24435
rect -1236 24415 -1234 24435
rect -1140 24415 -1138 24435
rect -876 24415 -874 24435
rect -780 24415 -778 24435
rect -564 24415 -562 24435
rect -468 24415 -466 24435
rect -12 24415 -10 24435
rect 84 24415 86 24435
rect 252 24415 254 24435
rect 348 24415 350 24435
rect 468 24415 470 24435
rect 492 24415 494 24435
rect 564 24415 566 24435
rect 588 24415 590 24435
rect 636 24415 638 24435
rect 660 24415 662 24435
rect 732 24415 734 24435
rect 948 24415 950 24435
rect 1044 24415 1046 24435
rect 1092 24415 1094 24435
rect 1140 24415 1142 24435
rect 1308 24415 1310 24435
rect 1356 24415 1358 24435
rect 1428 24415 1430 24435
rect 1572 24415 1574 24435
rect 1860 24415 1862 24435
rect 1956 24415 1958 24435
rect 2052 24415 2054 24435
rect 2148 24415 2150 24435
rect 2244 24415 2246 24435
rect 2460 24415 2462 24435
rect 2772 24415 2774 24435
rect 2868 24415 2870 24435
rect 2940 24415 2942 24435
rect 2988 24415 2990 24435
rect 3324 24415 3326 24435
rect 3540 24415 3542 24435
rect 3660 24415 3662 24435
rect 3780 24415 3782 24435
rect 4092 24415 4094 24435
rect 4188 24415 4190 24435
rect 4308 24415 4310 24435
rect 4404 24415 4406 24435
rect 4500 24415 4502 24435
rect 4596 24415 4598 24435
rect 4692 24415 4694 24435
rect 4932 24415 4934 24435
rect 4980 24415 4982 24435
rect 5028 24415 5030 24435
rect 5124 24415 5126 24435
rect 5220 24415 5222 24435
rect 5388 24415 5390 24435
rect 5508 24415 5510 24435
rect 5556 24415 5558 24435
rect 5652 24415 5654 24435
rect 5748 24415 5750 24435
rect 5796 24415 5798 24435
rect 5844 24415 5846 24435
rect 5892 24415 5894 24435
rect 6276 24415 6278 24435
rect 6289 24415 6347 24416
rect 6372 24415 6374 24435
rect 6420 24415 6422 24435
rect 6492 24415 6494 24435
rect 6516 24415 6518 24435
rect 6588 24415 6590 24435
rect 6612 24415 6614 24435
rect 6636 24415 6638 24435
rect 6684 24415 6686 24435
rect 6708 24415 6710 24435
rect 6804 24415 6806 24435
rect 6831 24432 6845 24435
rect 6855 24435 13925 24439
rect 6855 24432 6869 24435
rect 6900 24415 6902 24435
rect 7164 24415 7166 24435
rect 7236 24415 7238 24435
rect 7284 24415 7286 24435
rect 7380 24415 7382 24435
rect 7404 24415 7406 24435
rect 7476 24415 7478 24435
rect 7500 24415 7502 24435
rect 7572 24415 7574 24435
rect 7644 24432 7646 24435
rect 7644 24415 7647 24432
rect 7668 24415 7670 24435
rect 7908 24415 7910 24435
rect 8124 24415 8126 24435
rect 8220 24415 8222 24435
rect 8652 24415 8654 24435
rect 8700 24415 8702 24435
rect 8748 24415 8750 24435
rect 8796 24415 8798 24435
rect 8844 24415 8846 24435
rect 8868 24415 8870 24435
rect 9516 24415 9518 24435
rect 9660 24415 9662 24435
rect 9684 24415 9686 24435
rect 9780 24415 9782 24435
rect 9804 24415 9806 24435
rect 9828 24415 9830 24435
rect 10044 24415 10046 24435
rect 10140 24415 10142 24435
rect 10236 24415 10238 24435
rect 10332 24415 10334 24435
rect 10380 24415 10382 24435
rect 10428 24415 10430 24435
rect 10524 24415 10526 24435
rect 10548 24415 10550 24435
rect 10620 24415 10622 24435
rect 10644 24415 10646 24435
rect 10716 24415 10718 24435
rect 10753 24415 10811 24416
rect 10884 24415 10886 24435
rect 10956 24415 10958 24435
rect 11052 24415 11054 24435
rect 11100 24415 11102 24435
rect 11172 24415 11174 24435
rect 11220 24415 11222 24435
rect 11340 24415 11342 24435
rect 11436 24415 11438 24435
rect 11676 24415 11678 24435
rect 11724 24415 11726 24435
rect 11772 24415 11774 24435
rect 11796 24415 11798 24435
rect 12060 24415 12062 24435
rect 12276 24415 12278 24435
rect 12324 24415 12326 24435
rect 12372 24415 12374 24435
rect 12420 24415 12422 24435
rect 12468 24415 12470 24435
rect 12564 24415 12566 24435
rect 12780 24415 12782 24435
rect 12828 24415 12830 24435
rect 12876 24415 12878 24435
rect 12972 24415 12974 24435
rect 13044 24415 13046 24435
rect 13068 24415 13070 24435
rect 13153 24415 13211 24416
rect 13284 24415 13286 24435
rect 13332 24415 13334 24435
rect 13500 24415 13502 24435
rect 13572 24415 13574 24435
rect 13668 24415 13670 24435
rect 13716 24415 13718 24435
rect 13836 24415 13838 24435
rect 13911 24432 13925 24435
rect 13935 24435 21875 24439
rect 13935 24432 13949 24435
rect 13956 24432 13959 24435
rect 14004 24415 14006 24435
rect 14100 24415 14102 24435
rect 14940 24415 14942 24435
rect 15036 24415 15038 24435
rect 15276 24415 15278 24435
rect 15372 24415 15374 24435
rect 15420 24415 15422 24435
rect 15468 24415 15470 24435
rect 15564 24415 15566 24435
rect 15660 24415 15662 24435
rect 15708 24432 15710 24435
rect 15708 24415 15711 24432
rect 15732 24415 15734 24435
rect 15756 24415 15758 24435
rect 15804 24415 15806 24435
rect 15828 24415 15830 24435
rect 15852 24415 15854 24435
rect 15948 24415 15950 24435
rect 15972 24415 15974 24435
rect 16044 24415 16046 24435
rect 16068 24415 16070 24435
rect 16164 24415 16166 24435
rect 16260 24415 16262 24435
rect 16332 24415 16334 24435
rect 16380 24415 16382 24435
rect 16476 24415 16478 24435
rect 16548 24415 16550 24435
rect 16572 24415 16574 24435
rect 16668 24415 16670 24435
rect 16764 24415 16766 24435
rect 16812 24415 16814 24435
rect 16884 24415 16886 24435
rect 16908 24415 16910 24435
rect 17028 24415 17030 24435
rect 17124 24415 17126 24435
rect 17196 24415 17198 24435
rect 17220 24415 17222 24435
rect 17292 24415 17294 24435
rect 17316 24415 17318 24435
rect 17964 24415 17966 24435
rect 18060 24415 18062 24435
rect 18132 24415 18134 24435
rect 18228 24415 18230 24435
rect 18492 24415 18494 24435
rect 18540 24415 18542 24435
rect 18636 24415 18638 24435
rect 18732 24415 18734 24435
rect 18828 24415 18830 24435
rect 18924 24415 18926 24435
rect 18972 24415 18974 24435
rect 19020 24415 19022 24435
rect 19068 24415 19070 24435
rect 19140 24415 19142 24435
rect 19164 24415 19166 24435
rect 19236 24415 19238 24435
rect 19260 24415 19262 24435
rect 19788 24415 19790 24435
rect 19836 24415 19838 24435
rect 19860 24415 19862 24435
rect 19884 24415 19886 24435
rect 19956 24415 19958 24435
rect 19980 24415 19982 24435
rect 20004 24415 20006 24435
rect 20052 24415 20054 24435
rect 20076 24415 20078 24435
rect 20100 24415 20102 24435
rect 20172 24415 20174 24435
rect 20196 24415 20198 24435
rect 20292 24415 20294 24435
rect 20388 24415 20390 24435
rect 20412 24415 20414 24435
rect 20508 24415 20510 24435
rect 20532 24415 20534 24435
rect 20604 24415 20606 24435
rect 20628 24415 20630 24435
rect 20892 24415 20894 24435
rect 20964 24415 20966 24435
rect 20988 24415 20990 24435
rect 21108 24415 21110 24435
rect 21204 24415 21206 24435
rect 21300 24415 21302 24435
rect 21324 24415 21326 24435
rect 21444 24415 21446 24435
rect 21468 24415 21470 24435
rect 21564 24415 21566 24435
rect 21588 24415 21590 24435
rect 21684 24415 21686 24435
rect 21708 24415 21710 24435
rect 21721 24415 21755 24416
rect -8639 24411 -6835 24415
rect -8639 24408 -8635 24411
rect -8628 24408 -8625 24411
rect -8532 24408 -8530 24411
rect -8532 24392 -8529 24408
rect -8436 24392 -8434 24411
rect -8543 24391 -8509 24392
rect -8471 24391 -8413 24392
rect -8340 24391 -8338 24411
rect -8124 24391 -8122 24411
rect -7764 24391 -7762 24411
rect -7356 24391 -7354 24411
rect -7308 24391 -7306 24411
rect -7140 24391 -7138 24411
rect -6873 24408 -6859 24411
rect -6852 24408 -6835 24411
rect -6828 24411 -5467 24415
rect -6828 24408 -6811 24411
rect -6828 24391 -6826 24408
rect -6732 24391 -6730 24411
rect -6444 24391 -6442 24411
rect -6348 24391 -6346 24411
rect -6252 24391 -6250 24411
rect -5892 24391 -5890 24411
rect -5481 24408 -5467 24411
rect -5457 24411 15677 24415
rect -5457 24408 -5443 24411
rect -5436 24408 -5433 24411
rect -5340 24391 -5338 24411
rect -4716 24391 -4714 24411
rect -4500 24391 -4498 24411
rect -4284 24391 -4282 24411
rect -3876 24391 -3874 24411
rect -3540 24391 -3538 24411
rect -3468 24391 -3466 24411
rect -3324 24391 -3322 24411
rect -3108 24391 -3106 24411
rect -3012 24391 -3010 24411
rect -2964 24391 -2962 24411
rect -2916 24391 -2914 24411
rect -2868 24391 -2866 24411
rect -2772 24391 -2770 24411
rect -2745 24408 -2731 24411
rect -2601 24408 -2587 24411
rect -2364 24391 -2362 24411
rect -1908 24391 -1906 24411
rect -1452 24391 -1450 24411
rect -1356 24391 -1354 24411
rect -1260 24391 -1258 24411
rect -1236 24391 -1234 24411
rect -1140 24391 -1138 24411
rect -876 24391 -874 24411
rect -780 24391 -778 24411
rect -564 24391 -562 24411
rect -468 24391 -466 24411
rect -12 24391 -10 24411
rect 84 24391 86 24411
rect 207 24408 221 24411
rect 252 24391 254 24411
rect 348 24391 350 24411
rect 468 24391 470 24411
rect 492 24391 494 24411
rect 564 24391 566 24411
rect 588 24391 590 24411
rect 636 24391 638 24411
rect 660 24391 662 24411
rect 732 24391 734 24411
rect 948 24391 950 24411
rect 1044 24391 1046 24411
rect 1092 24391 1094 24411
rect 1140 24391 1142 24411
rect 1308 24391 1310 24411
rect 1356 24391 1358 24411
rect 1428 24391 1430 24411
rect 1572 24391 1574 24411
rect 1860 24391 1862 24411
rect 1956 24391 1958 24411
rect 2052 24391 2054 24411
rect 2148 24391 2150 24411
rect 2244 24391 2246 24411
rect 2460 24391 2462 24411
rect 2772 24391 2774 24411
rect 2868 24391 2870 24411
rect 2940 24391 2942 24411
rect 2988 24391 2990 24411
rect 3324 24391 3326 24411
rect 3540 24391 3542 24411
rect 3660 24391 3662 24411
rect 3780 24391 3782 24411
rect 4092 24391 4094 24411
rect 4188 24391 4190 24411
rect 4308 24391 4310 24411
rect 4404 24391 4406 24411
rect 4500 24391 4502 24411
rect 4596 24391 4598 24411
rect 4692 24391 4694 24411
rect 4932 24391 4934 24411
rect 4980 24391 4982 24411
rect 5028 24391 5030 24411
rect 5124 24391 5126 24411
rect 5220 24391 5222 24411
rect 5388 24392 5390 24411
rect 5353 24391 5411 24392
rect 5508 24391 5510 24411
rect 5556 24391 5558 24411
rect 5652 24391 5654 24411
rect 5748 24391 5750 24411
rect 5796 24391 5798 24411
rect 5844 24391 5846 24411
rect 5892 24391 5894 24411
rect 6276 24391 6278 24411
rect 6289 24406 6292 24411
rect 6299 24392 6302 24406
rect 6300 24391 6302 24392
rect 6372 24391 6374 24411
rect 6420 24408 6422 24411
rect 6396 24391 6399 24408
rect 6420 24391 6423 24408
rect 6492 24391 6494 24411
rect 6516 24391 6518 24411
rect 6588 24391 6590 24411
rect 6612 24391 6614 24411
rect 6636 24391 6638 24411
rect 6684 24391 6686 24411
rect 6708 24391 6710 24411
rect 6804 24391 6806 24411
rect 6900 24391 6902 24411
rect 7164 24391 7166 24411
rect 7236 24391 7238 24411
rect 7284 24391 7286 24411
rect 7380 24391 7382 24411
rect 7404 24391 7406 24411
rect 7476 24391 7478 24411
rect 7500 24391 7502 24411
rect 7572 24391 7574 24411
rect 7623 24408 7637 24411
rect 7644 24408 7647 24411
rect 7668 24391 7670 24411
rect 7908 24391 7910 24411
rect 8124 24391 8126 24411
rect 8220 24391 8222 24411
rect 8652 24391 8654 24411
rect 8700 24391 8702 24411
rect 8748 24391 8750 24411
rect 8796 24391 8798 24411
rect 8844 24391 8846 24411
rect 8868 24391 8870 24411
rect 9516 24391 9518 24411
rect 9660 24391 9662 24411
rect 9684 24391 9686 24411
rect 9780 24391 9782 24411
rect 9804 24391 9806 24411
rect 9828 24391 9830 24411
rect 10044 24391 10046 24411
rect 10140 24391 10142 24411
rect 10236 24391 10238 24411
rect 10332 24391 10334 24411
rect 10380 24391 10382 24411
rect 10428 24391 10430 24411
rect 10524 24391 10526 24411
rect 10548 24391 10550 24411
rect 10620 24391 10622 24411
rect 10644 24391 10646 24411
rect 10716 24391 10718 24411
rect 10884 24408 10886 24411
rect 10860 24391 10863 24408
rect 10884 24391 10887 24408
rect 10956 24391 10958 24411
rect 11052 24391 11054 24411
rect 11100 24391 11102 24411
rect 11172 24391 11174 24411
rect 11220 24391 11222 24411
rect 11340 24391 11342 24411
rect 11436 24391 11438 24411
rect 11676 24391 11678 24411
rect 11724 24391 11726 24411
rect 11772 24391 11774 24411
rect 11796 24391 11798 24411
rect 12060 24391 12062 24411
rect 12276 24391 12278 24411
rect 12324 24391 12326 24411
rect 12372 24391 12374 24411
rect 12420 24391 12422 24411
rect 12468 24391 12470 24411
rect 12564 24391 12566 24411
rect 12780 24391 12782 24411
rect 12828 24391 12830 24411
rect 12876 24391 12878 24411
rect 12972 24391 12974 24411
rect 13044 24391 13046 24411
rect 13068 24391 13070 24411
rect 13153 24406 13156 24411
rect 13284 24408 13286 24411
rect 13163 24392 13166 24406
rect 13164 24391 13166 24392
rect 13284 24391 13287 24408
rect 13332 24391 13334 24411
rect 13500 24391 13502 24411
rect 13572 24391 13574 24411
rect 13668 24391 13670 24411
rect 13716 24391 13718 24411
rect 13836 24391 13838 24411
rect 14004 24391 14006 24411
rect 14100 24391 14102 24411
rect 14940 24391 14942 24411
rect 15036 24391 15038 24411
rect 15276 24391 15278 24411
rect 15372 24391 15374 24411
rect 15420 24391 15422 24411
rect 15468 24391 15470 24411
rect 15564 24391 15566 24411
rect 15660 24391 15662 24411
rect 15663 24408 15677 24411
rect 15687 24411 21755 24415
rect 15687 24408 15701 24411
rect 15708 24408 15711 24411
rect 15732 24391 15734 24411
rect 15756 24391 15758 24411
rect 15804 24391 15806 24411
rect 15828 24391 15830 24411
rect 15852 24391 15854 24411
rect 15948 24391 15950 24411
rect 15972 24391 15974 24411
rect 16044 24391 16046 24411
rect 16068 24391 16070 24411
rect 16164 24391 16166 24411
rect 16177 24391 16235 24392
rect 16260 24391 16262 24411
rect 16332 24391 16334 24411
rect 16380 24391 16382 24411
rect 16476 24391 16478 24411
rect 16548 24391 16550 24411
rect 16572 24391 16574 24411
rect 16668 24391 16670 24411
rect 16764 24391 16766 24411
rect 16812 24391 16814 24411
rect 16884 24391 16886 24411
rect 16908 24391 16910 24411
rect 17028 24391 17030 24411
rect 17124 24391 17126 24411
rect 17196 24391 17198 24411
rect 17220 24391 17222 24411
rect 17292 24391 17294 24411
rect 17316 24391 17318 24411
rect 17964 24391 17966 24411
rect 18060 24391 18062 24411
rect 18132 24391 18134 24411
rect 18228 24391 18230 24411
rect 18492 24391 18494 24411
rect 18540 24391 18542 24411
rect 18636 24391 18638 24411
rect 18732 24391 18734 24411
rect 18828 24391 18830 24411
rect 18924 24391 18926 24411
rect 18972 24391 18974 24411
rect 19020 24391 19022 24411
rect 19068 24391 19070 24411
rect 19140 24391 19142 24411
rect 19164 24391 19166 24411
rect 19236 24391 19238 24411
rect 19260 24391 19262 24411
rect 19788 24391 19790 24411
rect 19836 24391 19838 24411
rect 19860 24391 19862 24411
rect 19884 24391 19886 24411
rect 19956 24391 19958 24411
rect 19980 24391 19982 24411
rect 20004 24391 20006 24411
rect 20052 24391 20054 24411
rect 20076 24391 20078 24411
rect 20100 24391 20102 24411
rect 20172 24391 20174 24411
rect 20196 24391 20198 24411
rect 20292 24391 20294 24411
rect 20388 24391 20390 24411
rect 20412 24391 20414 24411
rect 20508 24391 20510 24411
rect 20532 24391 20534 24411
rect 20604 24391 20606 24411
rect 20628 24391 20630 24411
rect 20892 24391 20894 24411
rect 20964 24391 20966 24411
rect 20988 24391 20990 24411
rect 21108 24391 21110 24411
rect 21204 24391 21206 24411
rect 21300 24391 21302 24411
rect 21324 24391 21326 24411
rect 21444 24391 21446 24411
rect 21468 24391 21470 24411
rect 21564 24391 21566 24411
rect 21588 24391 21590 24411
rect 21684 24391 21686 24411
rect 21708 24392 21710 24411
rect 21697 24391 21731 24392
rect -8543 24387 6389 24391
rect -8543 24384 -8539 24387
rect -8532 24384 -8529 24387
rect -8447 24382 -8444 24387
rect -8436 24384 -8434 24387
rect -8340 24384 -8338 24387
rect -8436 24382 -8433 24384
rect -8447 24374 -8443 24382
rect -8457 24368 -8447 24374
rect -8437 24368 -8433 24382
rect -8340 24368 -8337 24384
rect -8351 24367 -8317 24368
rect -8279 24367 -8245 24368
rect -8351 24363 -8245 24367
rect -8231 24367 -8197 24368
rect -8124 24367 -8122 24387
rect -7764 24367 -7762 24387
rect -7356 24367 -7354 24387
rect -7308 24367 -7306 24387
rect -7140 24367 -7138 24387
rect -6828 24367 -6826 24387
rect -6732 24367 -6730 24387
rect -6444 24367 -6442 24387
rect -6348 24367 -6346 24387
rect -6252 24367 -6250 24387
rect -5892 24367 -5890 24387
rect -5340 24367 -5338 24387
rect -4716 24367 -4714 24387
rect -4500 24367 -4498 24387
rect -4284 24367 -4282 24387
rect -3876 24367 -3874 24387
rect -3540 24367 -3538 24387
rect -3468 24367 -3466 24387
rect -3324 24367 -3322 24387
rect -3108 24367 -3106 24387
rect -3012 24367 -3010 24387
rect -2964 24367 -2962 24387
rect -2916 24367 -2914 24387
rect -2868 24367 -2866 24387
rect -2772 24367 -2770 24387
rect -2364 24367 -2362 24387
rect -1908 24367 -1906 24387
rect -1452 24367 -1450 24387
rect -1356 24367 -1354 24387
rect -1260 24367 -1258 24387
rect -1236 24367 -1234 24387
rect -1140 24367 -1138 24387
rect -876 24367 -874 24387
rect -780 24367 -778 24387
rect -564 24367 -562 24387
rect -468 24367 -466 24387
rect -12 24367 -10 24387
rect 84 24367 86 24387
rect 252 24367 254 24387
rect 348 24367 350 24387
rect 468 24367 470 24387
rect 492 24367 494 24387
rect 564 24367 566 24387
rect 588 24367 590 24387
rect 636 24367 638 24387
rect 660 24367 662 24387
rect 732 24367 734 24387
rect 948 24367 950 24387
rect 1044 24367 1046 24387
rect 1092 24367 1094 24387
rect 1140 24367 1142 24387
rect 1308 24367 1310 24387
rect 1356 24367 1358 24387
rect 1428 24367 1430 24387
rect 1572 24367 1574 24387
rect 1860 24367 1862 24387
rect 1956 24367 1958 24387
rect 2052 24367 2054 24387
rect 2148 24367 2150 24387
rect 2244 24367 2246 24387
rect 2460 24367 2462 24387
rect 2772 24367 2774 24387
rect 2868 24367 2870 24387
rect 2940 24367 2942 24387
rect 2988 24367 2990 24387
rect 3324 24367 3326 24387
rect 3540 24367 3542 24387
rect 3660 24367 3662 24387
rect 3780 24367 3782 24387
rect 4092 24367 4094 24387
rect 4188 24367 4190 24387
rect 4308 24367 4310 24387
rect 4404 24367 4406 24387
rect 4500 24367 4502 24387
rect 4596 24367 4598 24387
rect 4692 24367 4694 24387
rect 4932 24367 4934 24387
rect 4980 24367 4982 24387
rect 5028 24367 5030 24387
rect 5124 24367 5126 24387
rect 5220 24367 5222 24387
rect 5377 24382 5380 24387
rect 5388 24382 5390 24387
rect 5387 24368 5390 24382
rect 5460 24367 5463 24384
rect 5508 24367 5510 24387
rect 5556 24367 5558 24387
rect 5652 24367 5654 24387
rect 5748 24367 5750 24387
rect 5796 24367 5798 24387
rect 5844 24367 5846 24387
rect 5892 24367 5894 24387
rect 6276 24367 6278 24387
rect 6300 24367 6302 24387
rect 6372 24367 6374 24387
rect 6375 24384 6389 24387
rect 6396 24387 10853 24391
rect 6396 24384 6413 24387
rect 6420 24384 6423 24387
rect 6396 24367 6398 24384
rect 6492 24367 6494 24387
rect 6516 24367 6518 24387
rect 6588 24367 6590 24387
rect 6612 24367 6614 24387
rect 6636 24367 6638 24387
rect 6684 24367 6686 24387
rect 6708 24367 6710 24387
rect 6804 24367 6806 24387
rect 6900 24367 6902 24387
rect 7164 24367 7166 24387
rect 7236 24367 7238 24387
rect 7284 24367 7286 24387
rect 7380 24367 7382 24387
rect 7404 24367 7406 24387
rect 7476 24367 7478 24387
rect 7500 24367 7502 24387
rect 7572 24367 7574 24387
rect 7668 24367 7670 24387
rect 7908 24367 7910 24387
rect 8124 24367 8126 24387
rect 8220 24367 8222 24387
rect 8652 24367 8654 24387
rect 8700 24367 8702 24387
rect 8748 24367 8750 24387
rect 8796 24367 8798 24387
rect 8844 24367 8846 24387
rect 8868 24367 8870 24387
rect 9516 24367 9518 24387
rect 9660 24367 9662 24387
rect 9684 24367 9686 24387
rect 9780 24367 9782 24387
rect 9804 24367 9806 24387
rect 9828 24367 9830 24387
rect 10044 24367 10046 24387
rect 10140 24367 10142 24387
rect 10236 24367 10238 24387
rect 10332 24367 10334 24387
rect 10380 24367 10382 24387
rect 10428 24367 10430 24387
rect 10524 24367 10526 24387
rect 10548 24367 10550 24387
rect 10620 24367 10622 24387
rect 10644 24367 10646 24387
rect 10716 24367 10718 24387
rect 10839 24384 10853 24387
rect 10860 24387 13253 24391
rect 10860 24384 10877 24387
rect 10884 24384 10887 24387
rect 10860 24367 10862 24384
rect 10956 24367 10958 24387
rect 11052 24367 11054 24387
rect 11100 24367 11102 24387
rect 11172 24367 11174 24387
rect 11220 24367 11222 24387
rect 11340 24367 11342 24387
rect 11436 24367 11438 24387
rect 11676 24367 11678 24387
rect 11724 24367 11726 24387
rect 11772 24367 11774 24387
rect 11796 24367 11798 24387
rect 12060 24367 12062 24387
rect 12276 24367 12278 24387
rect 12324 24367 12326 24387
rect 12372 24367 12374 24387
rect 12420 24367 12422 24387
rect 12468 24367 12470 24387
rect 12564 24367 12566 24387
rect 12780 24367 12782 24387
rect 12828 24367 12830 24387
rect 12876 24367 12878 24387
rect 12972 24367 12974 24387
rect 13044 24367 13046 24387
rect 13068 24367 13070 24387
rect 13164 24367 13166 24387
rect 13239 24384 13253 24387
rect 13263 24387 21731 24391
rect 13263 24384 13277 24387
rect 13284 24384 13287 24387
rect 13332 24367 13334 24387
rect 13500 24367 13502 24387
rect 13572 24367 13574 24387
rect 13668 24367 13670 24387
rect 13716 24367 13718 24387
rect 13836 24367 13838 24387
rect 14004 24367 14006 24387
rect 14100 24367 14102 24387
rect 14940 24367 14942 24387
rect 15036 24367 15038 24387
rect 15276 24367 15278 24387
rect 15372 24367 15374 24387
rect 15420 24367 15422 24387
rect 15468 24367 15470 24387
rect 15564 24367 15566 24387
rect 15660 24367 15662 24387
rect 15732 24367 15734 24387
rect 15756 24367 15758 24387
rect 15804 24367 15806 24387
rect 15828 24367 15830 24387
rect 15852 24367 15854 24387
rect 15948 24367 15950 24387
rect 15972 24367 15974 24387
rect 16044 24367 16046 24387
rect 16068 24367 16070 24387
rect 16164 24367 16166 24387
rect 16260 24367 16262 24387
rect 16284 24367 16287 24384
rect 16332 24367 16334 24387
rect 16380 24367 16382 24387
rect 16476 24367 16478 24387
rect 16548 24367 16550 24387
rect 16572 24367 16574 24387
rect 16668 24367 16670 24387
rect 16764 24367 16766 24387
rect 16812 24367 16814 24387
rect 16884 24367 16886 24387
rect 16908 24367 16910 24387
rect 17028 24367 17030 24387
rect 17124 24367 17126 24387
rect 17196 24367 17198 24387
rect 17220 24367 17222 24387
rect 17292 24367 17294 24387
rect 17316 24367 17318 24387
rect 17964 24367 17966 24387
rect 18060 24367 18062 24387
rect 18132 24367 18134 24387
rect 18228 24367 18230 24387
rect 18492 24367 18494 24387
rect 18540 24367 18542 24387
rect 18636 24367 18638 24387
rect 18732 24367 18734 24387
rect 18828 24367 18830 24387
rect 18924 24367 18926 24387
rect 18972 24367 18974 24387
rect 19020 24367 19022 24387
rect 19068 24367 19070 24387
rect 19140 24367 19142 24387
rect 19164 24367 19166 24387
rect 19236 24367 19238 24387
rect 19260 24367 19262 24387
rect 19788 24367 19790 24387
rect 19836 24367 19838 24387
rect 19860 24367 19862 24387
rect 19884 24367 19886 24387
rect 19956 24367 19958 24387
rect 19980 24367 19982 24387
rect 20004 24367 20006 24387
rect 20052 24367 20054 24387
rect 20076 24367 20078 24387
rect 20100 24367 20102 24387
rect 20172 24367 20174 24387
rect 20196 24367 20198 24387
rect 20292 24367 20294 24387
rect 20388 24367 20390 24387
rect 20412 24367 20414 24387
rect 20508 24367 20510 24387
rect 20532 24367 20534 24387
rect 20604 24367 20606 24387
rect 20628 24367 20630 24387
rect 20892 24367 20894 24387
rect 20964 24367 20966 24387
rect 20988 24367 20990 24387
rect 21108 24367 21110 24387
rect 21204 24367 21206 24387
rect 21300 24367 21302 24387
rect 21324 24367 21326 24387
rect 21444 24367 21446 24387
rect 21468 24367 21470 24387
rect 21564 24367 21566 24387
rect 21588 24367 21590 24387
rect 21684 24368 21686 24387
rect 21697 24382 21700 24387
rect 21708 24382 21710 24387
rect 21707 24368 21710 24382
rect 21673 24367 21707 24368
rect -8231 24363 5453 24367
rect -8351 24360 -8347 24363
rect -8340 24360 -8337 24363
rect -8124 24360 -8122 24363
rect -8255 24350 -8251 24358
rect -8265 24344 -8255 24350
rect -8124 24344 -8121 24360
rect -8135 24343 -8101 24344
rect -7764 24343 -7762 24363
rect -7356 24343 -7354 24363
rect -7308 24343 -7306 24363
rect -7140 24343 -7138 24363
rect -6828 24343 -6826 24363
rect -6732 24343 -6730 24363
rect -6444 24343 -6442 24363
rect -6348 24343 -6346 24363
rect -6252 24343 -6250 24363
rect -5892 24343 -5890 24363
rect -5340 24343 -5338 24363
rect -4991 24343 -4957 24344
rect -4716 24343 -4714 24363
rect -4500 24343 -4498 24363
rect -4284 24343 -4282 24363
rect -3876 24343 -3874 24363
rect -3540 24343 -3538 24363
rect -3468 24343 -3466 24363
rect -3324 24343 -3322 24363
rect -3108 24343 -3106 24363
rect -3012 24343 -3010 24363
rect -2964 24343 -2962 24363
rect -2916 24343 -2914 24363
rect -2868 24343 -2866 24363
rect -2772 24343 -2770 24363
rect -2364 24343 -2362 24363
rect -1908 24343 -1906 24363
rect -1452 24343 -1450 24363
rect -1356 24343 -1354 24363
rect -1260 24343 -1258 24363
rect -1236 24343 -1234 24363
rect -1140 24343 -1138 24363
rect -876 24343 -874 24363
rect -780 24343 -778 24363
rect -564 24343 -562 24363
rect -468 24343 -466 24363
rect -12 24343 -10 24363
rect 84 24343 86 24363
rect 252 24343 254 24363
rect 348 24343 350 24363
rect 468 24343 470 24363
rect 492 24343 494 24363
rect 564 24343 566 24363
rect 588 24343 590 24363
rect 636 24343 638 24363
rect 660 24343 662 24363
rect 732 24343 734 24363
rect 948 24343 950 24363
rect 1044 24343 1046 24363
rect 1092 24343 1094 24363
rect 1140 24343 1142 24363
rect 1308 24343 1310 24363
rect 1356 24343 1358 24363
rect 1428 24343 1430 24363
rect 1572 24343 1574 24363
rect 1860 24343 1862 24363
rect 1956 24343 1958 24363
rect 2052 24343 2054 24363
rect 2148 24343 2150 24363
rect 2244 24343 2246 24363
rect 2460 24343 2462 24363
rect 2772 24343 2774 24363
rect 2868 24343 2870 24363
rect 2940 24343 2942 24363
rect 2988 24343 2990 24363
rect 3324 24343 3326 24363
rect 3540 24343 3542 24363
rect 3660 24343 3662 24363
rect 3780 24343 3782 24363
rect 4092 24343 4094 24363
rect 4188 24343 4190 24363
rect 4308 24343 4310 24363
rect 4404 24343 4406 24363
rect 4500 24343 4502 24363
rect 4596 24343 4598 24363
rect 4692 24343 4694 24363
rect 4932 24343 4934 24363
rect 4980 24343 4982 24363
rect 5028 24343 5030 24363
rect 5124 24343 5126 24363
rect 5220 24343 5222 24363
rect 5439 24360 5453 24363
rect 5460 24363 16277 24367
rect 5460 24360 5477 24363
rect 5460 24343 5462 24360
rect 5508 24343 5510 24363
rect 5556 24343 5558 24363
rect 5652 24343 5654 24363
rect 5748 24343 5750 24363
rect 5796 24343 5798 24363
rect 5844 24343 5846 24363
rect 5892 24343 5894 24363
rect 6276 24343 6278 24363
rect 6300 24343 6302 24363
rect 6372 24343 6374 24363
rect 6396 24343 6398 24363
rect 6492 24343 6494 24363
rect 6516 24343 6518 24363
rect 6588 24343 6590 24363
rect 6612 24343 6614 24363
rect 6636 24343 6638 24363
rect 6684 24343 6686 24363
rect 6708 24343 6710 24363
rect 6804 24343 6806 24363
rect 6900 24343 6902 24363
rect 7164 24343 7166 24363
rect 7236 24343 7238 24363
rect 7284 24343 7286 24363
rect 7380 24343 7382 24363
rect 7404 24343 7406 24363
rect 7476 24343 7478 24363
rect 7500 24343 7502 24363
rect 7572 24343 7574 24363
rect 7585 24343 7643 24344
rect 7668 24343 7670 24363
rect 7908 24343 7910 24363
rect 8124 24343 8126 24363
rect 8220 24343 8222 24363
rect 8652 24343 8654 24363
rect 8700 24343 8702 24363
rect 8748 24343 8750 24363
rect 8796 24343 8798 24363
rect 8844 24343 8846 24363
rect 8868 24343 8870 24363
rect 9516 24343 9518 24363
rect 9660 24343 9662 24363
rect 9684 24343 9686 24363
rect 9780 24343 9782 24363
rect 9804 24343 9806 24363
rect 9828 24343 9830 24363
rect 10044 24343 10046 24363
rect 10140 24343 10142 24363
rect 10236 24343 10238 24363
rect 10332 24343 10334 24363
rect 10380 24343 10382 24363
rect 10428 24343 10430 24363
rect 10524 24343 10526 24363
rect 10548 24343 10550 24363
rect 10620 24343 10622 24363
rect 10644 24343 10646 24363
rect 10716 24343 10718 24363
rect 10860 24343 10862 24363
rect 10956 24343 10958 24363
rect 11052 24343 11054 24363
rect 11100 24343 11102 24363
rect 11172 24343 11174 24363
rect 11220 24343 11222 24363
rect 11340 24343 11342 24363
rect 11436 24343 11438 24363
rect 11676 24343 11678 24363
rect 11724 24343 11726 24363
rect 11772 24343 11774 24363
rect 11796 24343 11798 24363
rect 12060 24343 12062 24363
rect 12276 24343 12278 24363
rect 12324 24343 12326 24363
rect 12372 24343 12374 24363
rect 12420 24343 12422 24363
rect 12468 24343 12470 24363
rect 12564 24343 12566 24363
rect 12780 24343 12782 24363
rect 12828 24343 12830 24363
rect 12876 24343 12878 24363
rect 12972 24343 12974 24363
rect 13044 24343 13046 24363
rect 13068 24343 13070 24363
rect 13164 24343 13166 24363
rect 13332 24343 13334 24363
rect 13500 24343 13502 24363
rect 13572 24343 13574 24363
rect 13668 24343 13670 24363
rect 13716 24343 13718 24363
rect 13836 24343 13838 24363
rect 14004 24343 14006 24363
rect 14100 24343 14102 24363
rect 14940 24343 14942 24363
rect 15036 24343 15038 24363
rect 15276 24343 15278 24363
rect 15372 24343 15374 24363
rect 15420 24343 15422 24363
rect 15468 24343 15470 24363
rect 15564 24343 15566 24363
rect 15660 24343 15662 24363
rect 15732 24343 15734 24363
rect 15756 24343 15758 24363
rect 15804 24343 15806 24363
rect 15828 24343 15830 24363
rect 15852 24343 15854 24363
rect 15948 24343 15950 24363
rect 15972 24343 15974 24363
rect 16044 24343 16046 24363
rect 16068 24343 16070 24363
rect 16164 24343 16166 24363
rect 16260 24343 16262 24363
rect 16263 24360 16277 24363
rect 16284 24363 21707 24367
rect 16284 24360 16301 24363
rect 16284 24343 16286 24360
rect 16332 24343 16334 24363
rect 16380 24343 16382 24363
rect 16476 24343 16478 24363
rect 16548 24343 16550 24363
rect 16572 24343 16574 24363
rect 16668 24343 16670 24363
rect 16764 24343 16766 24363
rect 16812 24343 16814 24363
rect 16884 24343 16886 24363
rect 16908 24343 16910 24363
rect 17028 24343 17030 24363
rect 17124 24343 17126 24363
rect 17196 24343 17198 24363
rect 17220 24343 17222 24363
rect 17292 24343 17294 24363
rect 17316 24343 17318 24363
rect 17964 24343 17966 24363
rect 18060 24343 18062 24363
rect 18132 24343 18134 24363
rect 18228 24343 18230 24363
rect 18492 24343 18494 24363
rect 18540 24343 18542 24363
rect 18636 24343 18638 24363
rect 18732 24343 18734 24363
rect 18828 24343 18830 24363
rect 18924 24343 18926 24363
rect 18972 24343 18974 24363
rect 19020 24343 19022 24363
rect 19068 24343 19070 24363
rect 19140 24343 19142 24363
rect 19164 24343 19166 24363
rect 19236 24343 19238 24363
rect 19260 24343 19262 24363
rect 19788 24343 19790 24363
rect 19836 24343 19838 24363
rect 19860 24343 19862 24363
rect 19884 24343 19886 24363
rect 19956 24343 19958 24363
rect 19980 24343 19982 24363
rect 20004 24343 20006 24363
rect 20052 24343 20054 24363
rect 20076 24343 20078 24363
rect 20100 24343 20102 24363
rect 20172 24343 20174 24363
rect 20196 24343 20198 24363
rect 20292 24343 20294 24363
rect 20388 24343 20390 24363
rect 20412 24343 20414 24363
rect 20508 24343 20510 24363
rect 20532 24343 20534 24363
rect 20604 24343 20606 24363
rect 20628 24343 20630 24363
rect 20892 24343 20894 24363
rect 20964 24343 20966 24363
rect 20988 24343 20990 24363
rect 21108 24343 21110 24363
rect 21204 24343 21206 24363
rect 21300 24343 21302 24363
rect 21324 24343 21326 24363
rect 21444 24343 21446 24363
rect 21468 24343 21470 24363
rect 21564 24343 21566 24363
rect 21588 24343 21590 24363
rect 21673 24358 21676 24363
rect 21684 24358 21686 24363
rect 21683 24344 21686 24358
rect 21601 24343 21635 24344
rect -8135 24339 21635 24343
rect -8135 24336 -8131 24339
rect -8124 24336 -8121 24339
rect -8015 24319 -7981 24320
rect -7764 24319 -7762 24339
rect -7356 24319 -7354 24339
rect -7308 24319 -7306 24339
rect -7140 24319 -7138 24339
rect -6828 24319 -6826 24339
rect -6732 24319 -6730 24339
rect -6444 24319 -6442 24339
rect -6348 24319 -6346 24339
rect -6252 24319 -6250 24339
rect -5892 24319 -5890 24339
rect -5340 24319 -5338 24339
rect -4716 24319 -4714 24339
rect -4500 24319 -4498 24339
rect -4284 24319 -4282 24339
rect -4055 24319 -3997 24320
rect -3876 24319 -3874 24339
rect -3540 24319 -3538 24339
rect -3468 24319 -3466 24339
rect -3324 24319 -3322 24339
rect -3108 24319 -3106 24339
rect -3012 24319 -3010 24339
rect -2964 24319 -2962 24339
rect -2916 24319 -2914 24339
rect -2868 24319 -2866 24339
rect -2772 24319 -2770 24339
rect -2364 24319 -2362 24339
rect -1908 24319 -1906 24339
rect -1452 24319 -1450 24339
rect -1356 24319 -1354 24339
rect -1260 24319 -1258 24339
rect -1236 24319 -1234 24339
rect -1140 24319 -1138 24339
rect -876 24319 -874 24339
rect -780 24319 -778 24339
rect -564 24319 -562 24339
rect -468 24319 -466 24339
rect -12 24319 -10 24339
rect 84 24319 86 24339
rect 145 24319 179 24320
rect 252 24319 254 24339
rect 348 24319 350 24339
rect 468 24319 470 24339
rect 492 24319 494 24339
rect 564 24319 566 24339
rect 588 24319 590 24339
rect 636 24319 638 24339
rect 660 24319 662 24339
rect 732 24319 734 24339
rect 948 24319 950 24339
rect 1044 24319 1046 24339
rect 1092 24319 1094 24339
rect 1140 24319 1142 24339
rect 1308 24319 1310 24339
rect 1356 24319 1358 24339
rect 1428 24319 1430 24339
rect 1572 24319 1574 24339
rect 1860 24319 1862 24339
rect 1956 24319 1958 24339
rect 2052 24319 2054 24339
rect 2148 24319 2150 24339
rect 2244 24319 2246 24339
rect 2460 24319 2462 24339
rect 2772 24319 2774 24339
rect 2868 24319 2870 24339
rect 2940 24319 2942 24339
rect 2988 24319 2990 24339
rect 3324 24319 3326 24339
rect 3540 24319 3542 24339
rect 3660 24319 3662 24339
rect 3780 24319 3782 24339
rect 4092 24319 4094 24339
rect 4188 24319 4190 24339
rect 4308 24319 4310 24339
rect 4404 24319 4406 24339
rect 4500 24319 4502 24339
rect 4596 24319 4598 24339
rect 4692 24319 4694 24339
rect 4932 24319 4934 24339
rect 4980 24319 4982 24339
rect 5028 24319 5030 24339
rect 5124 24319 5126 24339
rect 5220 24319 5222 24339
rect 5460 24319 5462 24339
rect 5508 24319 5510 24339
rect 5556 24319 5558 24339
rect 5652 24319 5654 24339
rect 5748 24319 5750 24339
rect 5796 24319 5798 24339
rect 5844 24319 5846 24339
rect 5892 24319 5894 24339
rect 6276 24319 6278 24339
rect 6300 24319 6302 24339
rect 6372 24319 6374 24339
rect 6396 24319 6398 24339
rect 6492 24319 6494 24339
rect 6516 24319 6518 24339
rect 6588 24319 6590 24339
rect 6612 24319 6614 24339
rect 6636 24319 6638 24339
rect 6684 24319 6686 24339
rect 6708 24319 6710 24339
rect 6804 24319 6806 24339
rect 6900 24319 6902 24339
rect 7164 24319 7166 24339
rect 7236 24319 7238 24339
rect 7284 24319 7286 24339
rect 7380 24319 7382 24339
rect 7404 24319 7406 24339
rect 7476 24319 7478 24339
rect 7500 24319 7502 24339
rect 7572 24319 7574 24339
rect 7585 24334 7588 24339
rect 7595 24320 7598 24334
rect 7596 24319 7598 24320
rect 7668 24319 7670 24339
rect 7692 24319 7695 24336
rect 7908 24319 7910 24339
rect 8124 24319 8126 24339
rect 8220 24319 8222 24339
rect 8521 24319 8579 24320
rect 8652 24319 8654 24339
rect 8700 24319 8702 24339
rect 8748 24319 8750 24339
rect 8796 24319 8798 24339
rect 8844 24319 8846 24339
rect 8868 24319 8870 24339
rect 9516 24319 9518 24339
rect 9660 24319 9662 24339
rect 9684 24319 9686 24339
rect 9780 24319 9782 24339
rect 9804 24319 9806 24339
rect 9828 24319 9830 24339
rect 10044 24319 10046 24339
rect 10140 24319 10142 24339
rect 10236 24319 10238 24339
rect 10332 24319 10334 24339
rect 10380 24319 10382 24339
rect 10428 24319 10430 24339
rect 10524 24319 10526 24339
rect 10548 24319 10550 24339
rect 10620 24319 10622 24339
rect 10644 24319 10646 24339
rect 10716 24319 10718 24339
rect 10860 24319 10862 24339
rect 10956 24319 10958 24339
rect 11052 24319 11054 24339
rect 11100 24319 11102 24339
rect 11172 24319 11174 24339
rect 11220 24319 11222 24339
rect 11340 24319 11342 24339
rect 11436 24319 11438 24339
rect 11676 24319 11678 24339
rect 11724 24319 11726 24339
rect 11772 24319 11774 24339
rect 11796 24319 11798 24339
rect 12060 24319 12062 24339
rect 12276 24319 12278 24339
rect 12324 24319 12326 24339
rect 12372 24319 12374 24339
rect 12420 24319 12422 24339
rect 12468 24319 12470 24339
rect 12564 24319 12566 24339
rect 12780 24319 12782 24339
rect 12828 24319 12830 24339
rect 12876 24319 12878 24339
rect 12972 24319 12974 24339
rect 13044 24319 13046 24339
rect 13068 24319 13070 24339
rect 13164 24319 13166 24339
rect 13332 24319 13334 24339
rect 13500 24319 13502 24339
rect 13572 24319 13574 24339
rect 13668 24319 13670 24339
rect 13716 24319 13718 24339
rect 13836 24319 13838 24339
rect 14004 24319 14006 24339
rect 14100 24319 14102 24339
rect 14940 24319 14942 24339
rect 15036 24319 15038 24339
rect 15276 24319 15278 24339
rect 15372 24319 15374 24339
rect 15420 24319 15422 24339
rect 15468 24319 15470 24339
rect 15564 24319 15566 24339
rect 15660 24319 15662 24339
rect 15732 24319 15734 24339
rect 15756 24319 15758 24339
rect 15804 24319 15806 24339
rect 15828 24319 15830 24339
rect 15852 24319 15854 24339
rect 15948 24319 15950 24339
rect 15972 24319 15974 24339
rect 16044 24319 16046 24339
rect 16068 24319 16070 24339
rect 16164 24319 16166 24339
rect 16260 24319 16262 24339
rect 16284 24319 16286 24339
rect 16332 24319 16334 24339
rect 16380 24319 16382 24339
rect 16476 24319 16478 24339
rect 16548 24319 16550 24339
rect 16572 24319 16574 24339
rect 16668 24319 16670 24339
rect 16764 24319 16766 24339
rect 16812 24319 16814 24339
rect 16884 24319 16886 24339
rect 16908 24319 16910 24339
rect 17028 24319 17030 24339
rect 17124 24319 17126 24339
rect 17196 24319 17198 24339
rect 17220 24319 17222 24339
rect 17292 24319 17294 24339
rect 17316 24319 17318 24339
rect 17964 24319 17966 24339
rect 18060 24319 18062 24339
rect 18132 24319 18134 24339
rect 18228 24319 18230 24339
rect 18492 24319 18494 24339
rect 18540 24319 18542 24339
rect 18636 24319 18638 24339
rect 18732 24319 18734 24339
rect 18828 24319 18830 24339
rect 18924 24319 18926 24339
rect 18972 24319 18974 24339
rect 19020 24319 19022 24339
rect 19068 24319 19070 24339
rect 19140 24319 19142 24339
rect 19164 24319 19166 24339
rect 19236 24319 19238 24339
rect 19260 24319 19262 24339
rect 19465 24319 19499 24320
rect 19788 24319 19790 24339
rect 19836 24319 19838 24339
rect 19860 24319 19862 24339
rect 19884 24319 19886 24339
rect 19956 24319 19958 24339
rect 19980 24319 19982 24339
rect 20004 24319 20006 24339
rect 20052 24319 20054 24339
rect 20076 24319 20078 24339
rect 20100 24319 20102 24339
rect 20172 24319 20174 24339
rect 20196 24319 20198 24339
rect 20292 24319 20294 24339
rect 20388 24319 20390 24339
rect 20412 24319 20414 24339
rect 20508 24319 20510 24339
rect 20532 24319 20534 24339
rect 20604 24319 20606 24339
rect 20628 24319 20630 24339
rect 20892 24319 20894 24339
rect 20964 24319 20966 24339
rect 20988 24319 20990 24339
rect 21108 24319 21110 24339
rect 21204 24319 21206 24339
rect 21300 24319 21302 24339
rect 21324 24319 21326 24339
rect 21444 24319 21446 24339
rect 21468 24319 21470 24339
rect 21564 24319 21566 24339
rect 21588 24320 21590 24339
rect 21577 24319 21611 24320
rect -8015 24315 7685 24319
rect -7871 24295 -7837 24296
rect -7764 24295 -7762 24315
rect -7356 24295 -7354 24315
rect -7308 24295 -7306 24315
rect -7140 24295 -7138 24315
rect -6828 24295 -6826 24315
rect -6732 24295 -6730 24315
rect -6444 24295 -6442 24315
rect -6348 24295 -6346 24315
rect -6252 24295 -6250 24315
rect -5892 24295 -5890 24315
rect -5340 24295 -5338 24315
rect -4905 24312 -4891 24315
rect -4716 24295 -4714 24315
rect -4500 24295 -4498 24315
rect -4284 24295 -4282 24315
rect -3935 24295 -3877 24296
rect -3876 24295 -3874 24315
rect -3540 24295 -3538 24315
rect -3468 24295 -3466 24315
rect -3324 24295 -3322 24315
rect -3108 24295 -3106 24315
rect -3012 24295 -3010 24315
rect -2964 24295 -2962 24315
rect -2916 24295 -2914 24315
rect -2868 24295 -2866 24315
rect -2772 24295 -2770 24315
rect -2663 24295 -2605 24296
rect -2364 24295 -2362 24315
rect -1908 24295 -1906 24315
rect -1452 24295 -1450 24315
rect -1356 24295 -1354 24315
rect -1260 24295 -1258 24315
rect -1236 24295 -1234 24315
rect -1140 24295 -1138 24315
rect -876 24295 -874 24315
rect -780 24295 -778 24315
rect -564 24295 -562 24315
rect -468 24295 -466 24315
rect -12 24295 -10 24315
rect 84 24295 86 24315
rect 252 24312 254 24315
rect 252 24295 255 24312
rect 348 24295 350 24315
rect 468 24295 470 24315
rect 492 24295 494 24315
rect 564 24295 566 24315
rect 588 24295 590 24315
rect 636 24295 638 24315
rect 660 24295 662 24315
rect 732 24295 734 24315
rect 948 24295 950 24315
rect 1044 24295 1046 24315
rect 1092 24295 1094 24315
rect 1140 24295 1142 24315
rect 1308 24295 1310 24315
rect 1356 24295 1358 24315
rect 1428 24295 1430 24315
rect 1572 24295 1574 24315
rect 1860 24295 1862 24315
rect 1956 24295 1958 24315
rect 2052 24295 2054 24315
rect 2148 24295 2150 24315
rect 2244 24295 2246 24315
rect 2460 24295 2462 24315
rect 2772 24295 2774 24315
rect 2868 24295 2870 24315
rect 2940 24295 2942 24315
rect 2988 24295 2990 24315
rect 3324 24295 3326 24315
rect 3540 24295 3542 24315
rect 3660 24295 3662 24315
rect 3780 24295 3782 24315
rect 4092 24295 4094 24315
rect 4188 24295 4190 24315
rect 4308 24295 4310 24315
rect 4404 24295 4406 24315
rect 4500 24295 4502 24315
rect 4596 24295 4598 24315
rect 4692 24295 4694 24315
rect 4932 24295 4934 24315
rect 4980 24295 4982 24315
rect 5028 24295 5030 24315
rect 5124 24295 5126 24315
rect 5220 24295 5222 24315
rect 5460 24295 5462 24315
rect 5508 24295 5510 24315
rect 5556 24295 5558 24315
rect 5652 24295 5654 24315
rect 5748 24295 5750 24315
rect 5796 24295 5798 24315
rect 5844 24295 5846 24315
rect 5892 24295 5894 24315
rect 6276 24295 6278 24315
rect 6300 24295 6302 24315
rect 6372 24295 6374 24315
rect 6396 24295 6398 24315
rect 6492 24295 6494 24315
rect 6516 24295 6518 24315
rect 6588 24295 6590 24315
rect 6612 24295 6614 24315
rect 6636 24295 6638 24315
rect 6684 24295 6686 24315
rect 6708 24295 6710 24315
rect 6804 24295 6806 24315
rect 6900 24295 6902 24315
rect 7164 24295 7166 24315
rect 7236 24295 7238 24315
rect 7284 24295 7286 24315
rect 7380 24295 7382 24315
rect 7404 24295 7406 24315
rect 7476 24295 7478 24315
rect 7500 24295 7502 24315
rect 7572 24295 7574 24315
rect 7596 24295 7598 24315
rect 7668 24295 7670 24315
rect 7671 24312 7685 24315
rect 7692 24315 21611 24319
rect 7692 24312 7709 24315
rect 7692 24295 7694 24312
rect 7908 24295 7910 24315
rect 8124 24295 8126 24315
rect 8220 24295 8222 24315
rect 8652 24312 8654 24315
rect 8305 24295 8363 24296
rect 8652 24295 8655 24312
rect 8700 24295 8702 24315
rect 8748 24295 8750 24315
rect 8796 24295 8798 24315
rect 8844 24295 8846 24315
rect 8868 24295 8870 24315
rect 9516 24295 9518 24315
rect 9660 24295 9662 24315
rect 9684 24295 9686 24315
rect 9780 24295 9782 24315
rect 9804 24295 9806 24315
rect 9828 24295 9830 24315
rect 10044 24295 10046 24315
rect 10140 24295 10142 24315
rect 10236 24295 10238 24315
rect 10332 24295 10334 24315
rect 10380 24295 10382 24315
rect 10428 24295 10430 24315
rect 10524 24295 10526 24315
rect 10548 24295 10550 24315
rect 10620 24295 10622 24315
rect 10644 24295 10646 24315
rect 10716 24295 10718 24315
rect 10860 24295 10862 24315
rect 10956 24295 10958 24315
rect 11052 24295 11054 24315
rect 11100 24295 11102 24315
rect 11172 24295 11174 24315
rect 11220 24295 11222 24315
rect 11340 24295 11342 24315
rect 11436 24295 11438 24315
rect 11676 24295 11678 24315
rect 11724 24295 11726 24315
rect 11772 24295 11774 24315
rect 11796 24295 11798 24315
rect 12060 24295 12062 24315
rect 12276 24295 12278 24315
rect 12324 24295 12326 24315
rect 12372 24295 12374 24315
rect 12420 24295 12422 24315
rect 12468 24295 12470 24315
rect 12564 24295 12566 24315
rect 12721 24295 12755 24296
rect 12780 24295 12782 24315
rect 12828 24295 12830 24315
rect 12876 24295 12878 24315
rect 12972 24295 12974 24315
rect 13044 24295 13046 24315
rect 13068 24295 13070 24315
rect 13164 24295 13166 24315
rect 13332 24295 13334 24315
rect 13500 24295 13502 24315
rect 13572 24295 13574 24315
rect 13668 24295 13670 24315
rect 13716 24295 13718 24315
rect 13836 24295 13838 24315
rect 14004 24295 14006 24315
rect 14100 24295 14102 24315
rect 14940 24295 14942 24315
rect 15036 24295 15038 24315
rect 15276 24295 15278 24315
rect 15372 24295 15374 24315
rect 15420 24295 15422 24315
rect 15468 24295 15470 24315
rect 15564 24295 15566 24315
rect 15660 24295 15662 24315
rect 15732 24295 15734 24315
rect 15756 24295 15758 24315
rect 15804 24295 15806 24315
rect 15828 24295 15830 24315
rect 15852 24295 15854 24315
rect 15948 24295 15950 24315
rect 15972 24295 15974 24315
rect 16044 24295 16046 24315
rect 16068 24295 16070 24315
rect 16164 24295 16166 24315
rect 16225 24295 16259 24296
rect 16260 24295 16262 24315
rect 16284 24295 16286 24315
rect 16332 24295 16334 24315
rect 16380 24295 16382 24315
rect 16476 24295 16478 24315
rect 16548 24295 16550 24315
rect 16572 24295 16574 24315
rect 16668 24295 16670 24315
rect 16681 24295 16739 24296
rect 16764 24295 16766 24315
rect 16812 24295 16814 24315
rect 16884 24295 16886 24315
rect 16908 24295 16910 24315
rect 17028 24295 17030 24315
rect 17124 24295 17126 24315
rect 17196 24295 17198 24315
rect 17220 24295 17222 24315
rect 17292 24295 17294 24315
rect 17316 24295 17318 24315
rect 17964 24295 17966 24315
rect 18060 24295 18062 24315
rect 18132 24295 18134 24315
rect 18228 24295 18230 24315
rect 18492 24295 18494 24315
rect 18540 24295 18542 24315
rect 18636 24295 18638 24315
rect 18732 24295 18734 24315
rect 18828 24295 18830 24315
rect 18924 24295 18926 24315
rect 18972 24295 18974 24315
rect 19020 24295 19022 24315
rect 19068 24295 19070 24315
rect 19140 24295 19142 24315
rect 19164 24295 19166 24315
rect 19236 24295 19238 24315
rect 19260 24295 19262 24315
rect 19788 24295 19790 24315
rect 19836 24295 19838 24315
rect 19860 24295 19862 24315
rect 19884 24295 19886 24315
rect 19956 24295 19958 24315
rect 19980 24295 19982 24315
rect 20004 24295 20006 24315
rect 20052 24295 20054 24315
rect 20076 24295 20078 24315
rect 20100 24295 20102 24315
rect 20172 24295 20174 24315
rect 20196 24295 20198 24315
rect 20292 24295 20294 24315
rect 20388 24295 20390 24315
rect 20412 24295 20414 24315
rect 20508 24295 20510 24315
rect 20532 24295 20534 24315
rect 20604 24295 20606 24315
rect 20628 24295 20630 24315
rect 20892 24295 20894 24315
rect 20964 24295 20966 24315
rect 20988 24295 20990 24315
rect 21108 24295 21110 24315
rect 21204 24295 21206 24315
rect 21300 24295 21302 24315
rect 21324 24295 21326 24315
rect 21444 24295 21446 24315
rect 21468 24296 21470 24315
rect 21564 24296 21566 24315
rect 21577 24310 21580 24315
rect 21588 24310 21590 24315
rect 21587 24296 21590 24310
rect 21457 24295 21515 24296
rect 21553 24295 21587 24296
rect -7871 24291 -3955 24295
rect -7764 24288 -7762 24291
rect -7764 24272 -7761 24288
rect -7775 24271 -7741 24272
rect -7356 24271 -7354 24291
rect -7308 24271 -7306 24291
rect -7140 24271 -7138 24291
rect -6828 24271 -6826 24291
rect -6732 24271 -6730 24291
rect -6647 24271 -6589 24272
rect -6444 24271 -6442 24291
rect -6348 24271 -6346 24291
rect -6252 24271 -6250 24291
rect -5892 24271 -5890 24291
rect -5340 24271 -5338 24291
rect -4716 24271 -4714 24291
rect -4500 24271 -4498 24291
rect -4284 24271 -4282 24291
rect -3969 24288 -3955 24291
rect -3945 24291 8621 24295
rect -3945 24288 -3931 24291
rect -3876 24271 -3874 24291
rect -3828 24271 -3825 24288
rect -3540 24271 -3538 24291
rect -3468 24271 -3466 24291
rect -3324 24271 -3322 24291
rect -3108 24271 -3106 24291
rect -3012 24271 -3010 24291
rect -2964 24271 -2962 24291
rect -2916 24271 -2914 24291
rect -2868 24271 -2866 24291
rect -2772 24271 -2770 24291
rect -2364 24271 -2362 24291
rect -1908 24271 -1906 24291
rect -1452 24271 -1450 24291
rect -1356 24271 -1354 24291
rect -1260 24271 -1258 24291
rect -1236 24271 -1234 24291
rect -1140 24271 -1138 24291
rect -876 24271 -874 24291
rect -780 24271 -778 24291
rect -564 24271 -562 24291
rect -468 24271 -466 24291
rect -12 24271 -10 24291
rect 84 24271 86 24291
rect 231 24288 245 24291
rect 252 24288 255 24291
rect 348 24271 350 24291
rect 468 24271 470 24291
rect 492 24271 494 24291
rect 564 24271 566 24291
rect 588 24271 590 24291
rect 636 24271 638 24291
rect 660 24271 662 24291
rect 732 24271 734 24291
rect 948 24271 950 24291
rect 1044 24271 1046 24291
rect 1092 24271 1094 24291
rect 1140 24271 1142 24291
rect 1308 24271 1310 24291
rect 1356 24271 1358 24291
rect 1428 24271 1430 24291
rect 1572 24271 1574 24291
rect 1860 24271 1862 24291
rect 1956 24271 1958 24291
rect 2052 24271 2054 24291
rect 2148 24271 2150 24291
rect 2244 24271 2246 24291
rect 2460 24271 2462 24291
rect 2772 24271 2774 24291
rect 2868 24271 2870 24291
rect 2940 24271 2942 24291
rect 2988 24271 2990 24291
rect 3324 24271 3326 24291
rect 3540 24271 3542 24291
rect 3660 24271 3662 24291
rect 3780 24271 3782 24291
rect 4092 24271 4094 24291
rect 4188 24271 4190 24291
rect 4308 24271 4310 24291
rect 4404 24271 4406 24291
rect 4500 24271 4502 24291
rect 4596 24271 4598 24291
rect 4692 24271 4694 24291
rect 4932 24271 4934 24291
rect 4980 24271 4982 24291
rect 5028 24271 5030 24291
rect 5124 24271 5126 24291
rect 5220 24271 5222 24291
rect 5460 24271 5462 24291
rect 5508 24271 5510 24291
rect 5556 24271 5558 24291
rect 5652 24271 5654 24291
rect 5748 24271 5750 24291
rect 5796 24271 5798 24291
rect 5844 24271 5846 24291
rect 5892 24271 5894 24291
rect 6276 24271 6278 24291
rect 6300 24271 6302 24291
rect 6372 24271 6374 24291
rect 6396 24271 6398 24291
rect 6492 24271 6494 24291
rect 6516 24271 6518 24291
rect 6588 24271 6590 24291
rect 6612 24271 6614 24291
rect 6636 24271 6638 24291
rect 6684 24271 6686 24291
rect 6708 24271 6710 24291
rect 6804 24271 6806 24291
rect 6900 24271 6902 24291
rect 7164 24271 7166 24291
rect 7236 24271 7238 24291
rect 7284 24271 7286 24291
rect 7380 24271 7382 24291
rect 7404 24271 7406 24291
rect 7476 24271 7478 24291
rect 7500 24271 7502 24291
rect 7572 24271 7574 24291
rect 7596 24271 7598 24291
rect 7668 24271 7670 24291
rect 7692 24271 7694 24291
rect 7908 24271 7910 24291
rect 8124 24271 8126 24291
rect 8220 24271 8222 24291
rect 8305 24286 8308 24291
rect 8607 24288 8621 24291
rect 8631 24291 21587 24295
rect 8631 24288 8645 24291
rect 8652 24288 8655 24291
rect 8315 24272 8318 24286
rect 8316 24271 8318 24272
rect 8412 24271 8415 24288
rect 8700 24271 8702 24291
rect 8748 24271 8750 24291
rect 8796 24271 8798 24291
rect 8844 24271 8846 24291
rect 8868 24271 8870 24291
rect 9516 24271 9518 24291
rect 9660 24271 9662 24291
rect 9684 24271 9686 24291
rect 9780 24271 9782 24291
rect 9804 24271 9806 24291
rect 9828 24271 9830 24291
rect 10044 24271 10046 24291
rect 10140 24271 10142 24291
rect 10236 24271 10238 24291
rect 10332 24271 10334 24291
rect 10380 24271 10382 24291
rect 10428 24271 10430 24291
rect 10524 24271 10526 24291
rect 10548 24271 10550 24291
rect 10620 24271 10622 24291
rect 10644 24271 10646 24291
rect 10716 24271 10718 24291
rect 10860 24271 10862 24291
rect 10956 24271 10958 24291
rect 11052 24271 11054 24291
rect 11100 24271 11102 24291
rect 11172 24271 11174 24291
rect 11220 24271 11222 24291
rect 11340 24271 11342 24291
rect 11436 24271 11438 24291
rect 11676 24271 11678 24291
rect 11724 24271 11726 24291
rect 11772 24271 11774 24291
rect 11796 24271 11798 24291
rect 12060 24271 12062 24291
rect 12276 24271 12278 24291
rect 12324 24271 12326 24291
rect 12372 24271 12374 24291
rect 12420 24271 12422 24291
rect 12468 24271 12470 24291
rect 12564 24271 12566 24291
rect 12780 24271 12782 24291
rect 12828 24288 12830 24291
rect 12828 24271 12831 24288
rect 12876 24271 12878 24291
rect 12972 24271 12974 24291
rect 13044 24271 13046 24291
rect 13068 24271 13070 24291
rect 13164 24271 13166 24291
rect 13332 24271 13334 24291
rect 13500 24271 13502 24291
rect 13572 24271 13574 24291
rect 13668 24271 13670 24291
rect 13716 24271 13718 24291
rect 13836 24271 13838 24291
rect 14004 24271 14006 24291
rect 14100 24271 14102 24291
rect 14940 24271 14942 24291
rect 15036 24271 15038 24291
rect 15276 24271 15278 24291
rect 15372 24271 15374 24291
rect 15420 24271 15422 24291
rect 15468 24271 15470 24291
rect 15564 24271 15566 24291
rect 15660 24271 15662 24291
rect 15732 24271 15734 24291
rect 15756 24271 15758 24291
rect 15804 24271 15806 24291
rect 15828 24271 15830 24291
rect 15852 24271 15854 24291
rect 15948 24271 15950 24291
rect 15972 24271 15974 24291
rect 16044 24271 16046 24291
rect 16068 24271 16070 24291
rect 16164 24271 16166 24291
rect 16260 24271 16262 24291
rect 16284 24271 16286 24291
rect 16332 24288 16334 24291
rect 16332 24271 16335 24288
rect 16380 24271 16382 24291
rect 16476 24271 16478 24291
rect 16548 24271 16550 24291
rect 16572 24271 16574 24291
rect 16668 24271 16670 24291
rect 16681 24286 16684 24291
rect 16691 24272 16694 24286
rect 16692 24271 16694 24272
rect 16764 24271 16766 24291
rect 16812 24288 16814 24291
rect 16788 24271 16791 24288
rect 16812 24271 16815 24288
rect 16884 24271 16886 24291
rect 16908 24271 16910 24291
rect 17028 24271 17030 24291
rect 17124 24271 17126 24291
rect 17196 24271 17198 24291
rect 17220 24271 17222 24291
rect 17292 24271 17294 24291
rect 17316 24271 17318 24291
rect 17964 24271 17966 24291
rect 18060 24271 18062 24291
rect 18132 24271 18134 24291
rect 18228 24271 18230 24291
rect 18492 24271 18494 24291
rect 18540 24271 18542 24291
rect 18636 24271 18638 24291
rect 18732 24271 18734 24291
rect 18828 24271 18830 24291
rect 18924 24271 18926 24291
rect 18972 24271 18974 24291
rect 19020 24271 19022 24291
rect 19068 24271 19070 24291
rect 19140 24271 19142 24291
rect 19164 24271 19166 24291
rect 19236 24271 19238 24291
rect 19260 24271 19262 24291
rect 19551 24288 19565 24291
rect 19788 24271 19790 24291
rect 19836 24271 19838 24291
rect 19860 24271 19862 24291
rect 19884 24271 19886 24291
rect 19956 24271 19958 24291
rect 19980 24271 19982 24291
rect 20004 24271 20006 24291
rect 20052 24271 20054 24291
rect 20076 24271 20078 24291
rect 20100 24271 20102 24291
rect 20172 24271 20174 24291
rect 20196 24271 20198 24291
rect 20292 24271 20294 24291
rect 20388 24271 20390 24291
rect 20412 24271 20414 24291
rect 20508 24271 20510 24291
rect 20532 24271 20534 24291
rect 20604 24271 20606 24291
rect 20628 24271 20630 24291
rect 20892 24271 20894 24291
rect 20964 24271 20966 24291
rect 20988 24271 20990 24291
rect 21108 24271 21110 24291
rect 21204 24271 21206 24291
rect 21300 24271 21302 24291
rect 21324 24271 21326 24291
rect 21444 24272 21446 24291
rect 21457 24286 21460 24291
rect 21468 24286 21470 24291
rect 21553 24286 21556 24291
rect 21564 24288 21566 24291
rect 21564 24286 21567 24288
rect 21467 24272 21470 24286
rect 21563 24278 21567 24286
rect 21577 24278 21581 24286
rect 21563 24272 21577 24278
rect 21433 24271 21467 24272
rect -7775 24267 -3835 24271
rect -7775 24264 -7771 24267
rect -7764 24264 -7761 24267
rect -7655 24247 -7621 24248
rect -7356 24247 -7354 24267
rect -7308 24248 -7306 24267
rect -7319 24247 -7285 24248
rect -7655 24243 -7285 24247
rect -7247 24247 -7213 24248
rect -7140 24247 -7138 24267
rect -6828 24247 -6826 24267
rect -6732 24247 -6730 24267
rect -6647 24262 -6644 24267
rect -6637 24248 -6634 24262
rect -6636 24247 -6634 24248
rect -6540 24247 -6537 24264
rect -6444 24247 -6442 24267
rect -6348 24247 -6346 24267
rect -6252 24247 -6250 24267
rect -5892 24247 -5890 24267
rect -5340 24247 -5338 24267
rect -4716 24247 -4714 24267
rect -4500 24247 -4498 24267
rect -4284 24247 -4282 24267
rect -3876 24247 -3874 24267
rect -3849 24264 -3835 24267
rect -3828 24267 -2563 24271
rect -3828 24264 -3811 24267
rect -3828 24247 -3826 24264
rect -3540 24247 -3538 24267
rect -3468 24247 -3466 24267
rect -3324 24247 -3322 24267
rect -3108 24247 -3106 24267
rect -3012 24247 -3010 24267
rect -2964 24247 -2962 24267
rect -2916 24247 -2914 24267
rect -2868 24247 -2866 24267
rect -2772 24247 -2770 24267
rect -2577 24264 -2563 24267
rect -2553 24267 8405 24271
rect -2553 24264 -2539 24267
rect -2364 24247 -2362 24267
rect -1908 24247 -1906 24267
rect -1452 24247 -1450 24267
rect -1356 24247 -1354 24267
rect -1260 24247 -1258 24267
rect -1236 24247 -1234 24267
rect -1140 24247 -1138 24267
rect -876 24247 -874 24267
rect -780 24247 -778 24267
rect -564 24247 -562 24267
rect -468 24247 -466 24267
rect -12 24247 -10 24267
rect 84 24247 86 24267
rect 348 24247 350 24267
rect 468 24247 470 24267
rect 492 24247 494 24267
rect 564 24247 566 24267
rect 588 24247 590 24267
rect 636 24247 638 24267
rect 660 24247 662 24267
rect 732 24247 734 24267
rect 948 24247 950 24267
rect 1044 24247 1046 24267
rect 1092 24247 1094 24267
rect 1140 24247 1142 24267
rect 1308 24247 1310 24267
rect 1356 24247 1358 24267
rect 1428 24247 1430 24267
rect 1572 24247 1574 24267
rect 1860 24247 1862 24267
rect 1956 24247 1958 24267
rect 2052 24247 2054 24267
rect 2148 24247 2150 24267
rect 2244 24247 2246 24267
rect 2460 24247 2462 24267
rect 2772 24247 2774 24267
rect 2868 24247 2870 24267
rect 2940 24247 2942 24267
rect 2988 24247 2990 24267
rect 3324 24247 3326 24267
rect 3540 24247 3542 24267
rect 3660 24247 3662 24267
rect 3780 24247 3782 24267
rect 4092 24247 4094 24267
rect 4188 24247 4190 24267
rect 4308 24247 4310 24267
rect 4404 24247 4406 24267
rect 4500 24247 4502 24267
rect 4596 24247 4598 24267
rect 4692 24247 4694 24267
rect 4932 24247 4934 24267
rect 4980 24247 4982 24267
rect 5028 24247 5030 24267
rect 5124 24247 5126 24267
rect 5220 24247 5222 24267
rect 5460 24247 5462 24267
rect 5508 24247 5510 24267
rect 5556 24247 5558 24267
rect 5652 24247 5654 24267
rect 5748 24247 5750 24267
rect 5796 24247 5798 24267
rect 5844 24247 5846 24267
rect 5892 24247 5894 24267
rect 6276 24247 6278 24267
rect 6300 24247 6302 24267
rect 6372 24247 6374 24267
rect 6396 24247 6398 24267
rect 6492 24247 6494 24267
rect 6516 24247 6518 24267
rect 6588 24247 6590 24267
rect 6612 24247 6614 24267
rect 6636 24247 6638 24267
rect 6684 24247 6686 24267
rect 6708 24247 6710 24267
rect 6804 24247 6806 24267
rect 6900 24247 6902 24267
rect 7164 24247 7166 24267
rect 7236 24247 7238 24267
rect 7284 24247 7286 24267
rect 7380 24247 7382 24267
rect 7404 24247 7406 24267
rect 7476 24247 7478 24267
rect 7500 24247 7502 24267
rect 7572 24247 7574 24267
rect 7596 24247 7598 24267
rect 7668 24247 7670 24267
rect 7692 24247 7694 24267
rect 7908 24247 7910 24267
rect 8124 24247 8126 24267
rect 8220 24247 8222 24267
rect 8316 24247 8318 24267
rect 8391 24264 8405 24267
rect 8412 24267 16781 24271
rect 8412 24264 8429 24267
rect 8412 24247 8414 24264
rect 8700 24247 8702 24267
rect 8748 24247 8750 24267
rect 8796 24247 8798 24267
rect 8844 24247 8846 24267
rect 8868 24247 8870 24267
rect 9516 24247 9518 24267
rect 9660 24247 9662 24267
rect 9684 24247 9686 24267
rect 9780 24247 9782 24267
rect 9804 24247 9806 24267
rect 9828 24247 9830 24267
rect 10044 24247 10046 24267
rect 10140 24247 10142 24267
rect 10236 24247 10238 24267
rect 10332 24247 10334 24267
rect 10380 24247 10382 24267
rect 10428 24247 10430 24267
rect 10524 24247 10526 24267
rect 10548 24247 10550 24267
rect 10620 24247 10622 24267
rect 10644 24247 10646 24267
rect 10716 24247 10718 24267
rect 10860 24247 10862 24267
rect 10956 24247 10958 24267
rect 11052 24247 11054 24267
rect 11100 24247 11102 24267
rect 11172 24247 11174 24267
rect 11220 24247 11222 24267
rect 11340 24247 11342 24267
rect 11436 24247 11438 24267
rect 11676 24247 11678 24267
rect 11724 24247 11726 24267
rect 11772 24247 11774 24267
rect 11796 24247 11798 24267
rect 12060 24247 12062 24267
rect 12276 24247 12278 24267
rect 12324 24247 12326 24267
rect 12372 24247 12374 24267
rect 12420 24247 12422 24267
rect 12468 24247 12470 24267
rect 12564 24247 12566 24267
rect 12780 24247 12782 24267
rect 12807 24264 12821 24267
rect 12828 24264 12831 24267
rect 12876 24247 12878 24267
rect 12972 24247 12974 24267
rect 13044 24247 13046 24267
rect 13068 24247 13070 24267
rect 13164 24247 13166 24267
rect 13332 24247 13334 24267
rect 13500 24247 13502 24267
rect 13572 24247 13574 24267
rect 13668 24247 13670 24267
rect 13716 24247 13718 24267
rect 13836 24247 13838 24267
rect 14004 24247 14006 24267
rect 14100 24247 14102 24267
rect 14940 24247 14942 24267
rect 15036 24247 15038 24267
rect 15276 24247 15278 24267
rect 15372 24247 15374 24267
rect 15420 24247 15422 24267
rect 15468 24247 15470 24267
rect 15564 24247 15566 24267
rect 15660 24247 15662 24267
rect 15732 24247 15734 24267
rect 15756 24247 15758 24267
rect 15804 24247 15806 24267
rect 15828 24247 15830 24267
rect 15852 24247 15854 24267
rect 15948 24247 15950 24267
rect 15972 24247 15974 24267
rect 16044 24247 16046 24267
rect 16068 24247 16070 24267
rect 16164 24247 16166 24267
rect 16260 24247 16262 24267
rect 16284 24247 16286 24267
rect 16311 24264 16325 24267
rect 16332 24264 16335 24267
rect 16380 24247 16382 24267
rect 16476 24247 16478 24267
rect 16548 24247 16550 24267
rect 16572 24247 16574 24267
rect 16668 24247 16670 24267
rect 16692 24247 16694 24267
rect 16764 24247 16766 24267
rect 16767 24264 16781 24267
rect 16788 24267 21467 24271
rect 16788 24264 16805 24267
rect 16812 24264 16815 24267
rect 16788 24247 16790 24264
rect 16884 24247 16886 24267
rect 16908 24247 16910 24267
rect 17028 24247 17030 24267
rect 17124 24247 17126 24267
rect 17196 24247 17198 24267
rect 17220 24247 17222 24267
rect 17292 24247 17294 24267
rect 17316 24247 17318 24267
rect 17964 24247 17966 24267
rect 18060 24247 18062 24267
rect 18132 24247 18134 24267
rect 18228 24247 18230 24267
rect 18492 24247 18494 24267
rect 18540 24247 18542 24267
rect 18636 24247 18638 24267
rect 18732 24247 18734 24267
rect 18828 24247 18830 24267
rect 18924 24247 18926 24267
rect 18972 24247 18974 24267
rect 19020 24247 19022 24267
rect 19068 24247 19070 24267
rect 19140 24247 19142 24267
rect 19164 24247 19166 24267
rect 19236 24247 19238 24267
rect 19260 24247 19262 24267
rect 19788 24247 19790 24267
rect 19836 24247 19838 24267
rect 19860 24247 19862 24267
rect 19884 24247 19886 24267
rect 19956 24247 19958 24267
rect 19980 24247 19982 24267
rect 20004 24247 20006 24267
rect 20052 24247 20054 24267
rect 20076 24247 20078 24267
rect 20100 24247 20102 24267
rect 20172 24247 20174 24267
rect 20196 24247 20198 24267
rect 20292 24247 20294 24267
rect 20388 24247 20390 24267
rect 20412 24247 20414 24267
rect 20508 24247 20510 24267
rect 20532 24247 20534 24267
rect 20604 24247 20606 24267
rect 20628 24247 20630 24267
rect 20892 24247 20894 24267
rect 20964 24247 20966 24267
rect 20988 24247 20990 24267
rect 21108 24247 21110 24267
rect 21204 24247 21206 24267
rect 21300 24247 21302 24267
rect 21324 24247 21326 24267
rect 21433 24262 21436 24267
rect 21444 24262 21446 24267
rect 21443 24248 21446 24262
rect 21361 24247 21395 24248
rect -7247 24243 -6547 24247
rect -7356 24224 -7354 24243
rect -7319 24238 -7316 24243
rect -7308 24238 -7306 24243
rect -7140 24240 -7138 24243
rect -7309 24224 -7306 24238
rect -7223 24230 -7219 24238
rect -7233 24224 -7223 24230
rect -7140 24224 -7137 24240
rect -7535 24223 -7501 24224
rect -7463 24223 -7429 24224
rect -7535 24219 -7429 24223
rect -7415 24223 -7381 24224
rect -7367 24223 -7333 24224
rect -7415 24219 -7333 24223
rect -7151 24223 -7117 24224
rect -6828 24223 -6826 24243
rect -6732 24223 -6730 24243
rect -6636 24223 -6634 24243
rect -6561 24240 -6547 24243
rect -6540 24243 21395 24247
rect -6540 24240 -6523 24243
rect -6540 24223 -6538 24240
rect -6444 24223 -6442 24243
rect -6348 24223 -6346 24243
rect -6252 24223 -6250 24243
rect -5892 24223 -5890 24243
rect -5340 24223 -5338 24243
rect -4716 24223 -4714 24243
rect -4500 24223 -4498 24243
rect -4284 24223 -4282 24243
rect -3876 24223 -3874 24243
rect -3828 24223 -3826 24243
rect -3540 24223 -3538 24243
rect -3468 24223 -3466 24243
rect -3324 24223 -3322 24243
rect -3108 24223 -3106 24243
rect -3095 24223 -3037 24224
rect -3012 24223 -3010 24243
rect -2964 24223 -2962 24243
rect -2916 24223 -2914 24243
rect -2868 24223 -2866 24243
rect -2772 24223 -2770 24243
rect -2364 24223 -2362 24243
rect -1908 24223 -1906 24243
rect -1452 24223 -1450 24243
rect -1356 24223 -1354 24243
rect -1260 24223 -1258 24243
rect -1236 24223 -1234 24243
rect -1140 24223 -1138 24243
rect -876 24223 -874 24243
rect -815 24223 -781 24224
rect -780 24223 -778 24243
rect -564 24223 -562 24243
rect -468 24223 -466 24243
rect -12 24223 -10 24243
rect 84 24223 86 24243
rect 348 24223 350 24243
rect 468 24223 470 24243
rect 492 24223 494 24243
rect 564 24223 566 24243
rect 588 24223 590 24243
rect 636 24223 638 24243
rect 660 24223 662 24243
rect 732 24223 734 24243
rect 948 24223 950 24243
rect 1044 24223 1046 24243
rect 1092 24223 1094 24243
rect 1140 24223 1142 24243
rect 1308 24223 1310 24243
rect 1356 24223 1358 24243
rect 1428 24223 1430 24243
rect 1572 24223 1574 24243
rect 1860 24223 1862 24243
rect 1956 24223 1958 24243
rect 2052 24223 2054 24243
rect 2148 24223 2150 24243
rect 2244 24223 2246 24243
rect 2460 24223 2462 24243
rect 2772 24223 2774 24243
rect 2868 24223 2870 24243
rect 2940 24223 2942 24243
rect 2988 24223 2990 24243
rect 3324 24223 3326 24243
rect 3540 24223 3542 24243
rect 3660 24223 3662 24243
rect 3780 24223 3782 24243
rect 4092 24223 4094 24243
rect 4188 24223 4190 24243
rect 4308 24223 4310 24243
rect 4404 24223 4406 24243
rect 4500 24223 4502 24243
rect 4596 24223 4598 24243
rect 4692 24223 4694 24243
rect 4932 24223 4934 24243
rect 4980 24223 4982 24243
rect 5028 24223 5030 24243
rect 5124 24223 5126 24243
rect 5220 24223 5222 24243
rect 5460 24223 5462 24243
rect 5508 24223 5510 24243
rect 5556 24223 5558 24243
rect 5652 24223 5654 24243
rect 5748 24223 5750 24243
rect 5796 24223 5798 24243
rect 5844 24223 5846 24243
rect 5892 24223 5894 24243
rect 6276 24223 6278 24243
rect 6300 24223 6302 24243
rect 6372 24223 6374 24243
rect 6396 24223 6398 24243
rect 6492 24223 6494 24243
rect 6516 24223 6518 24243
rect 6588 24223 6590 24243
rect 6612 24223 6614 24243
rect 6636 24223 6638 24243
rect 6684 24223 6686 24243
rect 6708 24223 6710 24243
rect 6804 24223 6806 24243
rect 6900 24223 6902 24243
rect 7164 24223 7166 24243
rect 7236 24223 7238 24243
rect 7284 24223 7286 24243
rect 7380 24223 7382 24243
rect 7404 24223 7406 24243
rect 7476 24223 7478 24243
rect 7500 24223 7502 24243
rect 7572 24223 7574 24243
rect 7596 24223 7598 24243
rect 7668 24223 7670 24243
rect 7692 24223 7694 24243
rect 7908 24223 7910 24243
rect 8124 24223 8126 24243
rect 8220 24223 8222 24243
rect 8316 24223 8318 24243
rect 8412 24223 8414 24243
rect 8700 24223 8702 24243
rect 8748 24223 8750 24243
rect 8796 24223 8798 24243
rect 8844 24223 8846 24243
rect 8868 24223 8870 24243
rect 9516 24223 9518 24243
rect 9660 24223 9662 24243
rect 9684 24223 9686 24243
rect 9780 24223 9782 24243
rect 9804 24223 9806 24243
rect 9828 24223 9830 24243
rect 10044 24223 10046 24243
rect 10140 24223 10142 24243
rect 10236 24223 10238 24243
rect 10332 24223 10334 24243
rect 10380 24223 10382 24243
rect 10428 24223 10430 24243
rect 10524 24223 10526 24243
rect 10548 24223 10550 24243
rect 10620 24223 10622 24243
rect 10644 24223 10646 24243
rect 10716 24223 10718 24243
rect 10860 24223 10862 24243
rect 10956 24223 10958 24243
rect 11052 24223 11054 24243
rect 11100 24223 11102 24243
rect 11172 24223 11174 24243
rect 11220 24223 11222 24243
rect 11340 24223 11342 24243
rect 11436 24223 11438 24243
rect 11676 24223 11678 24243
rect 11724 24223 11726 24243
rect 11772 24223 11774 24243
rect 11796 24223 11798 24243
rect 12060 24223 12062 24243
rect 12276 24223 12278 24243
rect 12324 24223 12326 24243
rect 12372 24223 12374 24243
rect 12420 24223 12422 24243
rect 12468 24223 12470 24243
rect 12564 24223 12566 24243
rect 12780 24223 12782 24243
rect 12876 24223 12878 24243
rect 12972 24223 12974 24243
rect 13044 24223 13046 24243
rect 13068 24223 13070 24243
rect 13164 24223 13166 24243
rect 13332 24223 13334 24243
rect 13500 24223 13502 24243
rect 13572 24223 13574 24243
rect 13668 24223 13670 24243
rect 13716 24223 13718 24243
rect 13836 24223 13838 24243
rect 14004 24223 14006 24243
rect 14100 24223 14102 24243
rect 14940 24223 14942 24243
rect 15036 24223 15038 24243
rect 15276 24223 15278 24243
rect 15372 24223 15374 24243
rect 15420 24223 15422 24243
rect 15468 24223 15470 24243
rect 15564 24223 15566 24243
rect 15660 24223 15662 24243
rect 15732 24223 15734 24243
rect 15756 24223 15758 24243
rect 15804 24223 15806 24243
rect 15828 24223 15830 24243
rect 15852 24223 15854 24243
rect 15948 24223 15950 24243
rect 15972 24223 15974 24243
rect 16044 24223 16046 24243
rect 16068 24223 16070 24243
rect 16164 24223 16166 24243
rect 16260 24223 16262 24243
rect 16284 24223 16286 24243
rect 16380 24223 16382 24243
rect 16476 24223 16478 24243
rect 16548 24223 16550 24243
rect 16572 24223 16574 24243
rect 16668 24223 16670 24243
rect 16692 24223 16694 24243
rect 16764 24223 16766 24243
rect 16788 24223 16790 24243
rect 16884 24223 16886 24243
rect 16908 24223 16910 24243
rect 17028 24223 17030 24243
rect 17124 24223 17126 24243
rect 17196 24223 17198 24243
rect 17220 24223 17222 24243
rect 17292 24223 17294 24243
rect 17316 24223 17318 24243
rect 17964 24223 17966 24243
rect 18060 24223 18062 24243
rect 18132 24223 18134 24243
rect 18228 24223 18230 24243
rect 18492 24223 18494 24243
rect 18540 24223 18542 24243
rect 18636 24223 18638 24243
rect 18732 24223 18734 24243
rect 18828 24223 18830 24243
rect 18924 24223 18926 24243
rect 18972 24223 18974 24243
rect 19020 24223 19022 24243
rect 19068 24223 19070 24243
rect 19140 24223 19142 24243
rect 19164 24223 19166 24243
rect 19236 24223 19238 24243
rect 19260 24223 19262 24243
rect 19788 24223 19790 24243
rect 19836 24223 19838 24243
rect 19860 24223 19862 24243
rect 19884 24223 19886 24243
rect 19956 24223 19958 24243
rect 19980 24223 19982 24243
rect 20004 24223 20006 24243
rect 20052 24223 20054 24243
rect 20076 24223 20078 24243
rect 20100 24223 20102 24243
rect 20172 24223 20174 24243
rect 20196 24223 20198 24243
rect 20292 24223 20294 24243
rect 20388 24223 20390 24243
rect 20412 24223 20414 24243
rect 20508 24223 20510 24243
rect 20532 24223 20534 24243
rect 20604 24223 20606 24243
rect 20628 24223 20630 24243
rect 20892 24223 20894 24243
rect 20964 24223 20966 24243
rect 20988 24223 20990 24243
rect 21108 24223 21110 24243
rect 21204 24223 21206 24243
rect 21300 24223 21302 24243
rect 21324 24223 21326 24243
rect 21337 24223 21371 24224
rect -7151 24219 21371 24223
rect -7367 24214 -7364 24219
rect -7356 24216 -7354 24219
rect -7151 24216 -7147 24219
rect -7140 24216 -7137 24219
rect -7356 24214 -7353 24216
rect -7439 24206 -7435 24214
rect -7449 24200 -7439 24206
rect -7357 24200 -7353 24214
rect -6828 24200 -6826 24219
rect -6935 24199 -6901 24200
rect -6863 24199 -6805 24200
rect -6732 24199 -6730 24219
rect -6636 24199 -6634 24219
rect -6540 24199 -6538 24219
rect -6444 24199 -6442 24219
rect -6348 24199 -6346 24219
rect -6252 24199 -6250 24219
rect -5892 24199 -5890 24219
rect -5340 24199 -5338 24219
rect -4716 24199 -4714 24219
rect -4500 24199 -4498 24219
rect -4284 24199 -4282 24219
rect -3876 24199 -3874 24219
rect -3828 24199 -3826 24219
rect -3540 24199 -3538 24219
rect -3468 24199 -3466 24219
rect -3324 24199 -3322 24219
rect -3108 24199 -3106 24219
rect -3012 24199 -3010 24219
rect -2964 24216 -2962 24219
rect -2988 24199 -2985 24216
rect -2964 24199 -2961 24216
rect -2916 24199 -2914 24219
rect -2868 24199 -2866 24219
rect -2772 24199 -2770 24219
rect -2364 24199 -2362 24219
rect -1908 24199 -1906 24219
rect -1452 24199 -1450 24219
rect -1356 24199 -1354 24219
rect -1260 24199 -1258 24219
rect -1236 24199 -1234 24219
rect -1140 24199 -1138 24219
rect -876 24199 -874 24219
rect -780 24199 -778 24219
rect -564 24199 -562 24219
rect -468 24199 -466 24219
rect -12 24199 -10 24219
rect 84 24199 86 24219
rect 348 24199 350 24219
rect 468 24199 470 24219
rect 492 24199 494 24219
rect 564 24199 566 24219
rect 588 24199 590 24219
rect 636 24199 638 24219
rect 660 24199 662 24219
rect 732 24199 734 24219
rect 948 24199 950 24219
rect 1044 24199 1046 24219
rect 1092 24199 1094 24219
rect 1140 24199 1142 24219
rect 1308 24199 1310 24219
rect 1356 24199 1358 24219
rect 1428 24199 1430 24219
rect 1572 24199 1574 24219
rect 1860 24199 1862 24219
rect 1956 24199 1958 24219
rect 2052 24199 2054 24219
rect 2148 24199 2150 24219
rect 2244 24199 2246 24219
rect 2460 24199 2462 24219
rect 2772 24199 2774 24219
rect 2868 24199 2870 24219
rect 2940 24199 2942 24219
rect 2988 24199 2990 24219
rect 3324 24199 3326 24219
rect 3540 24199 3542 24219
rect 3660 24199 3662 24219
rect 3780 24199 3782 24219
rect 4092 24199 4094 24219
rect 4188 24199 4190 24219
rect 4308 24199 4310 24219
rect 4404 24199 4406 24219
rect 4500 24199 4502 24219
rect 4596 24199 4598 24219
rect 4692 24199 4694 24219
rect 4932 24199 4934 24219
rect 4980 24199 4982 24219
rect 5028 24199 5030 24219
rect 5124 24199 5126 24219
rect 5220 24199 5222 24219
rect 5460 24199 5462 24219
rect 5508 24199 5510 24219
rect 5556 24199 5558 24219
rect 5652 24199 5654 24219
rect 5748 24199 5750 24219
rect 5796 24199 5798 24219
rect 5844 24199 5846 24219
rect 5892 24199 5894 24219
rect 6276 24199 6278 24219
rect 6300 24199 6302 24219
rect 6372 24199 6374 24219
rect 6396 24199 6398 24219
rect 6492 24199 6494 24219
rect 6516 24199 6518 24219
rect 6588 24199 6590 24219
rect 6612 24199 6614 24219
rect 6636 24199 6638 24219
rect 6684 24199 6686 24219
rect 6708 24199 6710 24219
rect 6804 24199 6806 24219
rect 6900 24199 6902 24219
rect 7164 24199 7166 24219
rect 7236 24199 7238 24219
rect 7284 24199 7286 24219
rect 7380 24199 7382 24219
rect 7404 24199 7406 24219
rect 7476 24199 7478 24219
rect 7500 24199 7502 24219
rect 7572 24199 7574 24219
rect 7596 24199 7598 24219
rect 7668 24199 7670 24219
rect 7692 24199 7694 24219
rect 7908 24199 7910 24219
rect 8124 24199 8126 24219
rect 8220 24199 8222 24219
rect 8316 24199 8318 24219
rect 8412 24199 8414 24219
rect 8700 24199 8702 24219
rect 8748 24199 8750 24219
rect 8796 24199 8798 24219
rect 8844 24199 8846 24219
rect 8868 24199 8870 24219
rect 9516 24199 9518 24219
rect 9660 24199 9662 24219
rect 9684 24199 9686 24219
rect 9780 24199 9782 24219
rect 9804 24199 9806 24219
rect 9828 24199 9830 24219
rect 10044 24199 10046 24219
rect 10140 24199 10142 24219
rect 10236 24199 10238 24219
rect 10332 24199 10334 24219
rect 10380 24199 10382 24219
rect 10428 24199 10430 24219
rect 10524 24199 10526 24219
rect 10548 24199 10550 24219
rect 10620 24199 10622 24219
rect 10644 24199 10646 24219
rect 10716 24199 10718 24219
rect 10860 24199 10862 24219
rect 10956 24199 10958 24219
rect 11052 24199 11054 24219
rect 11100 24199 11102 24219
rect 11172 24199 11174 24219
rect 11220 24199 11222 24219
rect 11340 24199 11342 24219
rect 11436 24199 11438 24219
rect 11676 24199 11678 24219
rect 11724 24199 11726 24219
rect 11772 24199 11774 24219
rect 11796 24199 11798 24219
rect 12060 24199 12062 24219
rect 12276 24199 12278 24219
rect 12324 24199 12326 24219
rect 12372 24199 12374 24219
rect 12420 24199 12422 24219
rect 12468 24199 12470 24219
rect 12564 24199 12566 24219
rect 12780 24199 12782 24219
rect 12876 24199 12878 24219
rect 12972 24199 12974 24219
rect 13044 24199 13046 24219
rect 13068 24199 13070 24219
rect 13164 24199 13166 24219
rect 13332 24199 13334 24219
rect 13500 24199 13502 24219
rect 13572 24199 13574 24219
rect 13668 24199 13670 24219
rect 13716 24199 13718 24219
rect 13836 24199 13838 24219
rect 13921 24199 13979 24200
rect 14004 24199 14006 24219
rect 14100 24199 14102 24219
rect 14940 24199 14942 24219
rect 15036 24199 15038 24219
rect 15276 24199 15278 24219
rect 15372 24199 15374 24219
rect 15420 24199 15422 24219
rect 15468 24199 15470 24219
rect 15564 24199 15566 24219
rect 15660 24199 15662 24219
rect 15732 24199 15734 24219
rect 15756 24199 15758 24219
rect 15804 24199 15806 24219
rect 15828 24199 15830 24219
rect 15852 24199 15854 24219
rect 15948 24199 15950 24219
rect 15972 24199 15974 24219
rect 16044 24199 16046 24219
rect 16068 24199 16070 24219
rect 16164 24199 16166 24219
rect 16260 24199 16262 24219
rect 16284 24199 16286 24219
rect 16380 24199 16382 24219
rect 16476 24199 16478 24219
rect 16548 24199 16550 24219
rect 16572 24199 16574 24219
rect 16668 24199 16670 24219
rect 16692 24199 16694 24219
rect 16764 24199 16766 24219
rect 16788 24199 16790 24219
rect 16884 24199 16886 24219
rect 16908 24199 16910 24219
rect 17028 24199 17030 24219
rect 17124 24199 17126 24219
rect 17196 24199 17198 24219
rect 17220 24199 17222 24219
rect 17292 24199 17294 24219
rect 17316 24199 17318 24219
rect 17964 24199 17966 24219
rect 18060 24199 18062 24219
rect 18132 24199 18134 24219
rect 18228 24199 18230 24219
rect 18492 24199 18494 24219
rect 18540 24199 18542 24219
rect 18636 24199 18638 24219
rect 18732 24199 18734 24219
rect 18828 24199 18830 24219
rect 18924 24199 18926 24219
rect 18972 24199 18974 24219
rect 19020 24199 19022 24219
rect 19068 24199 19070 24219
rect 19140 24199 19142 24219
rect 19164 24199 19166 24219
rect 19236 24199 19238 24219
rect 19260 24199 19262 24219
rect 19788 24199 19790 24219
rect 19836 24199 19838 24219
rect 19860 24199 19862 24219
rect 19884 24199 19886 24219
rect 19956 24199 19958 24219
rect 19980 24199 19982 24219
rect 20004 24199 20006 24219
rect 20052 24199 20054 24219
rect 20076 24199 20078 24219
rect 20100 24199 20102 24219
rect 20172 24199 20174 24219
rect 20196 24199 20198 24219
rect 20292 24199 20294 24219
rect 20388 24199 20390 24219
rect 20412 24199 20414 24219
rect 20508 24199 20510 24219
rect 20532 24199 20534 24219
rect 20604 24199 20606 24219
rect 20628 24199 20630 24219
rect 20892 24199 20894 24219
rect 20964 24199 20966 24219
rect 20988 24199 20990 24219
rect 21108 24199 21110 24219
rect 21204 24199 21206 24219
rect 21300 24199 21302 24219
rect 21324 24200 21326 24219
rect 21313 24199 21347 24200
rect -6935 24195 -2995 24199
rect -6839 24190 -6836 24195
rect -6828 24192 -6826 24195
rect -6732 24192 -6730 24195
rect -6828 24190 -6825 24192
rect -6839 24182 -6835 24190
rect -6849 24176 -6839 24182
rect -6829 24176 -6825 24190
rect -6732 24176 -6729 24192
rect -6636 24176 -6634 24195
rect -6743 24175 -6709 24176
rect -6671 24175 -6613 24176
rect -6540 24175 -6538 24195
rect -6444 24175 -6442 24195
rect -6348 24175 -6346 24195
rect -6252 24175 -6250 24195
rect -5892 24175 -5890 24195
rect -5615 24175 -5581 24176
rect -5340 24175 -5338 24195
rect -4716 24175 -4714 24195
rect -4500 24175 -4498 24195
rect -4284 24175 -4282 24195
rect -3876 24175 -3874 24195
rect -3828 24175 -3826 24195
rect -3540 24175 -3538 24195
rect -3468 24175 -3466 24195
rect -3324 24175 -3322 24195
rect -3108 24175 -3106 24195
rect -3012 24175 -3010 24195
rect -3009 24192 -2995 24195
rect -2988 24195 21347 24199
rect -2988 24192 -2971 24195
rect -2964 24192 -2961 24195
rect -2988 24175 -2986 24192
rect -2916 24175 -2914 24195
rect -2868 24175 -2866 24195
rect -2772 24175 -2770 24195
rect -2364 24175 -2362 24195
rect -1908 24175 -1906 24195
rect -1452 24175 -1450 24195
rect -1356 24175 -1354 24195
rect -1260 24175 -1258 24195
rect -1236 24175 -1234 24195
rect -1140 24175 -1138 24195
rect -876 24175 -874 24195
rect -780 24175 -778 24195
rect -729 24192 -715 24195
rect -564 24175 -562 24195
rect -468 24175 -466 24195
rect -12 24175 -10 24195
rect 84 24175 86 24195
rect 348 24175 350 24195
rect 468 24175 470 24195
rect 492 24175 494 24195
rect 564 24175 566 24195
rect 588 24175 590 24195
rect 636 24175 638 24195
rect 660 24175 662 24195
rect 732 24175 734 24195
rect 948 24175 950 24195
rect 1044 24175 1046 24195
rect 1092 24175 1094 24195
rect 1140 24175 1142 24195
rect 1308 24175 1310 24195
rect 1356 24175 1358 24195
rect 1428 24175 1430 24195
rect 1572 24175 1574 24195
rect 1860 24175 1862 24195
rect 1956 24175 1958 24195
rect 2052 24175 2054 24195
rect 2148 24175 2150 24195
rect 2244 24175 2246 24195
rect 2460 24175 2462 24195
rect 2772 24175 2774 24195
rect 2868 24175 2870 24195
rect 2940 24175 2942 24195
rect 2988 24175 2990 24195
rect 3324 24175 3326 24195
rect 3540 24175 3542 24195
rect 3660 24175 3662 24195
rect 3780 24175 3782 24195
rect 4092 24175 4094 24195
rect 4188 24175 4190 24195
rect 4308 24175 4310 24195
rect 4404 24175 4406 24195
rect 4500 24175 4502 24195
rect 4596 24175 4598 24195
rect 4692 24175 4694 24195
rect 4932 24175 4934 24195
rect 4980 24175 4982 24195
rect 5028 24175 5030 24195
rect 5124 24175 5126 24195
rect 5220 24175 5222 24195
rect 5460 24175 5462 24195
rect 5508 24175 5510 24195
rect 5556 24175 5558 24195
rect 5652 24175 5654 24195
rect 5748 24175 5750 24195
rect 5796 24175 5798 24195
rect 5844 24175 5846 24195
rect 5892 24175 5894 24195
rect 6276 24175 6278 24195
rect 6300 24175 6302 24195
rect 6372 24175 6374 24195
rect 6396 24175 6398 24195
rect 6492 24175 6494 24195
rect 6516 24175 6518 24195
rect 6588 24175 6590 24195
rect 6612 24175 6614 24195
rect 6636 24175 6638 24195
rect 6684 24175 6686 24195
rect 6708 24175 6710 24195
rect 6804 24175 6806 24195
rect 6900 24175 6902 24195
rect 7164 24175 7166 24195
rect 7236 24175 7238 24195
rect 7284 24175 7286 24195
rect 7380 24175 7382 24195
rect 7404 24175 7406 24195
rect 7476 24175 7478 24195
rect 7500 24175 7502 24195
rect 7572 24175 7574 24195
rect 7596 24175 7598 24195
rect 7668 24175 7670 24195
rect 7692 24175 7694 24195
rect 7908 24175 7910 24195
rect 8124 24175 8126 24195
rect 8220 24175 8222 24195
rect 8316 24175 8318 24195
rect 8412 24175 8414 24195
rect 8700 24175 8702 24195
rect 8748 24175 8750 24195
rect 8796 24175 8798 24195
rect 8844 24175 8846 24195
rect 8868 24175 8870 24195
rect 9516 24175 9518 24195
rect 9660 24175 9662 24195
rect 9684 24175 9686 24195
rect 9780 24175 9782 24195
rect 9804 24175 9806 24195
rect 9828 24175 9830 24195
rect 10044 24175 10046 24195
rect 10140 24175 10142 24195
rect 10236 24175 10238 24195
rect 10332 24175 10334 24195
rect 10380 24175 10382 24195
rect 10428 24175 10430 24195
rect 10524 24175 10526 24195
rect 10548 24175 10550 24195
rect 10620 24175 10622 24195
rect 10644 24175 10646 24195
rect 10716 24175 10718 24195
rect 10825 24175 10859 24176
rect 10860 24175 10862 24195
rect 10956 24175 10958 24195
rect 11052 24175 11054 24195
rect 11100 24175 11102 24195
rect 11172 24175 11174 24195
rect 11220 24175 11222 24195
rect 11340 24175 11342 24195
rect 11436 24175 11438 24195
rect 11676 24175 11678 24195
rect 11724 24175 11726 24195
rect 11772 24175 11774 24195
rect 11796 24175 11798 24195
rect 12060 24175 12062 24195
rect 12276 24175 12278 24195
rect 12324 24175 12326 24195
rect 12372 24175 12374 24195
rect 12420 24175 12422 24195
rect 12468 24175 12470 24195
rect 12564 24175 12566 24195
rect 12780 24175 12782 24195
rect 12876 24175 12878 24195
rect 12972 24175 12974 24195
rect 13044 24175 13046 24195
rect 13068 24175 13070 24195
rect 13164 24175 13166 24195
rect 13332 24175 13334 24195
rect 13500 24175 13502 24195
rect 13572 24175 13574 24195
rect 13668 24175 13670 24195
rect 13716 24175 13718 24195
rect 13836 24175 13838 24195
rect 13921 24190 13924 24195
rect 13931 24176 13934 24190
rect 13932 24175 13934 24176
rect 14004 24175 14006 24195
rect 14028 24175 14031 24192
rect 14100 24175 14102 24195
rect 14940 24175 14942 24195
rect 15036 24175 15038 24195
rect 15276 24175 15278 24195
rect 15372 24175 15374 24195
rect 15420 24175 15422 24195
rect 15468 24175 15470 24195
rect 15564 24175 15566 24195
rect 15660 24175 15662 24195
rect 15732 24175 15734 24195
rect 15756 24175 15758 24195
rect 15804 24175 15806 24195
rect 15828 24175 15830 24195
rect 15852 24175 15854 24195
rect 15948 24175 15950 24195
rect 15972 24175 15974 24195
rect 16044 24175 16046 24195
rect 16068 24175 16070 24195
rect 16164 24175 16166 24195
rect 16260 24175 16262 24195
rect 16284 24175 16286 24195
rect 16380 24175 16382 24195
rect 16476 24175 16478 24195
rect 16548 24175 16550 24195
rect 16572 24175 16574 24195
rect 16668 24175 16670 24195
rect 16692 24175 16694 24195
rect 16764 24175 16766 24195
rect 16788 24175 16790 24195
rect 16884 24175 16886 24195
rect 16908 24175 16910 24195
rect 17028 24175 17030 24195
rect 17124 24175 17126 24195
rect 17196 24175 17198 24195
rect 17220 24175 17222 24195
rect 17292 24175 17294 24195
rect 17316 24175 17318 24195
rect 17964 24175 17966 24195
rect 18060 24175 18062 24195
rect 18132 24175 18134 24195
rect 18228 24175 18230 24195
rect 18492 24175 18494 24195
rect 18540 24175 18542 24195
rect 18636 24175 18638 24195
rect 18732 24175 18734 24195
rect 18828 24175 18830 24195
rect 18924 24175 18926 24195
rect 18972 24175 18974 24195
rect 19020 24175 19022 24195
rect 19068 24175 19070 24195
rect 19140 24175 19142 24195
rect 19164 24175 19166 24195
rect 19236 24175 19238 24195
rect 19260 24175 19262 24195
rect 19788 24175 19790 24195
rect 19836 24175 19838 24195
rect 19860 24175 19862 24195
rect 19884 24175 19886 24195
rect 19956 24175 19958 24195
rect 19980 24175 19982 24195
rect 20004 24175 20006 24195
rect 20052 24175 20054 24195
rect 20076 24175 20078 24195
rect 20100 24175 20102 24195
rect 20172 24175 20174 24195
rect 20196 24175 20198 24195
rect 20292 24175 20294 24195
rect 20388 24175 20390 24195
rect 20412 24175 20414 24195
rect 20508 24175 20510 24195
rect 20532 24175 20534 24195
rect 20604 24175 20606 24195
rect 20628 24175 20630 24195
rect 20892 24175 20894 24195
rect 20964 24175 20966 24195
rect 20988 24175 20990 24195
rect 21108 24175 21110 24195
rect 21204 24175 21206 24195
rect 21300 24176 21302 24195
rect 21313 24190 21316 24195
rect 21324 24190 21326 24195
rect 21323 24176 21326 24190
rect 21289 24175 21323 24176
rect -6743 24171 14021 24175
rect -6743 24168 -6739 24171
rect -6732 24168 -6729 24171
rect -6647 24166 -6644 24171
rect -6636 24168 -6634 24171
rect -6540 24168 -6538 24171
rect -6636 24166 -6633 24168
rect -6647 24158 -6643 24166
rect -6657 24152 -6647 24158
rect -6637 24152 -6633 24166
rect -6540 24152 -6537 24168
rect -6551 24151 -6517 24152
rect -6444 24151 -6442 24171
rect -6348 24151 -6346 24171
rect -6252 24151 -6250 24171
rect -5892 24151 -5890 24171
rect -5340 24151 -5338 24171
rect -4716 24151 -4714 24171
rect -4500 24151 -4498 24171
rect -4284 24151 -4282 24171
rect -3876 24151 -3874 24171
rect -3828 24151 -3826 24171
rect -3540 24151 -3538 24171
rect -3468 24151 -3466 24171
rect -3324 24151 -3322 24171
rect -3108 24151 -3106 24171
rect -3012 24151 -3010 24171
rect -2988 24151 -2986 24171
rect -2916 24151 -2914 24171
rect -2868 24151 -2866 24171
rect -2772 24151 -2770 24171
rect -2364 24151 -2362 24171
rect -1908 24151 -1906 24171
rect -1452 24151 -1450 24171
rect -1356 24151 -1354 24171
rect -1260 24151 -1258 24171
rect -1236 24151 -1234 24171
rect -1140 24151 -1138 24171
rect -876 24151 -874 24171
rect -780 24151 -778 24171
rect -564 24151 -562 24171
rect -468 24151 -466 24171
rect -12 24151 -10 24171
rect 84 24151 86 24171
rect 348 24151 350 24171
rect 468 24151 470 24171
rect 492 24151 494 24171
rect 564 24151 566 24171
rect 588 24151 590 24171
rect 636 24151 638 24171
rect 660 24151 662 24171
rect 732 24151 734 24171
rect 948 24151 950 24171
rect 1044 24151 1046 24171
rect 1092 24151 1094 24171
rect 1140 24151 1142 24171
rect 1308 24151 1310 24171
rect 1356 24151 1358 24171
rect 1428 24151 1430 24171
rect 1572 24151 1574 24171
rect 1860 24151 1862 24171
rect 1956 24151 1958 24171
rect 2052 24151 2054 24171
rect 2148 24151 2150 24171
rect 2244 24151 2246 24171
rect 2460 24151 2462 24171
rect 2772 24151 2774 24171
rect 2868 24151 2870 24171
rect 2940 24151 2942 24171
rect 2988 24151 2990 24171
rect 3324 24151 3326 24171
rect 3540 24151 3542 24171
rect 3660 24151 3662 24171
rect 3780 24151 3782 24171
rect 4092 24151 4094 24171
rect 4188 24151 4190 24171
rect 4308 24151 4310 24171
rect 4404 24151 4406 24171
rect 4500 24151 4502 24171
rect 4596 24151 4598 24171
rect 4692 24151 4694 24171
rect 4932 24151 4934 24171
rect 4980 24151 4982 24171
rect 5028 24151 5030 24171
rect 5124 24151 5126 24171
rect 5220 24151 5222 24171
rect 5460 24151 5462 24171
rect 5508 24151 5510 24171
rect 5556 24151 5558 24171
rect 5652 24151 5654 24171
rect 5748 24151 5750 24171
rect 5796 24151 5798 24171
rect 5844 24151 5846 24171
rect 5892 24151 5894 24171
rect 6276 24151 6278 24171
rect 6300 24151 6302 24171
rect 6372 24151 6374 24171
rect 6396 24151 6398 24171
rect 6492 24151 6494 24171
rect 6516 24151 6518 24171
rect 6588 24151 6590 24171
rect 6612 24151 6614 24171
rect 6636 24151 6638 24171
rect 6684 24151 6686 24171
rect 6708 24151 6710 24171
rect 6804 24151 6806 24171
rect 6900 24151 6902 24171
rect 7164 24151 7166 24171
rect 7236 24151 7238 24171
rect 7284 24151 7286 24171
rect 7380 24151 7382 24171
rect 7404 24151 7406 24171
rect 7476 24151 7478 24171
rect 7500 24151 7502 24171
rect 7572 24151 7574 24171
rect 7596 24151 7598 24171
rect 7668 24151 7670 24171
rect 7692 24151 7694 24171
rect 7908 24151 7910 24171
rect 8124 24151 8126 24171
rect 8220 24151 8222 24171
rect 8316 24151 8318 24171
rect 8412 24151 8414 24171
rect 8700 24151 8702 24171
rect 8748 24151 8750 24171
rect 8796 24151 8798 24171
rect 8844 24151 8846 24171
rect 8868 24151 8870 24171
rect 9516 24151 9518 24171
rect 9660 24151 9662 24171
rect 9684 24151 9686 24171
rect 9780 24151 9782 24171
rect 9804 24151 9806 24171
rect 9828 24151 9830 24171
rect 10044 24151 10046 24171
rect 10140 24151 10142 24171
rect 10236 24151 10238 24171
rect 10332 24151 10334 24171
rect 10380 24151 10382 24171
rect 10428 24151 10430 24171
rect 10524 24151 10526 24171
rect 10548 24151 10550 24171
rect 10620 24151 10622 24171
rect 10644 24151 10646 24171
rect 10716 24151 10718 24171
rect 10860 24151 10862 24171
rect 10956 24151 10958 24171
rect 11052 24151 11054 24171
rect 11100 24151 11102 24171
rect 11172 24151 11174 24171
rect 11220 24151 11222 24171
rect 11340 24151 11342 24171
rect 11436 24151 11438 24171
rect 11676 24151 11678 24171
rect 11724 24151 11726 24171
rect 11772 24151 11774 24171
rect 11796 24151 11798 24171
rect 12060 24151 12062 24171
rect 12276 24151 12278 24171
rect 12324 24151 12326 24171
rect 12372 24151 12374 24171
rect 12420 24151 12422 24171
rect 12468 24151 12470 24171
rect 12564 24151 12566 24171
rect 12780 24151 12782 24171
rect 12876 24151 12878 24171
rect 12972 24151 12974 24171
rect 13044 24151 13046 24171
rect 13068 24151 13070 24171
rect 13164 24151 13166 24171
rect 13332 24151 13334 24171
rect 13500 24151 13502 24171
rect 13572 24151 13574 24171
rect 13668 24151 13670 24171
rect 13716 24152 13718 24171
rect 13705 24151 13739 24152
rect 13836 24151 13838 24171
rect 13932 24151 13934 24171
rect 14004 24151 14006 24171
rect 14007 24168 14021 24171
rect 14028 24171 21323 24175
rect 14028 24168 14045 24171
rect 14028 24151 14030 24168
rect 14100 24151 14102 24171
rect 14940 24151 14942 24171
rect 15036 24151 15038 24171
rect 15276 24151 15278 24171
rect 15372 24151 15374 24171
rect 15420 24151 15422 24171
rect 15468 24151 15470 24171
rect 15564 24151 15566 24171
rect 15660 24151 15662 24171
rect 15732 24151 15734 24171
rect 15756 24151 15758 24171
rect 15804 24151 15806 24171
rect 15828 24151 15830 24171
rect 15852 24151 15854 24171
rect 15948 24151 15950 24171
rect 15972 24151 15974 24171
rect 16044 24151 16046 24171
rect 16068 24151 16070 24171
rect 16164 24151 16166 24171
rect 16260 24151 16262 24171
rect 16284 24151 16286 24171
rect 16380 24151 16382 24171
rect 16476 24151 16478 24171
rect 16489 24151 16547 24152
rect 16548 24151 16550 24171
rect 16572 24151 16574 24171
rect 16668 24151 16670 24171
rect 16692 24151 16694 24171
rect 16764 24151 16766 24171
rect 16788 24151 16790 24171
rect 16884 24151 16886 24171
rect 16908 24151 16910 24171
rect 17028 24151 17030 24171
rect 17124 24151 17126 24171
rect 17196 24151 17198 24171
rect 17220 24151 17222 24171
rect 17292 24151 17294 24171
rect 17316 24151 17318 24171
rect 17964 24151 17966 24171
rect 18060 24151 18062 24171
rect 18132 24151 18134 24171
rect 18228 24151 18230 24171
rect 18492 24151 18494 24171
rect 18540 24151 18542 24171
rect 18636 24151 18638 24171
rect 18732 24151 18734 24171
rect 18828 24151 18830 24171
rect 18924 24151 18926 24171
rect 18972 24151 18974 24171
rect 19020 24151 19022 24171
rect 19068 24151 19070 24171
rect 19140 24151 19142 24171
rect 19164 24151 19166 24171
rect 19236 24151 19238 24171
rect 19260 24151 19262 24171
rect 19788 24151 19790 24171
rect 19836 24151 19838 24171
rect 19860 24151 19862 24171
rect 19884 24151 19886 24171
rect 19956 24151 19958 24171
rect 19980 24151 19982 24171
rect 20004 24151 20006 24171
rect 20052 24151 20054 24171
rect 20076 24151 20078 24171
rect 20100 24151 20102 24171
rect 20172 24151 20174 24171
rect 20196 24151 20198 24171
rect 20292 24151 20294 24171
rect 20388 24151 20390 24171
rect 20412 24151 20414 24171
rect 20508 24151 20510 24171
rect 20532 24151 20534 24171
rect 20604 24151 20606 24171
rect 20628 24151 20630 24171
rect 20892 24151 20894 24171
rect 20964 24151 20966 24171
rect 20988 24151 20990 24171
rect 21108 24151 21110 24171
rect 21204 24151 21206 24171
rect 21289 24166 21292 24171
rect 21300 24166 21302 24171
rect 21299 24152 21302 24166
rect 21217 24151 21251 24152
rect -6551 24147 21251 24151
rect -6551 24144 -6547 24147
rect -6540 24144 -6537 24147
rect -6444 24144 -6442 24147
rect -6444 24128 -6441 24144
rect -6348 24128 -6346 24147
rect -6455 24127 -6421 24128
rect -6407 24127 -6373 24128
rect -6455 24123 -6373 24127
rect -6359 24127 -6325 24128
rect -6252 24127 -6250 24147
rect -5892 24127 -5890 24147
rect -5529 24144 -5515 24147
rect -5340 24127 -5338 24147
rect -4716 24127 -4714 24147
rect -4500 24127 -4498 24147
rect -4284 24127 -4282 24147
rect -3876 24127 -3874 24147
rect -3828 24127 -3826 24147
rect -3540 24127 -3538 24147
rect -3468 24127 -3466 24147
rect -3324 24127 -3322 24147
rect -3108 24127 -3106 24147
rect -3012 24127 -3010 24147
rect -2988 24127 -2986 24147
rect -2916 24127 -2914 24147
rect -2868 24127 -2866 24147
rect -2772 24127 -2770 24147
rect -2364 24127 -2362 24147
rect -1908 24127 -1906 24147
rect -1487 24127 -1453 24128
rect -1452 24127 -1450 24147
rect -1356 24127 -1354 24147
rect -1260 24127 -1258 24147
rect -1236 24127 -1234 24147
rect -1140 24127 -1138 24147
rect -876 24127 -874 24147
rect -780 24127 -778 24147
rect -564 24127 -562 24147
rect -468 24127 -466 24147
rect -12 24127 -10 24147
rect 84 24127 86 24147
rect 348 24127 350 24147
rect 468 24127 470 24147
rect 492 24127 494 24147
rect 564 24127 566 24147
rect 588 24127 590 24147
rect 636 24127 638 24147
rect 660 24127 662 24147
rect 732 24127 734 24147
rect 948 24127 950 24147
rect 1044 24127 1046 24147
rect 1092 24127 1094 24147
rect 1140 24127 1142 24147
rect 1308 24127 1310 24147
rect 1356 24127 1358 24147
rect 1428 24127 1430 24147
rect 1572 24127 1574 24147
rect 1860 24127 1862 24147
rect 1956 24127 1958 24147
rect 2052 24127 2054 24147
rect 2148 24127 2150 24147
rect 2244 24127 2246 24147
rect 2460 24127 2462 24147
rect 2772 24127 2774 24147
rect 2868 24127 2870 24147
rect 2940 24127 2942 24147
rect 2988 24127 2990 24147
rect 3324 24127 3326 24147
rect 3540 24127 3542 24147
rect 3660 24127 3662 24147
rect 3780 24127 3782 24147
rect 4092 24127 4094 24147
rect 4188 24127 4190 24147
rect 4308 24127 4310 24147
rect 4404 24127 4406 24147
rect 4500 24127 4502 24147
rect 4596 24127 4598 24147
rect 4692 24127 4694 24147
rect 4932 24127 4934 24147
rect 4980 24127 4982 24147
rect 5028 24127 5030 24147
rect 5124 24127 5126 24147
rect 5220 24127 5222 24147
rect 5460 24127 5462 24147
rect 5508 24127 5510 24147
rect 5556 24127 5558 24147
rect 5652 24127 5654 24147
rect 5748 24127 5750 24147
rect 5796 24127 5798 24147
rect 5844 24127 5846 24147
rect 5892 24127 5894 24147
rect 6276 24127 6278 24147
rect 6300 24127 6302 24147
rect 6372 24127 6374 24147
rect 6396 24127 6398 24147
rect 6492 24127 6494 24147
rect 6516 24127 6518 24147
rect 6588 24127 6590 24147
rect 6612 24127 6614 24147
rect 6636 24127 6638 24147
rect 6684 24127 6686 24147
rect 6708 24127 6710 24147
rect 6804 24127 6806 24147
rect 6900 24127 6902 24147
rect 7129 24127 7163 24128
rect 7164 24127 7166 24147
rect 7236 24127 7238 24147
rect 7284 24127 7286 24147
rect 7380 24127 7382 24147
rect 7404 24127 7406 24147
rect 7476 24127 7478 24147
rect 7500 24127 7502 24147
rect 7572 24127 7574 24147
rect 7596 24127 7598 24147
rect 7668 24127 7670 24147
rect 7692 24127 7694 24147
rect 7908 24127 7910 24147
rect 8124 24127 8126 24147
rect 8220 24127 8222 24147
rect 8316 24127 8318 24147
rect 8412 24127 8414 24147
rect 8700 24127 8702 24147
rect 8748 24127 8750 24147
rect 8796 24127 8798 24147
rect 8844 24127 8846 24147
rect 8868 24127 8870 24147
rect 9516 24127 9518 24147
rect 9660 24127 9662 24147
rect 9684 24127 9686 24147
rect 9780 24127 9782 24147
rect 9804 24127 9806 24147
rect 9828 24127 9830 24147
rect 10044 24127 10046 24147
rect 10140 24127 10142 24147
rect 10236 24127 10238 24147
rect 10332 24127 10334 24147
rect 10380 24127 10382 24147
rect 10428 24127 10430 24147
rect 10524 24127 10526 24147
rect 10548 24127 10550 24147
rect 10620 24127 10622 24147
rect 10644 24127 10646 24147
rect 10716 24127 10718 24147
rect 10860 24127 10862 24147
rect 10911 24144 10925 24147
rect 10956 24127 10958 24147
rect 11052 24127 11054 24147
rect 11100 24127 11102 24147
rect 11172 24127 11174 24147
rect 11220 24127 11222 24147
rect 11340 24127 11342 24147
rect 11436 24127 11438 24147
rect 11676 24127 11678 24147
rect 11724 24127 11726 24147
rect 11772 24127 11774 24147
rect 11796 24127 11798 24147
rect 12060 24127 12062 24147
rect 12276 24127 12278 24147
rect 12324 24128 12326 24147
rect 12313 24127 12347 24128
rect 12372 24127 12374 24147
rect 12420 24127 12422 24147
rect 12468 24127 12470 24147
rect 12564 24127 12566 24147
rect 12780 24127 12782 24147
rect 12876 24127 12878 24147
rect 12972 24127 12974 24147
rect 13044 24127 13046 24147
rect 13068 24127 13070 24147
rect 13164 24127 13166 24147
rect 13332 24127 13334 24147
rect 13500 24127 13502 24147
rect 13572 24127 13574 24147
rect 13668 24128 13670 24147
rect 13705 24142 13708 24147
rect 13716 24142 13718 24147
rect 13715 24128 13718 24142
rect 13657 24127 13691 24128
rect 13836 24127 13838 24147
rect 13932 24127 13934 24147
rect 14004 24127 14006 24147
rect 14028 24127 14030 24147
rect 14100 24127 14102 24147
rect 14940 24127 14942 24147
rect 15001 24127 15035 24128
rect 15036 24127 15038 24147
rect 15276 24127 15278 24147
rect 15372 24127 15374 24147
rect 15420 24127 15422 24147
rect 15468 24127 15470 24147
rect 15564 24127 15566 24147
rect 15660 24127 15662 24147
rect 15732 24127 15734 24147
rect 15756 24127 15758 24147
rect 15804 24127 15806 24147
rect 15828 24127 15830 24147
rect 15852 24127 15854 24147
rect 15948 24127 15950 24147
rect 15972 24127 15974 24147
rect 16044 24127 16046 24147
rect 16068 24127 16070 24147
rect 16164 24127 16166 24147
rect 16260 24127 16262 24147
rect 16284 24127 16286 24147
rect 16380 24127 16382 24147
rect 16476 24127 16478 24147
rect 16548 24127 16550 24147
rect 16572 24127 16574 24147
rect 16596 24127 16599 24144
rect 16668 24127 16670 24147
rect 16692 24127 16694 24147
rect 16764 24127 16766 24147
rect 16788 24127 16790 24147
rect 16884 24127 16886 24147
rect 16908 24127 16910 24147
rect 17028 24127 17030 24147
rect 17124 24127 17126 24147
rect 17196 24127 17198 24147
rect 17220 24127 17222 24147
rect 17292 24127 17294 24147
rect 17316 24127 17318 24147
rect 17964 24127 17966 24147
rect 18060 24127 18062 24147
rect 18132 24127 18134 24147
rect 18228 24127 18230 24147
rect 18492 24127 18494 24147
rect 18540 24127 18542 24147
rect 18636 24127 18638 24147
rect 18732 24127 18734 24147
rect 18828 24127 18830 24147
rect 18924 24127 18926 24147
rect 18972 24127 18974 24147
rect 19020 24127 19022 24147
rect 19068 24127 19070 24147
rect 19140 24127 19142 24147
rect 19164 24127 19166 24147
rect 19236 24127 19238 24147
rect 19260 24127 19262 24147
rect 19788 24127 19790 24147
rect 19836 24127 19838 24147
rect 19860 24127 19862 24147
rect 19884 24127 19886 24147
rect 19956 24128 19958 24147
rect 19945 24127 19979 24128
rect 19980 24127 19982 24147
rect 20004 24127 20006 24147
rect 20052 24127 20054 24147
rect 20076 24127 20078 24147
rect 20100 24127 20102 24147
rect 20172 24127 20174 24147
rect 20196 24127 20198 24147
rect 20292 24127 20294 24147
rect 20388 24127 20390 24147
rect 20412 24127 20414 24147
rect 20508 24127 20510 24147
rect 20532 24127 20534 24147
rect 20604 24127 20606 24147
rect 20628 24127 20630 24147
rect 20892 24127 20894 24147
rect 20964 24127 20966 24147
rect 20988 24127 20990 24147
rect 21108 24127 21110 24147
rect 21204 24128 21206 24147
rect 21193 24127 21227 24128
rect -6359 24123 16589 24127
rect -6455 24120 -6451 24123
rect -6444 24120 -6441 24123
rect -6359 24118 -6356 24123
rect -6348 24120 -6346 24123
rect -6252 24120 -6250 24123
rect -6348 24118 -6345 24120
rect -6349 24104 -6345 24118
rect -6252 24104 -6249 24120
rect -6263 24103 -6229 24104
rect -5892 24103 -5890 24123
rect -5735 24103 -5701 24104
rect -6263 24099 -5701 24103
rect -5687 24103 -5653 24104
rect -5340 24103 -5338 24123
rect -4716 24103 -4714 24123
rect -4500 24103 -4498 24123
rect -4284 24103 -4282 24123
rect -3876 24103 -3874 24123
rect -3828 24103 -3826 24123
rect -3540 24103 -3538 24123
rect -3468 24103 -3466 24123
rect -3324 24103 -3322 24123
rect -3108 24103 -3106 24123
rect -3012 24103 -3010 24123
rect -2988 24103 -2986 24123
rect -2916 24103 -2914 24123
rect -2868 24103 -2866 24123
rect -2772 24103 -2770 24123
rect -2364 24103 -2362 24123
rect -1908 24103 -1906 24123
rect -1452 24103 -1450 24123
rect -1356 24103 -1354 24123
rect -1260 24103 -1258 24123
rect -1236 24103 -1234 24123
rect -1140 24103 -1138 24123
rect -876 24103 -874 24123
rect -780 24103 -778 24123
rect -564 24103 -562 24123
rect -468 24103 -466 24123
rect -12 24103 -10 24123
rect 84 24103 86 24123
rect 348 24103 350 24123
rect 468 24103 470 24123
rect 492 24103 494 24123
rect 564 24103 566 24123
rect 588 24103 590 24123
rect 636 24104 638 24123
rect 601 24103 659 24104
rect 660 24103 662 24123
rect 732 24103 734 24123
rect 948 24103 950 24123
rect 1044 24103 1046 24123
rect 1092 24103 1094 24123
rect 1140 24103 1142 24123
rect 1308 24103 1310 24123
rect 1356 24103 1358 24123
rect 1428 24103 1430 24123
rect 1572 24103 1574 24123
rect 1860 24103 1862 24123
rect 1956 24103 1958 24123
rect 2052 24103 2054 24123
rect 2148 24103 2150 24123
rect 2244 24103 2246 24123
rect 2460 24104 2462 24123
rect 2329 24103 2387 24104
rect 2425 24103 2483 24104
rect 2772 24103 2774 24123
rect 2868 24103 2870 24123
rect 2940 24103 2942 24123
rect 2988 24103 2990 24123
rect 3324 24103 3326 24123
rect 3540 24103 3542 24123
rect 3660 24103 3662 24123
rect 3780 24103 3782 24123
rect 4092 24103 4094 24123
rect 4188 24103 4190 24123
rect 4308 24103 4310 24123
rect 4404 24103 4406 24123
rect 4500 24103 4502 24123
rect 4596 24103 4598 24123
rect 4692 24103 4694 24123
rect 4932 24103 4934 24123
rect 4980 24103 4982 24123
rect 5028 24103 5030 24123
rect 5124 24103 5126 24123
rect 5220 24103 5222 24123
rect 5460 24103 5462 24123
rect 5508 24103 5510 24123
rect 5556 24103 5558 24123
rect 5652 24103 5654 24123
rect 5748 24103 5750 24123
rect 5796 24103 5798 24123
rect 5844 24103 5846 24123
rect 5892 24103 5894 24123
rect 6276 24103 6278 24123
rect 6300 24103 6302 24123
rect 6372 24103 6374 24123
rect 6396 24103 6398 24123
rect 6492 24103 6494 24123
rect 6516 24103 6518 24123
rect 6588 24103 6590 24123
rect 6612 24103 6614 24123
rect 6636 24103 6638 24123
rect 6684 24103 6686 24123
rect 6708 24103 6710 24123
rect 6804 24103 6806 24123
rect 6900 24103 6902 24123
rect 7164 24103 7166 24123
rect 7236 24120 7238 24123
rect 7236 24103 7239 24120
rect 7284 24103 7286 24123
rect 7380 24103 7382 24123
rect 7404 24103 7406 24123
rect 7476 24103 7478 24123
rect 7500 24103 7502 24123
rect 7572 24103 7574 24123
rect 7596 24103 7598 24123
rect 7668 24103 7670 24123
rect 7692 24103 7694 24123
rect 7908 24103 7910 24123
rect 8124 24103 8126 24123
rect 8220 24103 8222 24123
rect 8316 24103 8318 24123
rect 8412 24103 8414 24123
rect 8700 24103 8702 24123
rect 8748 24103 8750 24123
rect 8796 24103 8798 24123
rect 8844 24103 8846 24123
rect 8868 24103 8870 24123
rect 9516 24103 9518 24123
rect 9660 24103 9662 24123
rect 9684 24103 9686 24123
rect 9780 24103 9782 24123
rect 9804 24103 9806 24123
rect 9828 24103 9830 24123
rect 10044 24103 10046 24123
rect 10140 24103 10142 24123
rect 10236 24103 10238 24123
rect 10332 24103 10334 24123
rect 10380 24103 10382 24123
rect 10428 24103 10430 24123
rect 10524 24103 10526 24123
rect 10548 24103 10550 24123
rect 10620 24103 10622 24123
rect 10644 24103 10646 24123
rect 10716 24103 10718 24123
rect 10860 24103 10862 24123
rect 10956 24103 10958 24123
rect 11052 24103 11054 24123
rect 11100 24103 11102 24123
rect 11172 24103 11174 24123
rect 11220 24103 11222 24123
rect 11340 24103 11342 24123
rect 11436 24103 11438 24123
rect 11676 24103 11678 24123
rect 11724 24103 11726 24123
rect 11772 24103 11774 24123
rect 11796 24103 11798 24123
rect 12060 24103 12062 24123
rect 12276 24103 12278 24123
rect 12313 24118 12316 24123
rect 12324 24118 12326 24123
rect 12323 24104 12326 24118
rect 12372 24103 12374 24123
rect 12420 24120 12422 24123
rect 12420 24103 12423 24120
rect 12468 24103 12470 24123
rect 12564 24103 12566 24123
rect 12780 24103 12782 24123
rect 12876 24103 12878 24123
rect 12972 24103 12974 24123
rect 13044 24103 13046 24123
rect 13068 24103 13070 24123
rect 13164 24103 13166 24123
rect 13332 24103 13334 24123
rect 13500 24103 13502 24123
rect 13572 24103 13574 24123
rect 13657 24118 13660 24123
rect 13668 24118 13670 24123
rect 13791 24120 13805 24123
rect 13667 24104 13670 24118
rect 13836 24103 13838 24123
rect 13932 24103 13934 24123
rect 14004 24103 14006 24123
rect 14028 24103 14030 24123
rect 14100 24103 14102 24123
rect 14940 24103 14942 24123
rect 15036 24103 15038 24123
rect 15276 24103 15278 24123
rect 15372 24103 15374 24123
rect 15420 24103 15422 24123
rect 15468 24103 15470 24123
rect 15564 24103 15566 24123
rect 15660 24103 15662 24123
rect 15732 24103 15734 24123
rect 15756 24103 15758 24123
rect 15804 24103 15806 24123
rect 15828 24103 15830 24123
rect 15852 24103 15854 24123
rect 15948 24103 15950 24123
rect 15972 24103 15974 24123
rect 16044 24103 16046 24123
rect 16068 24103 16070 24123
rect 16164 24103 16166 24123
rect 16260 24103 16262 24123
rect 16284 24103 16286 24123
rect 16380 24103 16382 24123
rect 16476 24103 16478 24123
rect 16548 24103 16550 24123
rect 16572 24103 16574 24123
rect 16575 24120 16589 24123
rect 16596 24123 21227 24127
rect 16596 24120 16613 24123
rect 16596 24103 16598 24120
rect 16668 24103 16670 24123
rect 16692 24103 16694 24123
rect 16764 24103 16766 24123
rect 16788 24103 16790 24123
rect 16884 24103 16886 24123
rect 16908 24103 16910 24123
rect 17028 24103 17030 24123
rect 17124 24103 17126 24123
rect 17196 24103 17198 24123
rect 17220 24103 17222 24123
rect 17292 24103 17294 24123
rect 17316 24103 17318 24123
rect 17964 24103 17966 24123
rect 18060 24103 18062 24123
rect 18132 24103 18134 24123
rect 18228 24103 18230 24123
rect 18492 24103 18494 24123
rect 18540 24103 18542 24123
rect 18636 24103 18638 24123
rect 18732 24103 18734 24123
rect 18828 24103 18830 24123
rect 18924 24103 18926 24123
rect 18972 24103 18974 24123
rect 19020 24103 19022 24123
rect 19068 24103 19070 24123
rect 19140 24103 19142 24123
rect 19164 24103 19166 24123
rect 19236 24103 19238 24123
rect 19260 24103 19262 24123
rect 19788 24103 19790 24123
rect 19836 24103 19838 24123
rect 19860 24103 19862 24123
rect 19884 24103 19886 24123
rect 19945 24118 19948 24123
rect 19956 24118 19958 24123
rect 19955 24104 19958 24118
rect 19980 24103 19982 24123
rect 20004 24103 20006 24123
rect 20052 24120 20054 24123
rect 20052 24103 20055 24120
rect 20076 24103 20078 24123
rect 20100 24103 20102 24123
rect 20172 24103 20174 24123
rect 20196 24103 20198 24123
rect 20292 24103 20294 24123
rect 20388 24103 20390 24123
rect 20412 24103 20414 24123
rect 20508 24103 20510 24123
rect 20532 24103 20534 24123
rect 20604 24103 20606 24123
rect 20628 24103 20630 24123
rect 20892 24103 20894 24123
rect 20964 24103 20966 24123
rect 20988 24103 20990 24123
rect 21108 24104 21110 24123
rect 21193 24118 21196 24123
rect 21204 24118 21206 24123
rect 21203 24104 21206 24118
rect 21001 24103 21059 24104
rect 21097 24103 21131 24104
rect -5687 24099 21131 24103
rect -6263 24096 -6259 24099
rect -6252 24096 -6249 24099
rect -6143 24079 -6109 24080
rect -5892 24079 -5890 24099
rect -5879 24079 -5845 24080
rect -6143 24075 -5845 24079
rect -5567 24079 -5533 24080
rect -5340 24079 -5338 24099
rect -4716 24079 -4714 24099
rect -4500 24079 -4498 24099
rect -4284 24079 -4282 24099
rect -3876 24079 -3874 24099
rect -3828 24079 -3826 24099
rect -3540 24079 -3538 24099
rect -3468 24079 -3466 24099
rect -3324 24079 -3322 24099
rect -3108 24079 -3106 24099
rect -3012 24079 -3010 24099
rect -2988 24079 -2986 24099
rect -2916 24079 -2914 24099
rect -2868 24079 -2866 24099
rect -2772 24079 -2770 24099
rect -2364 24079 -2362 24099
rect -1908 24079 -1906 24099
rect -1452 24079 -1450 24099
rect -1401 24096 -1387 24099
rect -1356 24079 -1354 24099
rect -1260 24079 -1258 24099
rect -1236 24079 -1234 24099
rect -1140 24079 -1138 24099
rect -876 24079 -874 24099
rect -780 24079 -778 24099
rect -564 24079 -562 24099
rect -468 24079 -466 24099
rect -12 24079 -10 24099
rect 84 24079 86 24099
rect 348 24079 350 24099
rect 468 24079 470 24099
rect 492 24079 494 24099
rect 564 24079 566 24099
rect 588 24079 590 24099
rect 625 24094 628 24099
rect 636 24094 638 24099
rect 635 24080 638 24094
rect 660 24079 662 24099
rect 732 24096 734 24099
rect 732 24079 735 24096
rect 948 24079 950 24099
rect 1044 24079 1046 24099
rect 1092 24079 1094 24099
rect 1140 24079 1142 24099
rect 1308 24079 1310 24099
rect 1356 24079 1358 24099
rect 1428 24079 1430 24099
rect 1572 24079 1574 24099
rect 1860 24079 1862 24099
rect 1956 24079 1958 24099
rect 2052 24079 2054 24099
rect 2148 24079 2150 24099
rect 2244 24079 2246 24099
rect 2329 24094 2332 24099
rect 2449 24094 2452 24099
rect 2460 24096 2462 24099
rect 2460 24094 2463 24096
rect 2339 24080 2342 24094
rect 2435 24086 2439 24094
rect 2449 24086 2453 24094
rect 2435 24080 2449 24086
rect 2459 24080 2463 24094
rect 2340 24079 2342 24080
rect 2436 24079 2439 24080
rect 2532 24079 2535 24096
rect 2617 24079 2675 24080
rect 2772 24079 2774 24099
rect 2868 24079 2870 24099
rect 2940 24079 2942 24099
rect 2988 24079 2990 24099
rect 3324 24079 3326 24099
rect 3540 24079 3542 24099
rect 3660 24079 3662 24099
rect 3780 24079 3782 24099
rect 4092 24079 4094 24099
rect 4188 24079 4190 24099
rect 4308 24079 4310 24099
rect 4404 24079 4406 24099
rect 4500 24079 4502 24099
rect 4596 24079 4598 24099
rect 4692 24079 4694 24099
rect 4932 24079 4934 24099
rect 4980 24079 4982 24099
rect 5028 24079 5030 24099
rect 5124 24079 5126 24099
rect 5220 24079 5222 24099
rect 5460 24079 5462 24099
rect 5508 24079 5510 24099
rect 5556 24079 5558 24099
rect 5652 24079 5654 24099
rect 5748 24079 5750 24099
rect 5796 24079 5798 24099
rect 5844 24079 5846 24099
rect 5892 24079 5894 24099
rect 6276 24079 6278 24099
rect 6300 24079 6302 24099
rect 6372 24079 6374 24099
rect 6396 24079 6398 24099
rect 6492 24079 6494 24099
rect 6516 24079 6518 24099
rect 6588 24079 6590 24099
rect 6612 24079 6614 24099
rect 6636 24079 6638 24099
rect 6684 24079 6686 24099
rect 6708 24079 6710 24099
rect 6804 24079 6806 24099
rect 6900 24079 6902 24099
rect 7164 24079 7166 24099
rect 7215 24096 7229 24099
rect 7236 24096 7239 24099
rect 7284 24079 7286 24099
rect 7380 24079 7382 24099
rect 7404 24079 7406 24099
rect 7476 24079 7478 24099
rect 7500 24079 7502 24099
rect 7572 24079 7574 24099
rect 7596 24079 7598 24099
rect 7668 24079 7670 24099
rect 7692 24079 7694 24099
rect 7908 24079 7910 24099
rect 8124 24079 8126 24099
rect 8220 24079 8222 24099
rect 8316 24079 8318 24099
rect 8412 24079 8414 24099
rect 8700 24079 8702 24099
rect 8748 24079 8750 24099
rect 8796 24079 8798 24099
rect 8844 24079 8846 24099
rect 8868 24079 8870 24099
rect 9516 24079 9518 24099
rect 9660 24079 9662 24099
rect 9684 24079 9686 24099
rect 9780 24079 9782 24099
rect 9804 24079 9806 24099
rect 9828 24079 9830 24099
rect 10044 24079 10046 24099
rect 10140 24079 10142 24099
rect 10236 24079 10238 24099
rect 10332 24079 10334 24099
rect 10380 24079 10382 24099
rect 10428 24079 10430 24099
rect 10524 24079 10526 24099
rect 10548 24079 10550 24099
rect 10620 24079 10622 24099
rect 10644 24079 10646 24099
rect 10716 24079 10718 24099
rect 10860 24079 10862 24099
rect 10956 24079 10958 24099
rect 11052 24079 11054 24099
rect 11100 24079 11102 24099
rect 11172 24079 11174 24099
rect 11220 24079 11222 24099
rect 11340 24079 11342 24099
rect 11436 24079 11438 24099
rect 11676 24079 11678 24099
rect 11724 24079 11726 24099
rect 11772 24079 11774 24099
rect 11796 24079 11798 24099
rect 12060 24079 12062 24099
rect 12276 24079 12278 24099
rect 12372 24079 12374 24099
rect 12399 24096 12413 24099
rect 12420 24096 12423 24099
rect 12468 24079 12470 24099
rect 12564 24079 12566 24099
rect 12780 24079 12782 24099
rect 12876 24079 12878 24099
rect 12972 24079 12974 24099
rect 13044 24079 13046 24099
rect 13068 24079 13070 24099
rect 13164 24079 13166 24099
rect 13332 24079 13334 24099
rect 13500 24079 13502 24099
rect 13572 24079 13574 24099
rect 13743 24096 13757 24099
rect 13836 24079 13838 24099
rect 13932 24079 13934 24099
rect 14004 24079 14006 24099
rect 14028 24079 14030 24099
rect 14100 24079 14102 24099
rect 14940 24079 14942 24099
rect 15036 24079 15038 24099
rect 15087 24096 15101 24099
rect 15276 24079 15278 24099
rect 15372 24079 15374 24099
rect 15420 24079 15422 24099
rect 15468 24079 15470 24099
rect 15564 24079 15566 24099
rect 15660 24079 15662 24099
rect 15732 24079 15734 24099
rect 15756 24079 15758 24099
rect 15804 24079 15806 24099
rect 15828 24079 15830 24099
rect 15852 24079 15854 24099
rect 15948 24079 15950 24099
rect 15972 24079 15974 24099
rect 16044 24079 16046 24099
rect 16068 24079 16070 24099
rect 16164 24079 16166 24099
rect 16260 24079 16262 24099
rect 16284 24079 16286 24099
rect 16380 24079 16382 24099
rect 16476 24079 16478 24099
rect 16548 24079 16550 24099
rect 16572 24079 16574 24099
rect 16596 24079 16598 24099
rect 16668 24079 16670 24099
rect 16692 24079 16694 24099
rect 16764 24079 16766 24099
rect 16788 24079 16790 24099
rect 16884 24079 16886 24099
rect 16908 24079 16910 24099
rect 17028 24079 17030 24099
rect 17124 24079 17126 24099
rect 17196 24079 17198 24099
rect 17220 24079 17222 24099
rect 17292 24079 17294 24099
rect 17316 24079 17318 24099
rect 17964 24079 17966 24099
rect 18060 24079 18062 24099
rect 18132 24079 18134 24099
rect 18228 24079 18230 24099
rect 18492 24079 18494 24099
rect 18540 24079 18542 24099
rect 18636 24079 18638 24099
rect 18732 24079 18734 24099
rect 18828 24079 18830 24099
rect 18924 24079 18926 24099
rect 18972 24079 18974 24099
rect 19020 24079 19022 24099
rect 19068 24079 19070 24099
rect 19140 24079 19142 24099
rect 19164 24079 19166 24099
rect 19236 24079 19238 24099
rect 19260 24079 19262 24099
rect 19788 24079 19790 24099
rect 19836 24079 19838 24099
rect 19860 24079 19862 24099
rect 19884 24079 19886 24099
rect 19980 24079 19982 24099
rect 20004 24079 20006 24099
rect 20031 24096 20045 24099
rect 20052 24096 20055 24099
rect 20076 24079 20078 24099
rect 20100 24079 20102 24099
rect 20172 24079 20174 24099
rect 20196 24079 20198 24099
rect 20292 24079 20294 24099
rect 20388 24079 20390 24099
rect 20412 24079 20414 24099
rect 20508 24079 20510 24099
rect 20532 24079 20534 24099
rect 20604 24079 20606 24099
rect 20628 24079 20630 24099
rect 20892 24079 20894 24099
rect 20964 24079 20966 24099
rect 20988 24080 20990 24099
rect 21097 24094 21100 24099
rect 21108 24096 21110 24099
rect 21108 24094 21111 24096
rect 21107 24086 21111 24094
rect 21121 24086 21125 24094
rect 21107 24080 21121 24086
rect 20977 24079 21011 24080
rect -5567 24075 701 24079
rect -5892 24056 -5890 24075
rect -5999 24055 -5965 24056
rect -5903 24055 -5869 24056
rect -5999 24051 -5869 24055
rect -5447 24055 -5413 24056
rect -5340 24055 -5338 24075
rect -5183 24055 -5149 24056
rect -5447 24051 -5149 24055
rect -5063 24055 -5029 24056
rect -4716 24055 -4714 24075
rect -4500 24055 -4498 24075
rect -4284 24055 -4282 24075
rect -3876 24055 -3874 24075
rect -3828 24055 -3826 24075
rect -3540 24055 -3538 24075
rect -3468 24055 -3466 24075
rect -3324 24055 -3322 24075
rect -3108 24055 -3106 24075
rect -3012 24055 -3010 24075
rect -2988 24055 -2986 24075
rect -2916 24055 -2914 24075
rect -2868 24055 -2866 24075
rect -2772 24055 -2770 24075
rect -2364 24055 -2362 24075
rect -1908 24055 -1906 24075
rect -1452 24055 -1450 24075
rect -1356 24055 -1354 24075
rect -1260 24055 -1258 24075
rect -1236 24055 -1234 24075
rect -1140 24055 -1138 24075
rect -876 24055 -874 24075
rect -780 24055 -778 24075
rect -564 24055 -562 24075
rect -468 24055 -466 24075
rect -12 24055 -10 24075
rect 84 24055 86 24075
rect 348 24055 350 24075
rect 468 24055 470 24075
rect 492 24055 494 24075
rect 564 24055 566 24075
rect 588 24055 590 24075
rect 660 24055 662 24075
rect 687 24072 701 24075
rect 711 24075 2429 24079
rect 711 24072 725 24075
rect 732 24072 735 24075
rect 948 24055 950 24075
rect 1044 24055 1046 24075
rect 1092 24055 1094 24075
rect 1140 24055 1142 24075
rect 1308 24055 1310 24075
rect 1356 24055 1358 24075
rect 1428 24055 1430 24075
rect 1572 24055 1574 24075
rect 1860 24055 1862 24075
rect 1956 24055 1958 24075
rect 2052 24055 2054 24075
rect 2148 24055 2150 24075
rect 2244 24055 2246 24075
rect 2340 24055 2342 24075
rect 2415 24072 2429 24075
rect 2436 24075 2525 24079
rect 2436 24072 2453 24075
rect 2511 24072 2525 24075
rect 2532 24075 21011 24079
rect 2532 24072 2549 24075
rect 2436 24055 2438 24072
rect 2473 24055 2507 24056
rect 2532 24055 2534 24072
rect 2617 24070 2620 24075
rect 2627 24056 2630 24070
rect 2628 24055 2630 24056
rect 2724 24055 2727 24072
rect 2772 24056 2774 24075
rect 2761 24055 2795 24056
rect 2868 24055 2870 24075
rect 2940 24055 2942 24075
rect 2988 24055 2990 24075
rect 3324 24055 3326 24075
rect 3540 24055 3542 24075
rect 3660 24056 3662 24075
rect 3649 24055 3683 24056
rect 3780 24055 3782 24075
rect 4092 24055 4094 24075
rect 4188 24055 4190 24075
rect 4308 24055 4310 24075
rect 4404 24055 4406 24075
rect 4500 24055 4502 24075
rect 4596 24055 4598 24075
rect 4692 24055 4694 24075
rect 4932 24055 4934 24075
rect 4980 24055 4982 24075
rect 5028 24055 5030 24075
rect 5124 24055 5126 24075
rect 5220 24055 5222 24075
rect 5460 24055 5462 24075
rect 5508 24055 5510 24075
rect 5556 24055 5558 24075
rect 5652 24055 5654 24075
rect 5748 24055 5750 24075
rect 5796 24055 5798 24075
rect 5844 24055 5846 24075
rect 5892 24055 5894 24075
rect 6276 24055 6278 24075
rect 6300 24055 6302 24075
rect 6372 24055 6374 24075
rect 6396 24055 6398 24075
rect 6492 24055 6494 24075
rect 6516 24055 6518 24075
rect 6588 24055 6590 24075
rect 6612 24055 6614 24075
rect 6636 24055 6638 24075
rect 6684 24056 6686 24075
rect 6673 24055 6707 24056
rect 6708 24055 6710 24075
rect 6804 24055 6806 24075
rect 6900 24055 6902 24075
rect 7164 24055 7166 24075
rect 7284 24055 7286 24075
rect 7380 24055 7382 24075
rect 7404 24055 7406 24075
rect 7476 24055 7478 24075
rect 7500 24055 7502 24075
rect 7572 24055 7574 24075
rect 7596 24055 7598 24075
rect 7668 24055 7670 24075
rect 7692 24055 7694 24075
rect 7908 24055 7910 24075
rect 8124 24055 8126 24075
rect 8220 24055 8222 24075
rect 8316 24055 8318 24075
rect 8412 24055 8414 24075
rect 8700 24055 8702 24075
rect 8748 24055 8750 24075
rect 8796 24055 8798 24075
rect 8844 24055 8846 24075
rect 8868 24055 8870 24075
rect 9516 24055 9518 24075
rect 9660 24055 9662 24075
rect 9684 24055 9686 24075
rect 9780 24055 9782 24075
rect 9804 24055 9806 24075
rect 9828 24055 9830 24075
rect 10044 24055 10046 24075
rect 10140 24055 10142 24075
rect 10236 24055 10238 24075
rect 10332 24055 10334 24075
rect 10380 24055 10382 24075
rect 10428 24055 10430 24075
rect 10524 24055 10526 24075
rect 10548 24055 10550 24075
rect 10620 24055 10622 24075
rect 10644 24055 10646 24075
rect 10716 24055 10718 24075
rect 10860 24055 10862 24075
rect 10956 24055 10958 24075
rect 11052 24055 11054 24075
rect 11100 24055 11102 24075
rect 11172 24055 11174 24075
rect 11220 24055 11222 24075
rect 11340 24055 11342 24075
rect 11436 24055 11438 24075
rect 11676 24055 11678 24075
rect 11724 24055 11726 24075
rect 11772 24055 11774 24075
rect 11796 24055 11798 24075
rect 12060 24055 12062 24075
rect 12276 24055 12278 24075
rect 12372 24055 12374 24075
rect 12468 24055 12470 24075
rect 12564 24055 12566 24075
rect 12780 24055 12782 24075
rect 12876 24055 12878 24075
rect 12972 24055 12974 24075
rect 13044 24055 13046 24075
rect 13068 24055 13070 24075
rect 13164 24055 13166 24075
rect 13332 24055 13334 24075
rect 13500 24055 13502 24075
rect 13572 24055 13574 24075
rect 13836 24055 13838 24075
rect 13932 24055 13934 24075
rect 14004 24055 14006 24075
rect 14028 24055 14030 24075
rect 14100 24055 14102 24075
rect 14940 24055 14942 24075
rect 15036 24055 15038 24075
rect 15276 24055 15278 24075
rect 15372 24055 15374 24075
rect 15420 24055 15422 24075
rect 15468 24055 15470 24075
rect 15564 24055 15566 24075
rect 15660 24055 15662 24075
rect 15732 24055 15734 24075
rect 15756 24055 15758 24075
rect 15804 24055 15806 24075
rect 15828 24055 15830 24075
rect 15852 24055 15854 24075
rect 15948 24055 15950 24075
rect 15972 24055 15974 24075
rect 16044 24055 16046 24075
rect 16068 24055 16070 24075
rect 16164 24055 16166 24075
rect 16260 24055 16262 24075
rect 16284 24055 16286 24075
rect 16380 24055 16382 24075
rect 16476 24055 16478 24075
rect 16548 24055 16550 24075
rect 16572 24055 16574 24075
rect 16596 24055 16598 24075
rect 16668 24055 16670 24075
rect 16692 24055 16694 24075
rect 16764 24055 16766 24075
rect 16788 24055 16790 24075
rect 16884 24055 16886 24075
rect 16908 24055 16910 24075
rect 17028 24055 17030 24075
rect 17124 24055 17126 24075
rect 17196 24055 17198 24075
rect 17220 24055 17222 24075
rect 17292 24055 17294 24075
rect 17316 24055 17318 24075
rect 17964 24055 17966 24075
rect 18060 24055 18062 24075
rect 18132 24055 18134 24075
rect 18228 24055 18230 24075
rect 18492 24055 18494 24075
rect 18540 24055 18542 24075
rect 18636 24055 18638 24075
rect 18732 24055 18734 24075
rect 18828 24055 18830 24075
rect 18924 24055 18926 24075
rect 18972 24055 18974 24075
rect 19020 24055 19022 24075
rect 19068 24055 19070 24075
rect 19140 24055 19142 24075
rect 19164 24055 19166 24075
rect 19236 24055 19238 24075
rect 19260 24055 19262 24075
rect 19788 24055 19790 24075
rect 19836 24055 19838 24075
rect 19860 24055 19862 24075
rect 19884 24055 19886 24075
rect 19980 24055 19982 24075
rect 20004 24055 20006 24075
rect 20076 24055 20078 24075
rect 20100 24055 20102 24075
rect 20172 24055 20174 24075
rect 20196 24055 20198 24075
rect 20292 24055 20294 24075
rect 20388 24055 20390 24075
rect 20412 24055 20414 24075
rect 20508 24055 20510 24075
rect 20532 24055 20534 24075
rect 20604 24055 20606 24075
rect 20628 24056 20630 24075
rect 20892 24056 20894 24075
rect 20964 24056 20966 24075
rect 20977 24070 20980 24075
rect 20988 24070 20990 24075
rect 20987 24056 20990 24070
rect 20617 24055 20651 24056
rect -5063 24051 2717 24055
rect -5903 24046 -5900 24051
rect -5892 24048 -5890 24051
rect -5340 24048 -5338 24051
rect -5892 24046 -5889 24048
rect -5893 24032 -5889 24046
rect -5340 24032 -5337 24048
rect -5351 24031 -5317 24032
rect -5207 24031 -5173 24032
rect -5351 24027 -5173 24031
rect -4943 24031 -4909 24032
rect -4716 24031 -4714 24051
rect -4631 24031 -4573 24032
rect -4500 24031 -4498 24051
rect -4284 24031 -4282 24051
rect -3876 24031 -3874 24051
rect -3828 24031 -3826 24051
rect -3540 24031 -3538 24051
rect -3468 24031 -3466 24051
rect -3324 24031 -3322 24051
rect -3108 24031 -3106 24051
rect -3012 24031 -3010 24051
rect -2988 24031 -2986 24051
rect -2916 24031 -2914 24051
rect -2868 24031 -2866 24051
rect -2772 24031 -2770 24051
rect -2364 24031 -2362 24051
rect -1908 24031 -1906 24051
rect -1452 24031 -1450 24051
rect -1356 24031 -1354 24051
rect -1260 24031 -1258 24051
rect -1236 24031 -1234 24051
rect -1140 24031 -1138 24051
rect -876 24031 -874 24051
rect -780 24031 -778 24051
rect -564 24031 -562 24051
rect -468 24031 -466 24051
rect -12 24031 -10 24051
rect 84 24031 86 24051
rect 169 24031 227 24032
rect 348 24031 350 24051
rect 468 24031 470 24051
rect 492 24031 494 24051
rect 564 24031 566 24051
rect 588 24031 590 24051
rect 660 24031 662 24051
rect 948 24031 950 24051
rect 1044 24031 1046 24051
rect 1092 24031 1094 24051
rect 1140 24031 1142 24051
rect 1308 24031 1310 24051
rect 1356 24031 1358 24051
rect 1428 24031 1430 24051
rect 1572 24031 1574 24051
rect 1860 24031 1862 24051
rect 1956 24031 1958 24051
rect 2052 24031 2054 24051
rect 2148 24031 2150 24051
rect 2244 24031 2246 24051
rect 2340 24031 2342 24051
rect 2436 24031 2438 24051
rect 2532 24031 2534 24051
rect 2628 24031 2630 24051
rect 2703 24048 2717 24051
rect 2724 24051 20651 24055
rect 20785 24055 20819 24056
rect 20857 24055 20915 24056
rect 20953 24055 20987 24056
rect 20785 24051 20987 24055
rect 2724 24048 2741 24051
rect 2724 24031 2726 24048
rect 2761 24046 2764 24051
rect 2772 24046 2774 24051
rect 2771 24032 2774 24046
rect 2868 24048 2870 24051
rect 2868 24031 2871 24048
rect 2940 24031 2942 24051
rect 2988 24031 2990 24051
rect 3324 24031 3326 24051
rect 3540 24031 3542 24051
rect 3649 24046 3652 24051
rect 3660 24046 3662 24051
rect 3659 24032 3662 24046
rect 3780 24031 3782 24051
rect 3961 24031 4019 24032
rect 4092 24031 4094 24051
rect 4188 24031 4190 24051
rect 4308 24031 4310 24051
rect 4404 24031 4406 24051
rect 4500 24031 4502 24051
rect 4596 24031 4598 24051
rect 4692 24031 4694 24051
rect 4932 24031 4934 24051
rect 4980 24031 4982 24051
rect 5028 24031 5030 24051
rect 5124 24031 5126 24051
rect 5220 24031 5222 24051
rect 5460 24031 5462 24051
rect 5508 24031 5510 24051
rect 5556 24031 5558 24051
rect 5652 24031 5654 24051
rect 5748 24031 5750 24051
rect 5796 24031 5798 24051
rect 5844 24031 5846 24051
rect 5892 24031 5894 24051
rect 6276 24031 6278 24051
rect 6300 24031 6302 24051
rect 6372 24031 6374 24051
rect 6396 24031 6398 24051
rect 6492 24031 6494 24051
rect 6516 24031 6518 24051
rect 6588 24031 6590 24051
rect 6612 24031 6614 24051
rect 6636 24031 6638 24051
rect 6673 24046 6676 24051
rect 6684 24046 6686 24051
rect 6683 24032 6686 24046
rect 6708 24031 6710 24051
rect 6804 24031 6806 24051
rect 6900 24031 6902 24051
rect 7164 24031 7166 24051
rect 7284 24031 7286 24051
rect 7380 24031 7382 24051
rect 7404 24031 7406 24051
rect 7476 24031 7478 24051
rect 7500 24031 7502 24051
rect 7572 24031 7574 24051
rect 7596 24031 7598 24051
rect 7668 24031 7670 24051
rect 7692 24031 7694 24051
rect 7908 24031 7910 24051
rect 8124 24031 8126 24051
rect 8220 24031 8222 24051
rect 8316 24031 8318 24051
rect 8412 24031 8414 24051
rect 8700 24031 8702 24051
rect 8748 24031 8750 24051
rect 8796 24031 8798 24051
rect 8844 24031 8846 24051
rect 8868 24031 8870 24051
rect 9516 24031 9518 24051
rect 9660 24031 9662 24051
rect 9684 24031 9686 24051
rect 9780 24031 9782 24051
rect 9804 24031 9806 24051
rect 9828 24031 9830 24051
rect 10044 24031 10046 24051
rect 10140 24031 10142 24051
rect 10236 24031 10238 24051
rect 10332 24031 10334 24051
rect 10380 24031 10382 24051
rect 10428 24031 10430 24051
rect 10524 24031 10526 24051
rect 10548 24031 10550 24051
rect 10620 24031 10622 24051
rect 10644 24031 10646 24051
rect 10716 24031 10718 24051
rect 10860 24031 10862 24051
rect 10956 24031 10958 24051
rect 11052 24031 11054 24051
rect 11100 24031 11102 24051
rect 11172 24031 11174 24051
rect 11220 24031 11222 24051
rect 11340 24031 11342 24051
rect 11436 24031 11438 24051
rect 11676 24031 11678 24051
rect 11724 24031 11726 24051
rect 11772 24031 11774 24051
rect 11796 24031 11798 24051
rect 12060 24031 12062 24051
rect 12276 24031 12278 24051
rect 12372 24031 12374 24051
rect 12468 24031 12470 24051
rect 12564 24031 12566 24051
rect 12780 24031 12782 24051
rect 12876 24031 12878 24051
rect 12972 24031 12974 24051
rect 13044 24031 13046 24051
rect 13068 24031 13070 24051
rect 13164 24031 13166 24051
rect 13332 24031 13334 24051
rect 13500 24031 13502 24051
rect 13572 24031 13574 24051
rect 13836 24031 13838 24051
rect 13932 24031 13934 24051
rect 14004 24031 14006 24051
rect 14028 24031 14030 24051
rect 14100 24031 14102 24051
rect 14940 24031 14942 24051
rect 15036 24031 15038 24051
rect 15276 24031 15278 24051
rect 15372 24031 15374 24051
rect 15420 24031 15422 24051
rect 15468 24031 15470 24051
rect 15564 24031 15566 24051
rect 15660 24031 15662 24051
rect 15673 24031 15731 24032
rect 15732 24031 15734 24051
rect 15756 24031 15758 24051
rect 15804 24031 15806 24051
rect 15828 24031 15830 24051
rect 15852 24031 15854 24051
rect 15948 24031 15950 24051
rect 15972 24031 15974 24051
rect 16044 24031 16046 24051
rect 16068 24031 16070 24051
rect 16164 24031 16166 24051
rect 16260 24031 16262 24051
rect 16284 24031 16286 24051
rect 16380 24031 16382 24051
rect 16476 24031 16478 24051
rect 16548 24031 16550 24051
rect 16572 24031 16574 24051
rect 16596 24031 16598 24051
rect 16668 24031 16670 24051
rect 16692 24031 16694 24051
rect 16764 24031 16766 24051
rect 16788 24031 16790 24051
rect 16884 24031 16886 24051
rect 16908 24031 16910 24051
rect 17028 24031 17030 24051
rect 17124 24031 17126 24051
rect 17196 24031 17198 24051
rect 17220 24031 17222 24051
rect 17292 24031 17294 24051
rect 17316 24031 17318 24051
rect 17964 24031 17966 24051
rect 18060 24031 18062 24051
rect 18132 24031 18134 24051
rect 18228 24031 18230 24051
rect 18492 24031 18494 24051
rect 18540 24031 18542 24051
rect 18636 24031 18638 24051
rect 18732 24031 18734 24051
rect 18828 24031 18830 24051
rect 18924 24031 18926 24051
rect 18972 24031 18974 24051
rect 19020 24031 19022 24051
rect 19068 24031 19070 24051
rect 19140 24031 19142 24051
rect 19164 24031 19166 24051
rect 19236 24031 19238 24051
rect 19260 24031 19262 24051
rect 19788 24031 19790 24051
rect 19836 24031 19838 24051
rect 19860 24031 19862 24051
rect 19884 24031 19886 24051
rect 19980 24031 19982 24051
rect 20004 24031 20006 24051
rect 20076 24031 20078 24051
rect 20100 24031 20102 24051
rect 20172 24031 20174 24051
rect 20196 24031 20198 24051
rect 20292 24031 20294 24051
rect 20388 24031 20390 24051
rect 20412 24031 20414 24051
rect 20508 24031 20510 24051
rect 20532 24031 20534 24051
rect 20604 24032 20606 24051
rect 20617 24046 20620 24051
rect 20628 24046 20630 24051
rect 20627 24032 20630 24046
rect 20881 24046 20884 24051
rect 20892 24048 20894 24051
rect 20892 24046 20895 24048
rect 20953 24046 20956 24051
rect 20964 24048 20966 24051
rect 20964 24046 20967 24048
rect 20881 24038 20885 24046
rect 20871 24032 20881 24038
rect 20891 24032 20895 24046
rect 20963 24038 20967 24046
rect 20977 24038 20981 24046
rect 20963 24032 20977 24038
rect 20593 24031 20627 24032
rect -4943 24027 20627 24031
rect -5351 24024 -5347 24027
rect -5340 24024 -5337 24027
rect -4823 24007 -4789 24008
rect -4716 24007 -4714 24027
rect -4631 24022 -4628 24027
rect -4500 24024 -4498 24027
rect -4621 24008 -4618 24022
rect -4620 24007 -4618 24008
rect -4500 24007 -4497 24024
rect -4284 24007 -4282 24027
rect -3876 24007 -3874 24027
rect -3828 24007 -3826 24027
rect -3695 24007 -3661 24008
rect -3540 24007 -3538 24027
rect -3468 24007 -3466 24027
rect -3324 24007 -3322 24027
rect -3108 24007 -3106 24027
rect -3012 24007 -3010 24027
rect -2988 24007 -2986 24027
rect -2916 24007 -2914 24027
rect -2868 24007 -2866 24027
rect -2772 24007 -2770 24027
rect -2364 24007 -2362 24027
rect -1908 24007 -1906 24027
rect -1452 24007 -1450 24027
rect -1356 24007 -1354 24027
rect -1260 24007 -1258 24027
rect -1236 24007 -1234 24027
rect -1140 24007 -1138 24027
rect -876 24007 -874 24027
rect -780 24007 -778 24027
rect -564 24007 -562 24027
rect -468 24007 -466 24027
rect -12 24007 -10 24027
rect 84 24007 86 24027
rect 169 24022 172 24027
rect 179 24008 182 24022
rect 180 24007 182 24008
rect 348 24007 350 24027
rect 468 24007 470 24027
rect 492 24007 494 24027
rect 564 24007 566 24027
rect 588 24007 590 24027
rect 660 24007 662 24027
rect 948 24007 950 24027
rect 1044 24007 1046 24027
rect 1092 24007 1094 24027
rect 1140 24007 1142 24027
rect 1308 24007 1310 24027
rect 1356 24007 1358 24027
rect 1428 24008 1430 24027
rect 1417 24007 1451 24008
rect 1572 24007 1574 24027
rect 1860 24007 1862 24027
rect 1956 24007 1958 24027
rect 2052 24007 2054 24027
rect 2148 24007 2150 24027
rect 2244 24007 2246 24027
rect 2340 24007 2342 24027
rect 2436 24007 2438 24027
rect 2532 24007 2534 24027
rect 2559 24024 2573 24027
rect 2628 24007 2630 24027
rect 2724 24007 2726 24027
rect 2847 24024 2861 24027
rect 2868 24024 2871 24027
rect 2940 24007 2942 24027
rect 2988 24007 2990 24027
rect 3324 24007 3326 24027
rect 3540 24007 3542 24027
rect 3735 24024 3749 24027
rect 3780 24007 3782 24027
rect 4092 24024 4094 24027
rect 4092 24007 4095 24024
rect 4188 24007 4190 24027
rect 4308 24007 4310 24027
rect 4404 24008 4406 24027
rect 4393 24007 4427 24008
rect 4500 24007 4502 24027
rect 4596 24007 4598 24027
rect 4692 24007 4694 24027
rect 4932 24007 4934 24027
rect 4980 24007 4982 24027
rect 5028 24007 5030 24027
rect 5124 24007 5126 24027
rect 5220 24007 5222 24027
rect 5460 24007 5462 24027
rect 5508 24007 5510 24027
rect 5556 24007 5558 24027
rect 5652 24007 5654 24027
rect 5748 24007 5750 24027
rect 5796 24007 5798 24027
rect 5844 24007 5846 24027
rect 5892 24007 5894 24027
rect 6276 24007 6278 24027
rect 6300 24007 6302 24027
rect 6372 24007 6374 24027
rect 6396 24007 6398 24027
rect 6492 24007 6494 24027
rect 6516 24007 6518 24027
rect 6588 24007 6590 24027
rect 6612 24007 6614 24027
rect 6636 24007 6638 24027
rect 6708 24007 6710 24027
rect 6759 24024 6773 24027
rect 6804 24007 6806 24027
rect 6900 24007 6902 24027
rect 7164 24007 7166 24027
rect 7284 24007 7286 24027
rect 7380 24007 7382 24027
rect 7404 24007 7406 24027
rect 7476 24007 7478 24027
rect 7500 24007 7502 24027
rect 7572 24007 7574 24027
rect 7596 24007 7598 24027
rect 7668 24007 7670 24027
rect 7692 24007 7694 24027
rect 7908 24007 7910 24027
rect 8124 24007 8126 24027
rect 8220 24007 8222 24027
rect 8316 24007 8318 24027
rect 8412 24007 8414 24027
rect 8700 24007 8702 24027
rect 8748 24007 8750 24027
rect 8796 24007 8798 24027
rect 8844 24007 8846 24027
rect 8868 24007 8870 24027
rect 9001 24007 9035 24008
rect 9516 24007 9518 24027
rect 9660 24007 9662 24027
rect 9684 24007 9686 24027
rect 9780 24007 9782 24027
rect 9804 24007 9806 24027
rect 9828 24007 9830 24027
rect 10044 24007 10046 24027
rect 10140 24007 10142 24027
rect 10236 24007 10238 24027
rect 10332 24007 10334 24027
rect 10380 24007 10382 24027
rect 10428 24007 10430 24027
rect 10524 24007 10526 24027
rect 10548 24007 10550 24027
rect 10620 24007 10622 24027
rect 10644 24007 10646 24027
rect 10716 24007 10718 24027
rect 10860 24007 10862 24027
rect 10956 24007 10958 24027
rect 11052 24007 11054 24027
rect 11100 24007 11102 24027
rect 11172 24007 11174 24027
rect 11220 24007 11222 24027
rect 11340 24007 11342 24027
rect 11436 24007 11438 24027
rect 11676 24007 11678 24027
rect 11724 24007 11726 24027
rect 11772 24007 11774 24027
rect 11796 24007 11798 24027
rect 12060 24007 12062 24027
rect 12276 24007 12278 24027
rect 12372 24007 12374 24027
rect 12468 24007 12470 24027
rect 12564 24007 12566 24027
rect 12780 24007 12782 24027
rect 12876 24007 12878 24027
rect 12972 24007 12974 24027
rect 13044 24007 13046 24027
rect 13068 24007 13070 24027
rect 13164 24007 13166 24027
rect 13249 24007 13307 24008
rect 13332 24007 13334 24027
rect 13500 24007 13502 24027
rect 13572 24007 13574 24027
rect 13836 24007 13838 24027
rect 13932 24007 13934 24027
rect 14004 24007 14006 24027
rect 14028 24007 14030 24027
rect 14100 24007 14102 24027
rect 14940 24007 14942 24027
rect 15036 24007 15038 24027
rect 15276 24007 15278 24027
rect 15372 24007 15374 24027
rect 15420 24007 15422 24027
rect 15468 24007 15470 24027
rect 15564 24007 15566 24027
rect 15660 24007 15662 24027
rect 15673 24022 15676 24027
rect 15683 24008 15686 24022
rect 15684 24007 15686 24008
rect 15732 24007 15734 24027
rect 15756 24007 15758 24027
rect 15804 24024 15806 24027
rect 15804 24007 15807 24024
rect 15828 24007 15830 24027
rect 15852 24007 15854 24027
rect 15948 24007 15950 24027
rect 15972 24007 15974 24027
rect 16044 24007 16046 24027
rect 16068 24007 16070 24027
rect 16164 24007 16166 24027
rect 16260 24007 16262 24027
rect 16284 24007 16286 24027
rect 16380 24007 16382 24027
rect 16476 24007 16478 24027
rect 16548 24007 16550 24027
rect 16572 24007 16574 24027
rect 16596 24007 16598 24027
rect 16668 24007 16670 24027
rect 16692 24007 16694 24027
rect 16764 24007 16766 24027
rect 16788 24007 16790 24027
rect 16884 24007 16886 24027
rect 16908 24007 16910 24027
rect 17028 24007 17030 24027
rect 17124 24007 17126 24027
rect 17196 24007 17198 24027
rect 17220 24007 17222 24027
rect 17292 24007 17294 24027
rect 17316 24007 17318 24027
rect 17964 24007 17966 24027
rect 18060 24007 18062 24027
rect 18132 24007 18134 24027
rect 18228 24007 18230 24027
rect 18492 24007 18494 24027
rect 18540 24007 18542 24027
rect 18636 24007 18638 24027
rect 18732 24007 18734 24027
rect 18828 24007 18830 24027
rect 18924 24007 18926 24027
rect 18972 24007 18974 24027
rect 19020 24007 19022 24027
rect 19068 24007 19070 24027
rect 19140 24007 19142 24027
rect 19164 24007 19166 24027
rect 19236 24007 19238 24027
rect 19260 24007 19262 24027
rect 19788 24007 19790 24027
rect 19836 24007 19838 24027
rect 19860 24007 19862 24027
rect 19884 24007 19886 24027
rect 19980 24007 19982 24027
rect 20004 24007 20006 24027
rect 20076 24007 20078 24027
rect 20100 24007 20102 24027
rect 20172 24007 20174 24027
rect 20196 24007 20198 24027
rect 20292 24007 20294 24027
rect 20388 24007 20390 24027
rect 20412 24008 20414 24027
rect 20508 24008 20510 24027
rect 20532 24008 20534 24027
rect 20593 24022 20596 24027
rect 20604 24022 20606 24027
rect 20603 24008 20606 24022
rect 20401 24007 20459 24008
rect 20497 24007 20555 24008
rect 20569 24007 20603 24008
rect -4823 24003 -4531 24007
rect -4716 24000 -4714 24003
rect -4716 23984 -4713 24000
rect -4727 23983 -4693 23984
rect -4620 23983 -4618 24003
rect -4545 24000 -4531 24003
rect -4521 24003 269 24007
rect -4521 24000 -4507 24003
rect -4500 24000 -4497 24003
rect -4284 23983 -4282 24003
rect -3983 23983 -3949 23984
rect -3876 23983 -3874 24003
rect -3828 23983 -3826 24003
rect -3540 23983 -3538 24003
rect -3468 23983 -3466 24003
rect -3324 23983 -3322 24003
rect -3108 23983 -3106 24003
rect -3012 23983 -3010 24003
rect -2988 23983 -2986 24003
rect -2916 23983 -2914 24003
rect -2868 23983 -2866 24003
rect -2772 23983 -2770 24003
rect -2364 23983 -2362 24003
rect -1908 23983 -1906 24003
rect -1452 23983 -1450 24003
rect -1439 23983 -1381 23984
rect -1356 23983 -1354 24003
rect -1260 23983 -1258 24003
rect -1236 23983 -1234 24003
rect -1140 23983 -1138 24003
rect -876 23983 -874 24003
rect -780 23983 -778 24003
rect -564 23983 -562 24003
rect -468 23983 -466 24003
rect -12 23983 -10 24003
rect 84 23983 86 24003
rect 180 23983 182 24003
rect 255 24000 269 24003
rect 279 24003 4061 24007
rect 279 24000 293 24003
rect 348 23983 350 24003
rect 468 23983 470 24003
rect 492 23983 494 24003
rect 564 23983 566 24003
rect 588 23983 590 24003
rect 660 23983 662 24003
rect 948 23983 950 24003
rect 1044 23983 1046 24003
rect 1092 23983 1094 24003
rect 1140 23983 1142 24003
rect 1308 23983 1310 24003
rect 1356 23983 1358 24003
rect 1417 23998 1420 24003
rect 1428 23998 1430 24003
rect 1427 23984 1430 23998
rect 1572 23983 1574 24003
rect 1860 23983 1862 24003
rect 1956 23983 1958 24003
rect 2052 23983 2054 24003
rect 2148 23983 2150 24003
rect 2244 23983 2246 24003
rect 2340 23983 2342 24003
rect 2436 23983 2438 24003
rect 2532 23983 2534 24003
rect 2628 23983 2630 24003
rect 2724 23983 2726 24003
rect 2940 23983 2942 24003
rect 2988 23983 2990 24003
rect 3324 23983 3326 24003
rect 3540 23983 3542 24003
rect 3780 23983 3782 24003
rect 4047 24000 4061 24003
rect 4071 24003 15773 24007
rect 4071 24000 4085 24003
rect 4092 24000 4095 24003
rect 4188 23983 4190 24003
rect 4308 23983 4310 24003
rect 4393 23998 4396 24003
rect 4404 23998 4406 24003
rect 4403 23984 4406 23998
rect 4500 24000 4502 24003
rect 4500 23983 4503 24000
rect 4596 23984 4598 24003
rect 4561 23983 4619 23984
rect 4692 23983 4694 24003
rect 4932 23983 4934 24003
rect 4980 23983 4982 24003
rect 5028 23983 5030 24003
rect 5124 23983 5126 24003
rect 5220 23983 5222 24003
rect 5460 23983 5462 24003
rect 5508 23983 5510 24003
rect 5556 23983 5558 24003
rect 5652 23983 5654 24003
rect 5748 23983 5750 24003
rect 5796 23983 5798 24003
rect 5844 23983 5846 24003
rect 5892 23983 5894 24003
rect 6276 23983 6278 24003
rect 6300 23983 6302 24003
rect 6372 23983 6374 24003
rect 6396 23983 6398 24003
rect 6492 23983 6494 24003
rect 6516 23983 6518 24003
rect 6588 23983 6590 24003
rect 6612 23983 6614 24003
rect 6636 23983 6638 24003
rect 6708 23983 6710 24003
rect 6804 23983 6806 24003
rect 6900 23983 6902 24003
rect 7164 23983 7166 24003
rect 7284 23983 7286 24003
rect 7380 23983 7382 24003
rect 7404 23983 7406 24003
rect 7476 23983 7478 24003
rect 7500 23983 7502 24003
rect 7572 23983 7574 24003
rect 7596 23983 7598 24003
rect 7668 23983 7670 24003
rect 7692 23983 7694 24003
rect 7908 23983 7910 24003
rect 8124 23983 8126 24003
rect 8220 23983 8222 24003
rect 8316 23983 8318 24003
rect 8412 23983 8414 24003
rect 8700 23983 8702 24003
rect 8748 23983 8750 24003
rect 8796 23983 8798 24003
rect 8844 23983 8846 24003
rect 8868 23983 8870 24003
rect 9516 23983 9518 24003
rect 9660 23983 9662 24003
rect 9684 23983 9686 24003
rect 9780 23983 9782 24003
rect 9804 23983 9806 24003
rect 9828 23983 9830 24003
rect 10044 23983 10046 24003
rect 10140 23983 10142 24003
rect 10236 23983 10238 24003
rect 10332 23983 10334 24003
rect 10380 23983 10382 24003
rect 10428 23983 10430 24003
rect 10524 23983 10526 24003
rect 10548 23983 10550 24003
rect 10620 23983 10622 24003
rect 10644 23983 10646 24003
rect 10716 23983 10718 24003
rect 10860 23983 10862 24003
rect 10956 23983 10958 24003
rect 11052 23983 11054 24003
rect 11100 23983 11102 24003
rect 11172 23983 11174 24003
rect 11220 23983 11222 24003
rect 11340 23983 11342 24003
rect 11436 23983 11438 24003
rect 11676 23983 11678 24003
rect 11724 23983 11726 24003
rect 11772 23984 11774 24003
rect 11761 23983 11795 23984
rect 11796 23983 11798 24003
rect 12060 23983 12062 24003
rect 12276 23983 12278 24003
rect 12372 23983 12374 24003
rect 12409 23983 12443 23984
rect 12468 23983 12470 24003
rect 12564 23983 12566 24003
rect 12780 23983 12782 24003
rect 12876 23983 12878 24003
rect 12972 23983 12974 24003
rect 13044 23983 13046 24003
rect 13068 23983 13070 24003
rect 13164 23983 13166 24003
rect 13249 23998 13252 24003
rect 13259 23984 13262 23998
rect 13260 23983 13262 23984
rect 13332 23983 13334 24003
rect 13356 23983 13359 24000
rect 13500 23983 13502 24003
rect 13572 23983 13574 24003
rect 13836 23983 13838 24003
rect 13932 23983 13934 24003
rect 14004 23983 14006 24003
rect 14028 23983 14030 24003
rect 14100 23984 14102 24003
rect 14065 23983 14123 23984
rect 14940 23983 14942 24003
rect 15036 23983 15038 24003
rect 15276 23983 15278 24003
rect 15372 23983 15374 24003
rect 15420 23983 15422 24003
rect 15468 23983 15470 24003
rect 15564 23983 15566 24003
rect 15660 23983 15662 24003
rect 15684 23983 15686 24003
rect 15732 23983 15734 24003
rect 15756 23983 15758 24003
rect 15759 24000 15773 24003
rect 15783 24003 20603 24007
rect 15783 24000 15797 24003
rect 15804 24000 15807 24003
rect 15828 23983 15830 24003
rect 15852 23983 15854 24003
rect 15948 23983 15950 24003
rect 15972 23983 15974 24003
rect 16044 23983 16046 24003
rect 16068 23983 16070 24003
rect 16164 23983 16166 24003
rect 16260 23983 16262 24003
rect 16284 23983 16286 24003
rect 16380 23983 16382 24003
rect 16476 23983 16478 24003
rect 16548 23983 16550 24003
rect 16572 23983 16574 24003
rect 16596 23983 16598 24003
rect 16668 23983 16670 24003
rect 16692 23983 16694 24003
rect 16764 23983 16766 24003
rect 16788 23983 16790 24003
rect 16884 23983 16886 24003
rect 16908 23983 16910 24003
rect 17028 23983 17030 24003
rect 17124 23983 17126 24003
rect 17196 23983 17198 24003
rect 17220 23983 17222 24003
rect 17292 23983 17294 24003
rect 17316 23983 17318 24003
rect 17964 23983 17966 24003
rect 18060 23983 18062 24003
rect 18132 23983 18134 24003
rect 18228 23983 18230 24003
rect 18492 23983 18494 24003
rect 18540 23983 18542 24003
rect 18601 23983 18635 23984
rect 18636 23983 18638 24003
rect 18732 23983 18734 24003
rect 18828 23983 18830 24003
rect 18924 23983 18926 24003
rect 18972 23983 18974 24003
rect 19020 23983 19022 24003
rect 19068 23983 19070 24003
rect 19140 23983 19142 24003
rect 19164 23983 19166 24003
rect 19236 23983 19238 24003
rect 19260 23983 19262 24003
rect 19788 23983 19790 24003
rect 19836 23983 19838 24003
rect 19860 23983 19862 24003
rect 19884 23983 19886 24003
rect 19980 23983 19982 24003
rect 20004 23983 20006 24003
rect 20076 23983 20078 24003
rect 20100 23983 20102 24003
rect 20172 23983 20174 24003
rect 20196 23983 20198 24003
rect 20292 23984 20294 24003
rect 20388 23984 20390 24003
rect 20401 23998 20404 24003
rect 20412 23998 20414 24003
rect 20497 23998 20500 24003
rect 20508 24000 20510 24003
rect 20508 23998 20511 24000
rect 20411 23984 20414 23998
rect 20507 23990 20511 23998
rect 20521 23998 20524 24003
rect 20532 24000 20534 24003
rect 20532 23998 20535 24000
rect 20521 23990 20525 23998
rect 20507 23984 20521 23990
rect 20531 23984 20535 23998
rect 20593 23990 20597 23998
rect 20583 23984 20593 23990
rect 20281 23983 20339 23984
rect 20377 23983 20411 23984
rect -4727 23979 13349 23983
rect -4727 23976 -4723 23979
rect -4716 23976 -4713 23979
rect -4620 23976 -4618 23979
rect -4620 23960 -4617 23976
rect -4631 23959 -4597 23960
rect -4284 23959 -4282 23979
rect -3876 23976 -3874 23979
rect -3876 23959 -3873 23976
rect -3828 23959 -3826 23979
rect -3609 23976 -3595 23979
rect -3540 23959 -3538 23979
rect -3468 23959 -3466 23979
rect -3324 23959 -3322 23979
rect -3108 23959 -3106 23979
rect -3012 23959 -3010 23979
rect -2988 23959 -2986 23979
rect -2916 23959 -2914 23979
rect -2868 23959 -2866 23979
rect -2772 23959 -2770 23979
rect -2364 23959 -2362 23979
rect -1908 23959 -1906 23979
rect -1452 23959 -1450 23979
rect -1356 23959 -1354 23979
rect -1332 23959 -1329 23976
rect -1260 23959 -1258 23979
rect -1236 23959 -1234 23979
rect -1140 23959 -1138 23979
rect -876 23959 -874 23979
rect -780 23959 -778 23979
rect -564 23959 -562 23979
rect -468 23959 -466 23979
rect -12 23959 -10 23979
rect 84 23959 86 23979
rect 180 23959 182 23979
rect 348 23959 350 23979
rect 468 23959 470 23979
rect 492 23959 494 23979
rect 564 23959 566 23979
rect 588 23959 590 23979
rect 660 23959 662 23979
rect 948 23959 950 23979
rect 1044 23959 1046 23979
rect 1092 23959 1094 23979
rect 1140 23959 1142 23979
rect 1308 23959 1310 23979
rect 1356 23959 1358 23979
rect 1503 23976 1517 23979
rect 1572 23959 1574 23979
rect 1860 23959 1862 23979
rect 1956 23959 1958 23979
rect 2052 23959 2054 23979
rect 2148 23959 2150 23979
rect 2244 23959 2246 23979
rect 2340 23959 2342 23979
rect 2436 23959 2438 23979
rect 2532 23959 2534 23979
rect 2628 23959 2630 23979
rect 2724 23959 2726 23979
rect 2940 23959 2942 23979
rect 2988 23959 2990 23979
rect 3324 23959 3326 23979
rect 3540 23959 3542 23979
rect 3780 23959 3782 23979
rect 4057 23959 4115 23960
rect 4188 23959 4190 23979
rect 4308 23959 4310 23979
rect 4479 23976 4493 23979
rect 4500 23976 4503 23979
rect 4585 23974 4588 23979
rect 4596 23974 4598 23979
rect 4595 23960 4598 23974
rect 4692 23976 4694 23979
rect 4692 23959 4695 23976
rect 4932 23959 4934 23979
rect 4980 23959 4982 23979
rect 5028 23959 5030 23979
rect 5124 23959 5126 23979
rect 5220 23959 5222 23979
rect 5460 23959 5462 23979
rect 5508 23959 5510 23979
rect 5556 23959 5558 23979
rect 5652 23959 5654 23979
rect 5748 23959 5750 23979
rect 5796 23959 5798 23979
rect 5844 23959 5846 23979
rect 5892 23959 5894 23979
rect 6276 23959 6278 23979
rect 6300 23959 6302 23979
rect 6372 23959 6374 23979
rect 6396 23959 6398 23979
rect 6492 23959 6494 23979
rect 6516 23959 6518 23979
rect 6588 23959 6590 23979
rect 6612 23959 6614 23979
rect 6636 23959 6638 23979
rect 6708 23959 6710 23979
rect 6804 23959 6806 23979
rect 6900 23959 6902 23979
rect 7164 23959 7166 23979
rect 7284 23959 7286 23979
rect 7380 23959 7382 23979
rect 7404 23959 7406 23979
rect 7476 23959 7478 23979
rect 7500 23959 7502 23979
rect 7572 23959 7574 23979
rect 7596 23959 7598 23979
rect 7668 23959 7670 23979
rect 7692 23959 7694 23979
rect 7908 23959 7910 23979
rect 8124 23959 8126 23979
rect 8220 23959 8222 23979
rect 8316 23959 8318 23979
rect 8412 23959 8414 23979
rect 8700 23959 8702 23979
rect 8748 23959 8750 23979
rect 8796 23959 8798 23979
rect 8844 23959 8846 23979
rect 8868 23959 8870 23979
rect 9087 23976 9101 23979
rect 9516 23959 9518 23979
rect 9660 23959 9662 23979
rect 9684 23959 9686 23979
rect 9780 23959 9782 23979
rect 9804 23959 9806 23979
rect 9828 23959 9830 23979
rect 10044 23959 10046 23979
rect 10140 23959 10142 23979
rect 10236 23959 10238 23979
rect 10332 23959 10334 23979
rect 10380 23959 10382 23979
rect 10428 23959 10430 23979
rect 10524 23959 10526 23979
rect 10548 23959 10550 23979
rect 10620 23959 10622 23979
rect 10644 23959 10646 23979
rect 10716 23959 10718 23979
rect 10860 23959 10862 23979
rect 10956 23959 10958 23979
rect 11052 23959 11054 23979
rect 11100 23959 11102 23979
rect 11172 23959 11174 23979
rect 11220 23959 11222 23979
rect 11340 23959 11342 23979
rect 11436 23959 11438 23979
rect 11676 23959 11678 23979
rect 11724 23959 11726 23979
rect 11761 23974 11764 23979
rect 11772 23974 11774 23979
rect 11771 23960 11774 23974
rect 11796 23959 11798 23979
rect 12060 23959 12062 23979
rect 12276 23959 12278 23979
rect 12372 23959 12374 23979
rect 12468 23959 12470 23979
rect 12564 23959 12566 23979
rect 12780 23959 12782 23979
rect 12876 23959 12878 23979
rect 12972 23959 12974 23979
rect 13044 23959 13046 23979
rect 13068 23959 13070 23979
rect 13164 23959 13166 23979
rect 13260 23959 13262 23979
rect 13332 23959 13334 23979
rect 13335 23976 13349 23979
rect 13356 23979 20411 23983
rect 13356 23976 13373 23979
rect 13356 23959 13358 23976
rect 13500 23959 13502 23979
rect 13572 23959 13574 23979
rect 13836 23959 13838 23979
rect 13932 23959 13934 23979
rect 14004 23959 14006 23979
rect 14028 23959 14030 23979
rect 14089 23974 14092 23979
rect 14100 23974 14102 23979
rect 14099 23960 14102 23974
rect 14172 23959 14175 23976
rect 14940 23959 14942 23979
rect 15036 23959 15038 23979
rect 15276 23959 15278 23979
rect 15372 23959 15374 23979
rect 15420 23959 15422 23979
rect 15468 23959 15470 23979
rect 15564 23959 15566 23979
rect 15660 23959 15662 23979
rect 15684 23959 15686 23979
rect 15732 23959 15734 23979
rect 15756 23959 15758 23979
rect 15769 23959 15827 23960
rect 15828 23959 15830 23979
rect 15852 23959 15854 23979
rect 15948 23959 15950 23979
rect 15972 23959 15974 23979
rect 16044 23959 16046 23979
rect 16068 23959 16070 23979
rect 16164 23959 16166 23979
rect 16260 23959 16262 23979
rect 16284 23959 16286 23979
rect 16380 23959 16382 23979
rect 16476 23959 16478 23979
rect 16548 23959 16550 23979
rect 16572 23959 16574 23979
rect 16596 23959 16598 23979
rect 16668 23959 16670 23979
rect 16692 23959 16694 23979
rect 16764 23959 16766 23979
rect 16788 23959 16790 23979
rect 16884 23959 16886 23979
rect 16908 23959 16910 23979
rect 17028 23959 17030 23979
rect 17124 23959 17126 23979
rect 17196 23959 17198 23979
rect 17220 23959 17222 23979
rect 17292 23959 17294 23979
rect 17316 23959 17318 23979
rect 17964 23959 17966 23979
rect 18060 23959 18062 23979
rect 18132 23959 18134 23979
rect 18228 23959 18230 23979
rect 18492 23959 18494 23979
rect 18540 23959 18542 23979
rect 18636 23959 18638 23979
rect 18732 23959 18734 23979
rect 18828 23959 18830 23979
rect 18924 23959 18926 23979
rect 18972 23959 18974 23979
rect 19020 23959 19022 23979
rect 19068 23959 19070 23979
rect 19140 23959 19142 23979
rect 19164 23959 19166 23979
rect 19236 23959 19238 23979
rect 19260 23959 19262 23979
rect 19788 23959 19790 23979
rect 19836 23959 19838 23979
rect 19860 23959 19862 23979
rect 19884 23959 19886 23979
rect 19980 23959 19982 23979
rect 20004 23959 20006 23979
rect 20076 23959 20078 23979
rect 20100 23959 20102 23979
rect 20172 23959 20174 23979
rect 20196 23960 20198 23979
rect 20281 23974 20284 23979
rect 20292 23974 20294 23979
rect 20377 23974 20380 23979
rect 20388 23976 20390 23979
rect 20388 23974 20391 23976
rect 20291 23960 20294 23974
rect 20387 23966 20391 23974
rect 20401 23966 20405 23974
rect 20387 23960 20401 23966
rect 20185 23959 20219 23960
rect -4631 23955 -1339 23959
rect -4631 23952 -4627 23955
rect -4620 23952 -4617 23955
rect -4511 23935 -4477 23936
rect -4284 23935 -4282 23955
rect -3897 23952 -3883 23955
rect -3876 23952 -3873 23955
rect -3828 23935 -3826 23955
rect -3540 23935 -3538 23955
rect -3468 23935 -3466 23955
rect -3324 23935 -3322 23955
rect -3108 23935 -3106 23955
rect -3012 23935 -3010 23955
rect -2988 23935 -2986 23955
rect -2916 23935 -2914 23955
rect -2868 23935 -2866 23955
rect -2772 23935 -2770 23955
rect -2615 23935 -2581 23936
rect -2364 23935 -2362 23955
rect -1908 23935 -1906 23955
rect -1452 23935 -1450 23955
rect -1356 23935 -1354 23955
rect -1353 23952 -1339 23955
rect -1332 23955 4661 23959
rect -1332 23952 -1315 23955
rect -1332 23935 -1330 23952
rect -1260 23935 -1258 23955
rect -1236 23935 -1234 23955
rect -1140 23935 -1138 23955
rect -876 23935 -874 23955
rect -780 23935 -778 23955
rect -564 23935 -562 23955
rect -468 23935 -466 23955
rect -12 23935 -10 23955
rect 84 23935 86 23955
rect 180 23935 182 23955
rect 348 23935 350 23955
rect 468 23935 470 23955
rect 492 23935 494 23955
rect 564 23935 566 23955
rect 588 23935 590 23955
rect 660 23935 662 23955
rect 948 23935 950 23955
rect 1044 23935 1046 23955
rect 1092 23935 1094 23955
rect 1140 23935 1142 23955
rect 1308 23935 1310 23955
rect 1356 23935 1358 23955
rect 1572 23935 1574 23955
rect 1860 23935 1862 23955
rect 1956 23935 1958 23955
rect 2052 23935 2054 23955
rect 2148 23935 2150 23955
rect 2244 23935 2246 23955
rect 2340 23935 2342 23955
rect 2436 23935 2438 23955
rect 2532 23935 2534 23955
rect 2628 23935 2630 23955
rect 2665 23935 2699 23936
rect 2724 23935 2726 23955
rect 2940 23935 2942 23955
rect 2988 23935 2990 23955
rect 3324 23935 3326 23955
rect 3540 23935 3542 23955
rect 3780 23935 3782 23955
rect 4057 23950 4060 23955
rect 4188 23952 4190 23955
rect 4067 23936 4070 23950
rect 4068 23935 4070 23936
rect 4188 23935 4191 23952
rect 4308 23935 4310 23955
rect 4647 23952 4661 23955
rect 4671 23955 14165 23959
rect 4671 23952 4685 23955
rect 4692 23952 4695 23955
rect 4932 23935 4934 23955
rect 4980 23935 4982 23955
rect 5028 23935 5030 23955
rect 5124 23935 5126 23955
rect 5220 23935 5222 23955
rect 5460 23935 5462 23955
rect 5508 23935 5510 23955
rect 5556 23935 5558 23955
rect 5652 23935 5654 23955
rect 5748 23935 5750 23955
rect 5796 23935 5798 23955
rect 5844 23935 5846 23955
rect 5892 23935 5894 23955
rect 6276 23935 6278 23955
rect 6300 23935 6302 23955
rect 6372 23935 6374 23955
rect 6396 23935 6398 23955
rect 6492 23935 6494 23955
rect 6516 23935 6518 23955
rect 6588 23935 6590 23955
rect 6612 23935 6614 23955
rect 6636 23935 6638 23955
rect 6708 23935 6710 23955
rect 6804 23935 6806 23955
rect 6900 23935 6902 23955
rect 7009 23935 7043 23936
rect 7164 23935 7166 23955
rect 7284 23935 7286 23955
rect 7380 23935 7382 23955
rect 7404 23935 7406 23955
rect 7476 23935 7478 23955
rect 7500 23935 7502 23955
rect 7572 23935 7574 23955
rect 7596 23935 7598 23955
rect 7668 23935 7670 23955
rect 7692 23935 7694 23955
rect 7908 23935 7910 23955
rect 8124 23935 8126 23955
rect 8220 23935 8222 23955
rect 8316 23935 8318 23955
rect 8412 23935 8414 23955
rect 8700 23935 8702 23955
rect 8748 23935 8750 23955
rect 8796 23935 8798 23955
rect 8844 23935 8846 23955
rect 8868 23935 8870 23955
rect 9516 23935 9518 23955
rect 9660 23935 9662 23955
rect 9684 23935 9686 23955
rect 9780 23935 9782 23955
rect 9804 23935 9806 23955
rect 9828 23935 9830 23955
rect 10044 23935 10046 23955
rect 10140 23935 10142 23955
rect 10236 23935 10238 23955
rect 10332 23935 10334 23955
rect 10380 23935 10382 23955
rect 10428 23935 10430 23955
rect 10524 23935 10526 23955
rect 10548 23935 10550 23955
rect 10620 23935 10622 23955
rect 10644 23935 10646 23955
rect 10716 23935 10718 23955
rect 10860 23935 10862 23955
rect 10956 23935 10958 23955
rect 11052 23935 11054 23955
rect 11100 23935 11102 23955
rect 11172 23935 11174 23955
rect 11220 23935 11222 23955
rect 11340 23935 11342 23955
rect 11436 23935 11438 23955
rect 11676 23935 11678 23955
rect 11724 23935 11726 23955
rect 11796 23935 11798 23955
rect 11847 23952 11861 23955
rect 12060 23935 12062 23955
rect 12276 23935 12278 23955
rect 12372 23935 12374 23955
rect 12468 23935 12470 23955
rect 12495 23952 12509 23955
rect 12564 23935 12566 23955
rect 12780 23935 12782 23955
rect 12876 23935 12878 23955
rect 12972 23936 12974 23955
rect 12961 23935 12995 23936
rect 13044 23935 13046 23955
rect 13068 23935 13070 23955
rect 13164 23935 13166 23955
rect 13260 23935 13262 23955
rect 13332 23935 13334 23955
rect 13356 23935 13358 23955
rect 13500 23935 13502 23955
rect 13572 23935 13574 23955
rect 13836 23935 13838 23955
rect 13932 23935 13934 23955
rect 14004 23935 14006 23955
rect 14028 23935 14030 23955
rect 14151 23952 14165 23955
rect 14172 23955 20219 23959
rect 14172 23952 14189 23955
rect 14172 23935 14174 23952
rect 14940 23935 14942 23955
rect 15036 23935 15038 23955
rect 15276 23935 15278 23955
rect 15372 23935 15374 23955
rect 15420 23935 15422 23955
rect 15468 23935 15470 23955
rect 15564 23935 15566 23955
rect 15660 23935 15662 23955
rect 15684 23935 15686 23955
rect 15732 23935 15734 23955
rect 15756 23935 15758 23955
rect 15769 23950 15772 23955
rect 15779 23936 15782 23950
rect 15780 23935 15782 23936
rect 15828 23935 15830 23955
rect 15852 23935 15854 23955
rect 15876 23935 15879 23952
rect 15948 23935 15950 23955
rect 15972 23935 15974 23955
rect 16044 23935 16046 23955
rect 16068 23935 16070 23955
rect 16164 23935 16166 23955
rect 16260 23935 16262 23955
rect 16284 23935 16286 23955
rect 16380 23935 16382 23955
rect 16476 23935 16478 23955
rect 16548 23935 16550 23955
rect 16572 23935 16574 23955
rect 16596 23935 16598 23955
rect 16668 23935 16670 23955
rect 16692 23935 16694 23955
rect 16764 23935 16766 23955
rect 16788 23935 16790 23955
rect 16884 23935 16886 23955
rect 16908 23935 16910 23955
rect 17028 23935 17030 23955
rect 17124 23935 17126 23955
rect 17196 23935 17198 23955
rect 17220 23935 17222 23955
rect 17292 23935 17294 23955
rect 17316 23935 17318 23955
rect 17964 23935 17966 23955
rect 18060 23935 18062 23955
rect 18132 23935 18134 23955
rect 18228 23935 18230 23955
rect 18492 23935 18494 23955
rect 18540 23935 18542 23955
rect 18636 23935 18638 23955
rect 18687 23952 18701 23955
rect 18732 23935 18734 23955
rect 18828 23935 18830 23955
rect 18924 23935 18926 23955
rect 18972 23935 18974 23955
rect 19020 23935 19022 23955
rect 19068 23935 19070 23955
rect 19140 23935 19142 23955
rect 19164 23935 19166 23955
rect 19236 23935 19238 23955
rect 19260 23935 19262 23955
rect 19788 23935 19790 23955
rect 19836 23935 19838 23955
rect 19860 23935 19862 23955
rect 19884 23935 19886 23955
rect 19980 23935 19982 23955
rect 20004 23935 20006 23955
rect 20076 23935 20078 23955
rect 20100 23936 20102 23955
rect 20172 23936 20174 23955
rect 20185 23950 20188 23955
rect 20196 23950 20198 23955
rect 20195 23936 20198 23950
rect 20089 23935 20147 23936
rect 20161 23935 20195 23936
rect -4511 23931 4157 23935
rect -4284 23912 -4282 23931
rect -4391 23911 -4357 23912
rect -4319 23911 -4261 23912
rect -3828 23911 -3826 23931
rect -3540 23911 -3538 23931
rect -3468 23911 -3466 23931
rect -3455 23911 -3397 23912
rect -3324 23911 -3322 23931
rect -3108 23911 -3106 23931
rect -3012 23911 -3010 23931
rect -2988 23911 -2986 23931
rect -2916 23911 -2914 23931
rect -2868 23911 -2866 23931
rect -2772 23911 -2770 23931
rect -2364 23911 -2362 23931
rect -1908 23911 -1906 23931
rect -1452 23911 -1450 23931
rect -1356 23911 -1354 23931
rect -1332 23911 -1330 23931
rect -1260 23911 -1258 23931
rect -1236 23911 -1234 23931
rect -1140 23911 -1138 23931
rect -876 23911 -874 23931
rect -780 23911 -778 23931
rect -564 23911 -562 23931
rect -468 23911 -466 23931
rect -12 23911 -10 23931
rect 84 23911 86 23931
rect 180 23911 182 23931
rect 241 23911 275 23912
rect 348 23911 350 23931
rect 468 23911 470 23931
rect 492 23911 494 23931
rect 564 23911 566 23931
rect 588 23911 590 23931
rect 660 23911 662 23931
rect 697 23911 755 23912
rect 948 23911 950 23931
rect 1044 23911 1046 23931
rect 1092 23911 1094 23931
rect 1140 23911 1142 23931
rect 1308 23911 1310 23931
rect 1356 23911 1358 23931
rect 1572 23911 1574 23931
rect 1860 23911 1862 23931
rect 1956 23911 1958 23931
rect 2052 23911 2054 23931
rect 2148 23911 2150 23931
rect 2244 23911 2246 23931
rect 2340 23911 2342 23931
rect 2436 23911 2438 23931
rect 2532 23911 2534 23931
rect 2628 23911 2630 23931
rect 2724 23911 2726 23931
rect 2940 23911 2942 23931
rect 2988 23911 2990 23931
rect 3324 23911 3326 23931
rect 3540 23911 3542 23931
rect 3780 23911 3782 23931
rect 4068 23911 4070 23931
rect 4143 23928 4157 23931
rect 4167 23931 15869 23935
rect 4167 23928 4181 23931
rect 4188 23928 4191 23931
rect 4308 23911 4310 23931
rect 4932 23911 4934 23931
rect 4980 23911 4982 23931
rect 5028 23911 5030 23931
rect 5124 23911 5126 23931
rect 5137 23911 5195 23912
rect 5220 23911 5222 23931
rect 5460 23911 5462 23931
rect 5508 23911 5510 23931
rect 5556 23911 5558 23931
rect 5652 23911 5654 23931
rect 5748 23911 5750 23931
rect 5796 23911 5798 23931
rect 5844 23911 5846 23931
rect 5892 23911 5894 23931
rect 6276 23911 6278 23931
rect 6300 23911 6302 23931
rect 6372 23911 6374 23931
rect 6396 23911 6398 23931
rect 6492 23911 6494 23931
rect 6516 23911 6518 23931
rect 6588 23911 6590 23931
rect 6612 23911 6614 23931
rect 6636 23911 6638 23931
rect 6708 23911 6710 23931
rect 6804 23911 6806 23931
rect 6900 23911 6902 23931
rect 7164 23911 7166 23931
rect 7284 23911 7286 23931
rect 7380 23911 7382 23931
rect 7404 23911 7406 23931
rect 7476 23911 7478 23931
rect 7500 23911 7502 23931
rect 7572 23911 7574 23931
rect 7596 23911 7598 23931
rect 7668 23911 7670 23931
rect 7692 23911 7694 23931
rect 7908 23911 7910 23931
rect 8124 23911 8126 23931
rect 8220 23911 8222 23931
rect 8316 23911 8318 23931
rect 8412 23911 8414 23931
rect 8700 23911 8702 23931
rect 8748 23911 8750 23931
rect 8796 23911 8798 23931
rect 8844 23911 8846 23931
rect 8868 23911 8870 23931
rect 9516 23911 9518 23931
rect 9660 23911 9662 23931
rect 9684 23911 9686 23931
rect 9780 23911 9782 23931
rect 9804 23911 9806 23931
rect 9828 23911 9830 23931
rect 10044 23911 10046 23931
rect 10140 23911 10142 23931
rect 10236 23911 10238 23931
rect 10332 23911 10334 23931
rect 10380 23911 10382 23931
rect 10428 23911 10430 23931
rect 10524 23911 10526 23931
rect 10548 23911 10550 23931
rect 10620 23911 10622 23931
rect 10644 23911 10646 23931
rect 10716 23911 10718 23931
rect 10860 23911 10862 23931
rect 10956 23911 10958 23931
rect 11052 23911 11054 23931
rect 11100 23911 11102 23931
rect 11172 23911 11174 23931
rect 11220 23911 11222 23931
rect 11340 23911 11342 23931
rect 11436 23912 11438 23931
rect 11401 23911 11459 23912
rect 11676 23911 11678 23931
rect 11724 23911 11726 23931
rect 11796 23911 11798 23931
rect 12060 23911 12062 23931
rect 12276 23911 12278 23931
rect 12372 23911 12374 23931
rect 12468 23911 12470 23931
rect 12564 23911 12566 23931
rect 12780 23911 12782 23931
rect 12876 23911 12878 23931
rect 12961 23926 12964 23931
rect 12972 23926 12974 23931
rect 12971 23912 12974 23926
rect 13044 23911 13046 23931
rect 13068 23928 13070 23931
rect 13068 23911 13071 23928
rect 13164 23911 13166 23931
rect 13260 23911 13262 23931
rect 13332 23911 13334 23931
rect 13356 23911 13358 23931
rect 13500 23911 13502 23931
rect 13572 23911 13574 23931
rect 13836 23911 13838 23931
rect 13932 23911 13934 23931
rect 14004 23911 14006 23931
rect 14028 23911 14030 23931
rect 14172 23911 14174 23931
rect 14940 23911 14942 23931
rect 15036 23911 15038 23931
rect 15276 23911 15278 23931
rect 15372 23911 15374 23931
rect 15420 23911 15422 23931
rect 15468 23911 15470 23931
rect 15564 23911 15566 23931
rect 15660 23911 15662 23931
rect 15684 23911 15686 23931
rect 15732 23911 15734 23931
rect 15756 23911 15758 23931
rect 15780 23911 15782 23931
rect 15828 23911 15830 23931
rect 15852 23911 15854 23931
rect 15855 23928 15869 23931
rect 15876 23931 20195 23935
rect 15876 23928 15893 23931
rect 15876 23911 15878 23928
rect 15948 23911 15950 23931
rect 15972 23911 15974 23931
rect 16044 23911 16046 23931
rect 16068 23911 16070 23931
rect 16164 23911 16166 23931
rect 16260 23911 16262 23931
rect 16284 23911 16286 23931
rect 16380 23911 16382 23931
rect 16476 23911 16478 23931
rect 16548 23911 16550 23931
rect 16572 23912 16574 23931
rect 16561 23911 16595 23912
rect 16596 23911 16598 23931
rect 16668 23911 16670 23931
rect 16692 23911 16694 23931
rect 16764 23911 16766 23931
rect 16788 23911 16790 23931
rect 16884 23911 16886 23931
rect 16908 23911 16910 23931
rect 17028 23911 17030 23931
rect 17124 23911 17126 23931
rect 17196 23911 17198 23931
rect 17220 23911 17222 23931
rect 17292 23911 17294 23931
rect 17316 23911 17318 23931
rect 17964 23911 17966 23931
rect 18060 23911 18062 23931
rect 18132 23911 18134 23931
rect 18228 23911 18230 23931
rect 18492 23911 18494 23931
rect 18540 23911 18542 23931
rect 18636 23911 18638 23931
rect 18732 23911 18734 23931
rect 18828 23911 18830 23931
rect 18924 23911 18926 23931
rect 18972 23911 18974 23931
rect 19020 23911 19022 23931
rect 19068 23911 19070 23931
rect 19140 23911 19142 23931
rect 19164 23911 19166 23931
rect 19236 23911 19238 23931
rect 19260 23911 19262 23931
rect 19788 23911 19790 23931
rect 19836 23911 19838 23931
rect 19860 23912 19862 23931
rect 19849 23911 19883 23912
rect 19884 23911 19886 23931
rect 19980 23911 19982 23931
rect 20004 23911 20006 23931
rect 20076 23912 20078 23931
rect 20089 23926 20092 23931
rect 20100 23926 20102 23931
rect 20161 23926 20164 23931
rect 20172 23926 20174 23931
rect 20099 23912 20102 23926
rect 20171 23912 20174 23926
rect 20185 23918 20189 23926
rect 20175 23912 20185 23918
rect 20065 23911 20099 23912
rect -4391 23907 20099 23911
rect -4295 23902 -4292 23907
rect -4284 23904 -4282 23907
rect -4284 23902 -4281 23904
rect -4295 23894 -4291 23902
rect -4305 23888 -4295 23894
rect -4285 23888 -4281 23902
rect -3828 23888 -3826 23907
rect -4175 23887 -4141 23888
rect -4103 23887 -4069 23888
rect -4175 23883 -4069 23887
rect -4055 23887 -4021 23888
rect -3839 23887 -3805 23888
rect -4055 23883 -3805 23887
rect -3767 23887 -3733 23888
rect -3540 23887 -3538 23907
rect -3468 23887 -3466 23907
rect -3455 23902 -3452 23907
rect -3324 23904 -3322 23907
rect -3445 23888 -3442 23902
rect -3444 23887 -3442 23888
rect -3324 23887 -3321 23904
rect -3108 23887 -3106 23907
rect -3012 23887 -3010 23907
rect -2988 23888 -2986 23907
rect -2916 23888 -2914 23907
rect -2868 23888 -2866 23907
rect -2999 23887 -2941 23888
rect -2927 23887 -2893 23888
rect -3767 23883 -3355 23887
rect -3839 23878 -3836 23883
rect -3828 23878 -3826 23883
rect -4079 23870 -4075 23878
rect -4089 23864 -4079 23870
rect -3829 23864 -3826 23878
rect -3743 23870 -3739 23878
rect -3753 23864 -3743 23870
rect -3540 23864 -3538 23883
rect -3468 23864 -3466 23883
rect -3444 23864 -3442 23883
rect -3369 23880 -3355 23883
rect -3345 23883 -2893 23887
rect -2879 23887 -2845 23888
rect -2772 23887 -2770 23907
rect -2529 23904 -2515 23907
rect -2364 23887 -2362 23907
rect -1908 23887 -1906 23907
rect -1452 23887 -1450 23907
rect -1356 23887 -1354 23907
rect -1332 23887 -1330 23907
rect -1260 23887 -1258 23907
rect -1236 23887 -1234 23907
rect -1140 23887 -1138 23907
rect -876 23887 -874 23907
rect -780 23887 -778 23907
rect -564 23887 -562 23907
rect -468 23887 -466 23907
rect -12 23887 -10 23907
rect 84 23887 86 23907
rect 180 23887 182 23907
rect 348 23904 350 23907
rect 348 23887 351 23904
rect 468 23887 470 23907
rect 492 23887 494 23907
rect 564 23887 566 23907
rect 588 23887 590 23907
rect 660 23887 662 23907
rect 697 23902 700 23907
rect 707 23888 710 23902
rect 708 23887 710 23888
rect 948 23887 950 23907
rect 1044 23887 1046 23907
rect 1092 23887 1094 23907
rect 1140 23887 1142 23907
rect 1308 23887 1310 23907
rect 1356 23887 1358 23907
rect 1572 23887 1574 23907
rect 1860 23887 1862 23907
rect 1956 23887 1958 23907
rect 2052 23887 2054 23907
rect 2148 23887 2150 23907
rect 2244 23887 2246 23907
rect 2340 23887 2342 23907
rect 2436 23887 2438 23907
rect 2532 23887 2534 23907
rect 2628 23887 2630 23907
rect 2724 23887 2726 23907
rect 2751 23904 2765 23907
rect 2940 23887 2942 23907
rect 2988 23887 2990 23907
rect 3169 23887 3203 23888
rect 3324 23887 3326 23907
rect 3540 23887 3542 23907
rect 3721 23887 3755 23888
rect 3780 23887 3782 23907
rect 4068 23887 4070 23907
rect 4308 23887 4310 23907
rect 4932 23887 4934 23907
rect 4980 23887 4982 23907
rect 5028 23887 5030 23907
rect 5124 23887 5126 23907
rect 5137 23902 5140 23907
rect 5147 23888 5150 23902
rect 5148 23887 5150 23888
rect 5220 23887 5222 23907
rect 5244 23887 5247 23904
rect 5460 23887 5462 23907
rect 5508 23887 5510 23907
rect 5556 23887 5558 23907
rect 5652 23887 5654 23907
rect 5748 23887 5750 23907
rect 5796 23887 5798 23907
rect 5844 23887 5846 23907
rect 5892 23887 5894 23907
rect 6276 23887 6278 23907
rect 6300 23887 6302 23907
rect 6372 23887 6374 23907
rect 6396 23887 6398 23907
rect 6492 23887 6494 23907
rect 6516 23887 6518 23907
rect 6588 23887 6590 23907
rect 6612 23887 6614 23907
rect 6636 23887 6638 23907
rect 6708 23887 6710 23907
rect 6804 23887 6806 23907
rect 6900 23887 6902 23907
rect 7095 23904 7109 23907
rect 7164 23887 7166 23907
rect 7225 23887 7259 23888
rect 7284 23887 7286 23907
rect 7380 23887 7382 23907
rect 7404 23887 7406 23907
rect 7476 23887 7478 23907
rect 7500 23887 7502 23907
rect 7572 23887 7574 23907
rect 7596 23887 7598 23907
rect 7668 23887 7670 23907
rect 7692 23887 7694 23907
rect 7908 23887 7910 23907
rect 8124 23887 8126 23907
rect 8220 23887 8222 23907
rect 8316 23887 8318 23907
rect 8412 23887 8414 23907
rect 8700 23887 8702 23907
rect 8748 23887 8750 23907
rect 8796 23887 8798 23907
rect 8844 23887 8846 23907
rect 8868 23887 8870 23907
rect 9516 23887 9518 23907
rect 9553 23887 9587 23888
rect 9660 23887 9662 23907
rect 9684 23887 9686 23907
rect 9780 23887 9782 23907
rect 9804 23887 9806 23907
rect 9828 23887 9830 23907
rect 10044 23887 10046 23907
rect 10140 23887 10142 23907
rect 10236 23887 10238 23907
rect 10332 23887 10334 23907
rect 10380 23887 10382 23907
rect 10428 23887 10430 23907
rect 10524 23887 10526 23907
rect 10548 23887 10550 23907
rect 10620 23887 10622 23907
rect 10644 23887 10646 23907
rect 10716 23887 10718 23907
rect 10860 23887 10862 23907
rect 10956 23887 10958 23907
rect 11052 23887 11054 23907
rect 11100 23887 11102 23907
rect 11172 23887 11174 23907
rect 11220 23887 11222 23907
rect 11340 23887 11342 23907
rect 11425 23902 11428 23907
rect 11436 23902 11438 23907
rect 11435 23888 11438 23902
rect 11508 23887 11511 23904
rect 11676 23887 11678 23907
rect 11724 23887 11726 23907
rect 11796 23887 11798 23907
rect 12060 23887 12062 23907
rect 12276 23887 12278 23907
rect 12372 23887 12374 23907
rect 12468 23887 12470 23907
rect 12564 23887 12566 23907
rect 12780 23887 12782 23907
rect 12876 23887 12878 23907
rect 13044 23887 13046 23907
rect 13047 23904 13061 23907
rect 13068 23904 13071 23907
rect 13164 23887 13166 23907
rect 13260 23887 13262 23907
rect 13332 23887 13334 23907
rect 13356 23887 13358 23907
rect 13500 23887 13502 23907
rect 13572 23887 13574 23907
rect 13836 23887 13838 23907
rect 13932 23887 13934 23907
rect 14004 23887 14006 23907
rect 14028 23887 14030 23907
rect 14172 23887 14174 23907
rect 14940 23887 14942 23907
rect 15036 23887 15038 23907
rect 15276 23887 15278 23907
rect 15372 23887 15374 23907
rect 15420 23888 15422 23907
rect 15409 23887 15443 23888
rect 15468 23887 15470 23907
rect 15564 23887 15566 23907
rect 15660 23887 15662 23907
rect 15684 23887 15686 23907
rect 15732 23887 15734 23907
rect 15756 23887 15758 23907
rect 15780 23887 15782 23907
rect 15828 23887 15830 23907
rect 15852 23887 15854 23907
rect 15876 23887 15878 23907
rect 15948 23887 15950 23907
rect 15972 23887 15974 23907
rect 16044 23887 16046 23907
rect 16068 23887 16070 23907
rect 16164 23887 16166 23907
rect 16260 23887 16262 23907
rect 16284 23887 16286 23907
rect 16380 23887 16382 23907
rect 16476 23887 16478 23907
rect 16548 23887 16550 23907
rect 16561 23902 16564 23907
rect 16572 23902 16574 23907
rect 16571 23888 16574 23902
rect 16596 23887 16598 23907
rect 16668 23904 16670 23907
rect 16668 23887 16671 23904
rect 16692 23887 16694 23907
rect 16764 23887 16766 23907
rect 16788 23887 16790 23907
rect 16884 23887 16886 23907
rect 16908 23887 16910 23907
rect 17028 23887 17030 23907
rect 17124 23887 17126 23907
rect 17196 23887 17198 23907
rect 17220 23887 17222 23907
rect 17292 23887 17294 23907
rect 17316 23887 17318 23907
rect 17964 23887 17966 23907
rect 18060 23887 18062 23907
rect 18132 23887 18134 23907
rect 18228 23887 18230 23907
rect 18492 23887 18494 23907
rect 18540 23887 18542 23907
rect 18636 23887 18638 23907
rect 18732 23887 18734 23907
rect 18828 23887 18830 23907
rect 18924 23887 18926 23907
rect 18972 23887 18974 23907
rect 19020 23887 19022 23907
rect 19068 23887 19070 23907
rect 19140 23887 19142 23907
rect 19164 23887 19166 23907
rect 19236 23887 19238 23907
rect 19260 23887 19262 23907
rect 19788 23887 19790 23907
rect 19836 23887 19838 23907
rect 19849 23902 19852 23907
rect 19860 23902 19862 23907
rect 19859 23888 19862 23902
rect 19884 23888 19886 23907
rect 19980 23888 19982 23907
rect 20004 23888 20006 23907
rect 20065 23902 20068 23907
rect 20076 23902 20078 23907
rect 20075 23888 20078 23902
rect 19873 23887 19931 23888
rect 19969 23887 20027 23888
rect 20041 23887 20075 23888
rect -2879 23883 797 23887
rect -3345 23880 -3331 23883
rect -3324 23880 -3321 23883
rect -3108 23864 -3106 23883
rect -3012 23864 -3010 23883
rect -2999 23878 -2996 23883
rect -2988 23878 -2986 23883
rect -2927 23878 -2924 23883
rect -2916 23878 -2914 23883
rect -2879 23878 -2876 23883
rect -2868 23880 -2866 23883
rect -2772 23880 -2770 23883
rect -2868 23878 -2865 23880
rect -2989 23864 -2986 23878
rect -2917 23864 -2914 23878
rect -2903 23870 -2899 23878
rect -2913 23864 -2903 23870
rect -2869 23864 -2865 23878
rect -2772 23864 -2769 23880
rect -3935 23863 -3901 23864
rect -3887 23863 -3853 23864
rect -3935 23859 -3853 23863
rect -3647 23863 -3613 23864
rect -3575 23863 -3517 23864
rect -3479 23863 -3421 23864
rect -3119 23863 -3061 23864
rect -3023 23863 -2989 23864
rect -3647 23859 -2989 23863
rect -2783 23863 -2749 23864
rect -2364 23863 -2362 23883
rect -1908 23863 -1906 23883
rect -1452 23863 -1450 23883
rect -1356 23863 -1354 23883
rect -1332 23863 -1330 23883
rect -1260 23863 -1258 23883
rect -1236 23863 -1234 23883
rect -1140 23863 -1138 23883
rect -876 23863 -874 23883
rect -780 23863 -778 23883
rect -564 23863 -562 23883
rect -468 23863 -466 23883
rect -12 23863 -10 23883
rect 84 23863 86 23883
rect 180 23863 182 23883
rect 327 23880 341 23883
rect 348 23880 351 23883
rect 468 23863 470 23883
rect 492 23863 494 23883
rect 564 23863 566 23883
rect 588 23863 590 23883
rect 660 23863 662 23883
rect 708 23863 710 23883
rect 783 23880 797 23883
rect 807 23883 5237 23887
rect 807 23880 821 23883
rect 948 23863 950 23883
rect 1044 23863 1046 23883
rect 1092 23863 1094 23883
rect 1140 23863 1142 23883
rect 1308 23863 1310 23883
rect 1356 23863 1358 23883
rect 1572 23863 1574 23883
rect 1860 23863 1862 23883
rect 1956 23863 1958 23883
rect 2052 23863 2054 23883
rect 2148 23863 2150 23883
rect 2244 23863 2246 23883
rect 2340 23863 2342 23883
rect 2436 23863 2438 23883
rect 2532 23863 2534 23883
rect 2628 23863 2630 23883
rect 2724 23863 2726 23883
rect 2940 23863 2942 23883
rect 2988 23863 2990 23883
rect 3324 23863 3326 23883
rect 3540 23863 3542 23883
rect 3780 23863 3782 23883
rect 4068 23863 4070 23883
rect 4308 23863 4310 23883
rect 4932 23863 4934 23883
rect 4980 23863 4982 23883
rect 5028 23863 5030 23883
rect 5124 23863 5126 23883
rect 5148 23863 5150 23883
rect 5220 23863 5222 23883
rect 5223 23880 5237 23883
rect 5244 23883 11501 23887
rect 5244 23880 5261 23883
rect 5244 23863 5246 23880
rect 5460 23863 5462 23883
rect 5508 23863 5510 23883
rect 5556 23863 5558 23883
rect 5652 23863 5654 23883
rect 5748 23863 5750 23883
rect 5796 23863 5798 23883
rect 5844 23863 5846 23883
rect 5892 23863 5894 23883
rect 6276 23863 6278 23883
rect 6300 23863 6302 23883
rect 6372 23863 6374 23883
rect 6396 23863 6398 23883
rect 6492 23863 6494 23883
rect 6516 23863 6518 23883
rect 6588 23863 6590 23883
rect 6612 23863 6614 23883
rect 6636 23863 6638 23883
rect 6708 23863 6710 23883
rect 6804 23863 6806 23883
rect 6900 23863 6902 23883
rect 7164 23863 7166 23883
rect 7284 23863 7286 23883
rect 7380 23863 7382 23883
rect 7404 23863 7406 23883
rect 7476 23863 7478 23883
rect 7500 23863 7502 23883
rect 7572 23863 7574 23883
rect 7596 23863 7598 23883
rect 7668 23863 7670 23883
rect 7692 23863 7694 23883
rect 7908 23863 7910 23883
rect 8124 23863 8126 23883
rect 8220 23863 8222 23883
rect 8316 23863 8318 23883
rect 8412 23863 8414 23883
rect 8700 23863 8702 23883
rect 8748 23863 8750 23883
rect 8796 23863 8798 23883
rect 8844 23863 8846 23883
rect 8868 23863 8870 23883
rect 9516 23863 9518 23883
rect 9660 23880 9662 23883
rect 9660 23863 9663 23880
rect 9684 23863 9686 23883
rect 9780 23863 9782 23883
rect 9804 23863 9806 23883
rect 9828 23863 9830 23883
rect 10044 23863 10046 23883
rect 10140 23863 10142 23883
rect 10236 23863 10238 23883
rect 10332 23863 10334 23883
rect 10380 23863 10382 23883
rect 10428 23863 10430 23883
rect 10524 23863 10526 23883
rect 10548 23863 10550 23883
rect 10620 23863 10622 23883
rect 10644 23863 10646 23883
rect 10716 23863 10718 23883
rect 10860 23863 10862 23883
rect 10956 23863 10958 23883
rect 11052 23863 11054 23883
rect 11100 23863 11102 23883
rect 11172 23863 11174 23883
rect 11220 23863 11222 23883
rect 11340 23863 11342 23883
rect 11487 23880 11501 23883
rect 11508 23883 20075 23887
rect 11508 23880 11525 23883
rect 11508 23863 11510 23880
rect 11676 23863 11678 23883
rect 11724 23863 11726 23883
rect 11796 23863 11798 23883
rect 12060 23863 12062 23883
rect 12276 23863 12278 23883
rect 12372 23863 12374 23883
rect 12468 23863 12470 23883
rect 12564 23863 12566 23883
rect 12780 23863 12782 23883
rect 12876 23863 12878 23883
rect 13044 23863 13046 23883
rect 13164 23863 13166 23883
rect 13260 23863 13262 23883
rect 13332 23863 13334 23883
rect 13356 23863 13358 23883
rect 13500 23863 13502 23883
rect 13572 23863 13574 23883
rect 13836 23863 13838 23883
rect 13932 23863 13934 23883
rect 14004 23863 14006 23883
rect 14028 23863 14030 23883
rect 14172 23863 14174 23883
rect 14940 23863 14942 23883
rect 15036 23863 15038 23883
rect 15276 23863 15278 23883
rect 15372 23863 15374 23883
rect 15409 23878 15412 23883
rect 15420 23878 15422 23883
rect 15419 23864 15422 23878
rect 15468 23863 15470 23883
rect 15564 23863 15566 23883
rect 15660 23863 15662 23883
rect 15684 23863 15686 23883
rect 15732 23863 15734 23883
rect 15756 23863 15758 23883
rect 15780 23863 15782 23883
rect 15828 23863 15830 23883
rect 15852 23863 15854 23883
rect 15876 23863 15878 23883
rect 15948 23863 15950 23883
rect 15972 23863 15974 23883
rect 16044 23863 16046 23883
rect 16068 23863 16070 23883
rect 16164 23863 16166 23883
rect 16260 23863 16262 23883
rect 16284 23863 16286 23883
rect 16380 23863 16382 23883
rect 16476 23863 16478 23883
rect 16548 23863 16550 23883
rect 16596 23863 16598 23883
rect 16647 23880 16661 23883
rect 16668 23880 16671 23883
rect 16692 23863 16694 23883
rect 16764 23863 16766 23883
rect 16788 23863 16790 23883
rect 16884 23863 16886 23883
rect 16908 23863 16910 23883
rect 17028 23863 17030 23883
rect 17124 23863 17126 23883
rect 17196 23863 17198 23883
rect 17220 23863 17222 23883
rect 17292 23863 17294 23883
rect 17316 23863 17318 23883
rect 17964 23863 17966 23883
rect 18060 23863 18062 23883
rect 18132 23863 18134 23883
rect 18228 23863 18230 23883
rect 18492 23863 18494 23883
rect 18540 23863 18542 23883
rect 18636 23863 18638 23883
rect 18732 23863 18734 23883
rect 18828 23863 18830 23883
rect 18924 23863 18926 23883
rect 18972 23863 18974 23883
rect 19020 23863 19022 23883
rect 19068 23863 19070 23883
rect 19140 23863 19142 23883
rect 19164 23863 19166 23883
rect 19236 23863 19238 23883
rect 19260 23863 19262 23883
rect 19788 23864 19790 23883
rect 19836 23864 19838 23883
rect 19873 23878 19876 23883
rect 19884 23878 19886 23883
rect 19935 23880 19949 23883
rect 19969 23878 19972 23883
rect 19980 23880 19982 23883
rect 19980 23878 19983 23880
rect 19883 23864 19886 23878
rect 19979 23870 19983 23878
rect 19993 23878 19996 23883
rect 20004 23880 20006 23883
rect 20004 23878 20007 23880
rect 19993 23870 19997 23878
rect 19979 23864 19993 23870
rect 20003 23864 20007 23878
rect 20065 23870 20069 23878
rect 20055 23864 20065 23870
rect 19753 23863 19811 23864
rect 19825 23863 19859 23864
rect -2783 23859 19859 23863
rect -3551 23854 -3548 23859
rect -3540 23856 -3538 23859
rect -3540 23854 -3537 23856
rect -3479 23854 -3476 23859
rect -3468 23856 -3466 23859
rect -3468 23854 -3465 23856
rect -3551 23846 -3547 23854
rect -3561 23840 -3551 23846
rect -3541 23840 -3537 23854
rect -3469 23846 -3465 23854
rect -3455 23854 -3452 23859
rect -3444 23856 -3442 23859
rect -3444 23854 -3441 23856
rect -3119 23854 -3116 23859
rect -3108 23854 -3106 23859
rect -3023 23854 -3020 23859
rect -3012 23856 -3010 23859
rect -2783 23856 -2779 23859
rect -2772 23856 -2769 23859
rect -3012 23854 -3009 23856
rect -3455 23846 -3451 23854
rect -3469 23840 -3455 23846
rect -3445 23840 -3441 23854
rect -3109 23840 -3106 23854
rect -3013 23846 -3009 23854
rect -2999 23846 -2995 23854
rect -3013 23840 -2999 23846
rect -2364 23840 -2362 23859
rect -3335 23839 -3301 23840
rect -3263 23839 -3229 23840
rect -3335 23835 -3229 23839
rect -3215 23839 -3181 23840
rect -3143 23839 -3109 23840
rect -3215 23835 -3109 23839
rect -2663 23839 -2629 23840
rect -2471 23839 -2413 23840
rect -2375 23839 -2341 23840
rect -2663 23835 -2341 23839
rect -2327 23839 -2293 23840
rect -2063 23839 -2029 23840
rect -2327 23835 -2029 23839
rect -2015 23839 -1981 23840
rect -1908 23839 -1906 23859
rect -1452 23839 -1450 23859
rect -1356 23839 -1354 23859
rect -1332 23839 -1330 23859
rect -1260 23839 -1258 23859
rect -1236 23839 -1234 23859
rect -1140 23839 -1138 23859
rect -876 23839 -874 23859
rect -780 23839 -778 23859
rect -564 23839 -562 23859
rect -468 23839 -466 23859
rect -12 23839 -10 23859
rect 84 23839 86 23859
rect 180 23839 182 23859
rect 468 23839 470 23859
rect 492 23839 494 23859
rect 564 23839 566 23859
rect 588 23839 590 23859
rect 660 23839 662 23859
rect 708 23839 710 23859
rect 948 23839 950 23859
rect 1044 23839 1046 23859
rect 1092 23839 1094 23859
rect 1140 23839 1142 23859
rect 1308 23839 1310 23859
rect 1356 23839 1358 23859
rect 1572 23839 1574 23859
rect 1860 23839 1862 23859
rect 1956 23839 1958 23859
rect 2052 23839 2054 23859
rect 2148 23839 2150 23859
rect 2244 23839 2246 23859
rect 2340 23839 2342 23859
rect 2436 23839 2438 23859
rect 2532 23839 2534 23859
rect 2628 23839 2630 23859
rect 2724 23839 2726 23859
rect 2940 23839 2942 23859
rect 2988 23839 2990 23859
rect 3255 23856 3269 23859
rect 3324 23839 3326 23859
rect 3540 23839 3542 23859
rect 3780 23839 3782 23859
rect 3807 23856 3821 23859
rect 4068 23839 4070 23859
rect 4308 23839 4310 23859
rect 4932 23839 4934 23859
rect 4980 23839 4982 23859
rect 5028 23839 5030 23859
rect 5124 23839 5126 23859
rect 5148 23839 5150 23859
rect 5220 23839 5222 23859
rect 5244 23839 5246 23859
rect 5460 23839 5462 23859
rect 5508 23839 5510 23859
rect 5556 23839 5558 23859
rect 5652 23839 5654 23859
rect 5748 23839 5750 23859
rect 5796 23839 5798 23859
rect 5844 23839 5846 23859
rect 5892 23839 5894 23859
rect 6276 23839 6278 23859
rect 6300 23839 6302 23859
rect 6372 23839 6374 23859
rect 6396 23839 6398 23859
rect 6492 23839 6494 23859
rect 6516 23839 6518 23859
rect 6588 23839 6590 23859
rect 6612 23839 6614 23859
rect 6636 23839 6638 23859
rect 6708 23839 6710 23859
rect 6804 23839 6806 23859
rect 6900 23839 6902 23859
rect 7164 23839 7166 23859
rect 7284 23839 7286 23859
rect 7311 23856 7325 23859
rect 7380 23839 7382 23859
rect 7404 23839 7406 23859
rect 7476 23839 7478 23859
rect 7500 23839 7502 23859
rect 7572 23839 7574 23859
rect 7596 23839 7598 23859
rect 7668 23839 7670 23859
rect 7692 23839 7694 23859
rect 7908 23839 7910 23859
rect 8124 23839 8126 23859
rect 8220 23839 8222 23859
rect 8316 23839 8318 23859
rect 8412 23839 8414 23859
rect 8700 23839 8702 23859
rect 8748 23839 8750 23859
rect 8796 23839 8798 23859
rect 8844 23839 8846 23859
rect 8868 23839 8870 23859
rect 9516 23839 9518 23859
rect 9639 23856 9653 23859
rect 9660 23856 9663 23859
rect 9684 23839 9686 23859
rect 9780 23839 9782 23859
rect 9804 23839 9806 23859
rect 9828 23839 9830 23859
rect 10044 23839 10046 23859
rect 10140 23839 10142 23859
rect 10236 23839 10238 23859
rect 10332 23839 10334 23859
rect 10380 23839 10382 23859
rect 10428 23839 10430 23859
rect 10524 23839 10526 23859
rect 10548 23839 10550 23859
rect 10620 23839 10622 23859
rect 10644 23839 10646 23859
rect 10716 23839 10718 23859
rect 10860 23839 10862 23859
rect 10956 23839 10958 23859
rect 11052 23839 11054 23859
rect 11100 23839 11102 23859
rect 11172 23839 11174 23859
rect 11220 23839 11222 23859
rect 11340 23839 11342 23859
rect 11508 23839 11510 23859
rect 11676 23839 11678 23859
rect 11724 23839 11726 23859
rect 11796 23839 11798 23859
rect 12060 23839 12062 23859
rect 12276 23839 12278 23859
rect 12372 23839 12374 23859
rect 12468 23839 12470 23859
rect 12564 23839 12566 23859
rect 12780 23839 12782 23859
rect 12876 23839 12878 23859
rect 13044 23839 13046 23859
rect 13164 23839 13166 23859
rect 13260 23839 13262 23859
rect 13332 23839 13334 23859
rect 13356 23839 13358 23859
rect 13500 23839 13502 23859
rect 13572 23839 13574 23859
rect 13836 23839 13838 23859
rect 13932 23839 13934 23859
rect 14004 23839 14006 23859
rect 14028 23839 14030 23859
rect 14172 23839 14174 23859
rect 14940 23839 14942 23859
rect 15036 23839 15038 23859
rect 15276 23839 15278 23859
rect 15372 23839 15374 23859
rect 15468 23839 15470 23859
rect 15495 23856 15509 23859
rect 15564 23839 15566 23859
rect 15660 23839 15662 23859
rect 15684 23839 15686 23859
rect 15732 23839 15734 23859
rect 15756 23839 15758 23859
rect 15780 23839 15782 23859
rect 15828 23839 15830 23859
rect 15852 23839 15854 23859
rect 15876 23839 15878 23859
rect 15948 23839 15950 23859
rect 15972 23839 15974 23859
rect 16044 23839 16046 23859
rect 16068 23839 16070 23859
rect 16164 23839 16166 23859
rect 16260 23839 16262 23859
rect 16284 23839 16286 23859
rect 16380 23839 16382 23859
rect 16476 23839 16478 23859
rect 16548 23839 16550 23859
rect 16596 23839 16598 23859
rect 16692 23839 16694 23859
rect 16764 23839 16766 23859
rect 16788 23839 16790 23859
rect 16884 23839 16886 23859
rect 16908 23839 16910 23859
rect 17028 23839 17030 23859
rect 17124 23839 17126 23859
rect 17196 23839 17198 23859
rect 17220 23839 17222 23859
rect 17292 23839 17294 23859
rect 17316 23839 17318 23859
rect 17964 23839 17966 23859
rect 18060 23839 18062 23859
rect 18132 23839 18134 23859
rect 18228 23839 18230 23859
rect 18492 23839 18494 23859
rect 18540 23839 18542 23859
rect 18636 23839 18638 23859
rect 18732 23839 18734 23859
rect 18828 23839 18830 23859
rect 18924 23839 18926 23859
rect 18972 23839 18974 23859
rect 19020 23839 19022 23859
rect 19068 23839 19070 23859
rect 19140 23839 19142 23859
rect 19164 23839 19166 23859
rect 19236 23839 19238 23859
rect 19260 23839 19262 23859
rect 19777 23854 19780 23859
rect 19788 23854 19790 23859
rect 19825 23854 19828 23859
rect 19836 23854 19838 23859
rect 19787 23840 19790 23854
rect 19835 23840 19838 23854
rect 19849 23846 19853 23854
rect 19839 23840 19849 23846
rect 19729 23839 19763 23840
rect -2015 23835 19763 23839
rect -2375 23830 -2372 23835
rect -2364 23832 -2362 23835
rect -1908 23832 -1906 23835
rect -2364 23830 -2361 23832
rect -3239 23822 -3235 23830
rect -3119 23822 -3115 23830
rect -2365 23822 -2361 23830
rect -2351 23822 -2347 23830
rect -3249 23816 -3239 23822
rect -3129 23816 -3119 23822
rect -2365 23816 -2351 23822
rect -1908 23816 -1905 23832
rect -2135 23815 -2101 23816
rect -2087 23815 -2053 23816
rect -2135 23811 -2053 23815
rect -1919 23815 -1885 23816
rect -1703 23815 -1645 23816
rect -1452 23815 -1450 23835
rect -1356 23815 -1354 23835
rect -1332 23815 -1330 23835
rect -1260 23815 -1258 23835
rect -1236 23815 -1234 23835
rect -1140 23816 -1138 23835
rect -1151 23815 -1117 23816
rect -1919 23811 -1117 23815
rect -1103 23815 -1069 23816
rect -876 23815 -874 23835
rect -780 23815 -778 23835
rect -564 23815 -562 23835
rect -468 23815 -466 23835
rect -407 23815 -373 23816
rect -143 23815 -85 23816
rect -12 23815 -10 23835
rect 84 23815 86 23835
rect 180 23815 182 23835
rect 468 23815 470 23835
rect 492 23815 494 23835
rect 564 23815 566 23835
rect 588 23815 590 23835
rect 660 23815 662 23835
rect 708 23815 710 23835
rect 948 23815 950 23835
rect 1044 23815 1046 23835
rect 1092 23815 1094 23835
rect 1140 23815 1142 23835
rect 1308 23815 1310 23835
rect 1356 23815 1358 23835
rect 1572 23815 1574 23835
rect 1860 23815 1862 23835
rect 1956 23815 1958 23835
rect 2052 23815 2054 23835
rect 2148 23815 2150 23835
rect 2244 23815 2246 23835
rect 2340 23815 2342 23835
rect 2436 23815 2438 23835
rect 2532 23815 2534 23835
rect 2628 23815 2630 23835
rect 2724 23815 2726 23835
rect 2940 23815 2942 23835
rect 2988 23815 2990 23835
rect 3324 23815 3326 23835
rect 3540 23815 3542 23835
rect 3780 23815 3782 23835
rect 4068 23815 4070 23835
rect 4308 23815 4310 23835
rect 4932 23815 4934 23835
rect 4980 23815 4982 23835
rect 5028 23815 5030 23835
rect 5124 23815 5126 23835
rect 5148 23815 5150 23835
rect 5220 23815 5222 23835
rect 5244 23815 5246 23835
rect 5460 23815 5462 23835
rect 5508 23815 5510 23835
rect 5556 23815 5558 23835
rect 5652 23815 5654 23835
rect 5665 23815 5723 23816
rect 5748 23815 5750 23835
rect 5796 23815 5798 23835
rect 5844 23815 5846 23835
rect 5892 23815 5894 23835
rect 6276 23815 6278 23835
rect 6300 23815 6302 23835
rect 6372 23815 6374 23835
rect 6396 23815 6398 23835
rect 6492 23815 6494 23835
rect 6516 23815 6518 23835
rect 6588 23815 6590 23835
rect 6612 23815 6614 23835
rect 6636 23815 6638 23835
rect 6708 23815 6710 23835
rect 6804 23815 6806 23835
rect 6900 23815 6902 23835
rect 7164 23815 7166 23835
rect 7284 23815 7286 23835
rect 7380 23815 7382 23835
rect 7404 23815 7406 23835
rect 7476 23815 7478 23835
rect 7500 23815 7502 23835
rect 7572 23815 7574 23835
rect 7596 23815 7598 23835
rect 7668 23815 7670 23835
rect 7692 23815 7694 23835
rect 7908 23815 7910 23835
rect 8124 23815 8126 23835
rect 8220 23815 8222 23835
rect 8316 23815 8318 23835
rect 8412 23815 8414 23835
rect 8700 23815 8702 23835
rect 8748 23815 8750 23835
rect 8796 23815 8798 23835
rect 8844 23815 8846 23835
rect 8868 23815 8870 23835
rect 9516 23815 9518 23835
rect 9684 23815 9686 23835
rect 9780 23815 9782 23835
rect 9804 23815 9806 23835
rect 9828 23815 9830 23835
rect 10044 23815 10046 23835
rect 10140 23815 10142 23835
rect 10236 23815 10238 23835
rect 10332 23815 10334 23835
rect 10380 23815 10382 23835
rect 10428 23815 10430 23835
rect 10524 23815 10526 23835
rect 10548 23815 10550 23835
rect 10620 23815 10622 23835
rect 10644 23815 10646 23835
rect 10716 23815 10718 23835
rect 10860 23815 10862 23835
rect 10956 23815 10958 23835
rect 11052 23815 11054 23835
rect 11100 23815 11102 23835
rect 11172 23816 11174 23835
rect 11137 23815 11195 23816
rect 11220 23815 11222 23835
rect 11340 23815 11342 23835
rect 11508 23815 11510 23835
rect 11676 23815 11678 23835
rect 11724 23815 11726 23835
rect 11796 23815 11798 23835
rect 12060 23815 12062 23835
rect 12276 23815 12278 23835
rect 12372 23815 12374 23835
rect 12468 23815 12470 23835
rect 12564 23815 12566 23835
rect 12780 23815 12782 23835
rect 12876 23815 12878 23835
rect 13044 23815 13046 23835
rect 13164 23815 13166 23835
rect 13260 23815 13262 23835
rect 13332 23815 13334 23835
rect 13356 23815 13358 23835
rect 13500 23815 13502 23835
rect 13572 23815 13574 23835
rect 13836 23815 13838 23835
rect 13932 23815 13934 23835
rect 14004 23815 14006 23835
rect 14028 23815 14030 23835
rect 14172 23815 14174 23835
rect 14940 23815 14942 23835
rect 15036 23815 15038 23835
rect 15276 23815 15278 23835
rect 15372 23815 15374 23835
rect 15468 23815 15470 23835
rect 15564 23815 15566 23835
rect 15660 23815 15662 23835
rect 15684 23815 15686 23835
rect 15732 23815 15734 23835
rect 15756 23815 15758 23835
rect 15780 23815 15782 23835
rect 15828 23815 15830 23835
rect 15852 23815 15854 23835
rect 15876 23815 15878 23835
rect 15948 23815 15950 23835
rect 15972 23815 15974 23835
rect 16044 23815 16046 23835
rect 16068 23815 16070 23835
rect 16164 23815 16166 23835
rect 16260 23815 16262 23835
rect 16284 23815 16286 23835
rect 16380 23815 16382 23835
rect 16476 23815 16478 23835
rect 16548 23815 16550 23835
rect 16596 23815 16598 23835
rect 16692 23815 16694 23835
rect 16764 23815 16766 23835
rect 16788 23815 16790 23835
rect 16884 23815 16886 23835
rect 16908 23815 16910 23835
rect 17028 23815 17030 23835
rect 17124 23815 17126 23835
rect 17196 23815 17198 23835
rect 17220 23815 17222 23835
rect 17292 23815 17294 23835
rect 17316 23815 17318 23835
rect 17964 23815 17966 23835
rect 18060 23815 18062 23835
rect 18132 23815 18134 23835
rect 18228 23815 18230 23835
rect 18492 23815 18494 23835
rect 18540 23815 18542 23835
rect 18636 23815 18638 23835
rect 18732 23815 18734 23835
rect 18828 23815 18830 23835
rect 18924 23815 18926 23835
rect 18972 23815 18974 23835
rect 19020 23815 19022 23835
rect 19068 23815 19070 23835
rect 19140 23815 19142 23835
rect 19164 23815 19166 23835
rect 19236 23815 19238 23835
rect 19260 23815 19262 23835
rect 19705 23815 19739 23816
rect -1103 23811 19739 23815
rect -1919 23808 -1915 23811
rect -1908 23808 -1905 23811
rect -1452 23792 -1450 23811
rect -1559 23791 -1525 23792
rect -1463 23791 -1429 23792
rect -1356 23791 -1354 23811
rect -1332 23791 -1330 23811
rect -1260 23791 -1258 23811
rect -1236 23792 -1234 23811
rect -1151 23806 -1148 23811
rect -1140 23806 -1138 23811
rect -1141 23792 -1138 23806
rect -1247 23791 -1213 23792
rect -1559 23787 -1213 23791
rect -983 23791 -949 23792
rect -876 23791 -874 23811
rect -780 23791 -778 23811
rect -564 23791 -562 23811
rect -468 23791 -466 23811
rect -143 23806 -140 23811
rect -12 23808 -10 23811
rect -133 23792 -130 23806
rect -132 23791 -130 23792
rect -12 23791 -9 23808
rect 84 23791 86 23811
rect 180 23791 182 23811
rect 468 23791 470 23811
rect 492 23791 494 23811
rect 564 23791 566 23811
rect 588 23791 590 23811
rect 660 23791 662 23811
rect 708 23791 710 23811
rect 948 23791 950 23811
rect 1044 23791 1046 23811
rect 1092 23791 1094 23811
rect 1140 23791 1142 23811
rect 1308 23791 1310 23811
rect 1356 23791 1358 23811
rect 1572 23791 1574 23811
rect 1860 23791 1862 23811
rect 1956 23791 1958 23811
rect 2052 23791 2054 23811
rect 2148 23791 2150 23811
rect 2244 23791 2246 23811
rect 2340 23791 2342 23811
rect 2436 23791 2438 23811
rect 2532 23791 2534 23811
rect 2628 23791 2630 23811
rect 2724 23791 2726 23811
rect 2940 23791 2942 23811
rect 2988 23791 2990 23811
rect 3324 23791 3326 23811
rect 3540 23791 3542 23811
rect 3780 23791 3782 23811
rect 4068 23791 4070 23811
rect 4308 23791 4310 23811
rect 4932 23791 4934 23811
rect 4980 23791 4982 23811
rect 5028 23791 5030 23811
rect 5124 23791 5126 23811
rect 5148 23791 5150 23811
rect 5220 23791 5222 23811
rect 5244 23791 5246 23811
rect 5460 23791 5462 23811
rect 5508 23791 5510 23811
rect 5556 23791 5558 23811
rect 5652 23791 5654 23811
rect 5748 23791 5750 23811
rect 5796 23808 5798 23811
rect 5796 23791 5799 23808
rect 5844 23791 5846 23811
rect 5892 23791 5894 23811
rect 6276 23791 6278 23811
rect 6300 23791 6302 23811
rect 6372 23791 6374 23811
rect 6396 23791 6398 23811
rect 6492 23791 6494 23811
rect 6516 23791 6518 23811
rect 6588 23791 6590 23811
rect 6612 23791 6614 23811
rect 6636 23791 6638 23811
rect 6708 23791 6710 23811
rect 6804 23791 6806 23811
rect 6900 23791 6902 23811
rect 7164 23791 7166 23811
rect 7284 23791 7286 23811
rect 7380 23791 7382 23811
rect 7404 23791 7406 23811
rect 7476 23791 7478 23811
rect 7500 23791 7502 23811
rect 7572 23791 7574 23811
rect 7596 23791 7598 23811
rect 7668 23791 7670 23811
rect 7692 23791 7694 23811
rect 7908 23791 7910 23811
rect 8124 23791 8126 23811
rect 8220 23791 8222 23811
rect 8316 23791 8318 23811
rect 8412 23791 8414 23811
rect 8700 23791 8702 23811
rect 8748 23791 8750 23811
rect 8796 23791 8798 23811
rect 8844 23791 8846 23811
rect 8868 23791 8870 23811
rect 9516 23791 9518 23811
rect 9684 23791 9686 23811
rect 9780 23791 9782 23811
rect 9804 23791 9806 23811
rect 9828 23791 9830 23811
rect 10044 23791 10046 23811
rect 10140 23791 10142 23811
rect 10236 23791 10238 23811
rect 10332 23791 10334 23811
rect 10380 23791 10382 23811
rect 10428 23791 10430 23811
rect 10524 23791 10526 23811
rect 10548 23791 10550 23811
rect 10620 23791 10622 23811
rect 10644 23791 10646 23811
rect 10716 23791 10718 23811
rect 10860 23791 10862 23811
rect 10956 23791 10958 23811
rect 11052 23791 11054 23811
rect 11100 23791 11102 23811
rect 11137 23806 11140 23811
rect 11161 23806 11164 23811
rect 11172 23806 11174 23811
rect 11147 23792 11150 23806
rect 11171 23792 11174 23806
rect 11148 23791 11150 23792
rect 11220 23791 11222 23811
rect 11244 23791 11247 23808
rect 11340 23791 11342 23811
rect 11508 23791 11510 23811
rect 11676 23791 11678 23811
rect 11724 23791 11726 23811
rect 11796 23791 11798 23811
rect 12060 23791 12062 23811
rect 12276 23791 12278 23811
rect 12372 23791 12374 23811
rect 12468 23791 12470 23811
rect 12564 23791 12566 23811
rect 12780 23791 12782 23811
rect 12876 23791 12878 23811
rect 13044 23791 13046 23811
rect 13164 23791 13166 23811
rect 13260 23791 13262 23811
rect 13332 23791 13334 23811
rect 13356 23791 13358 23811
rect 13500 23791 13502 23811
rect 13572 23791 13574 23811
rect 13836 23791 13838 23811
rect 13932 23791 13934 23811
rect 14004 23791 14006 23811
rect 14028 23791 14030 23811
rect 14172 23791 14174 23811
rect 14473 23791 14507 23792
rect 14940 23791 14942 23811
rect 15036 23791 15038 23811
rect 15276 23791 15278 23811
rect 15372 23791 15374 23811
rect 15468 23791 15470 23811
rect 15564 23791 15566 23811
rect 15660 23791 15662 23811
rect 15684 23791 15686 23811
rect 15732 23791 15734 23811
rect 15756 23791 15758 23811
rect 15780 23791 15782 23811
rect 15828 23791 15830 23811
rect 15852 23791 15854 23811
rect 15876 23791 15878 23811
rect 15948 23791 15950 23811
rect 15972 23791 15974 23811
rect 16044 23791 16046 23811
rect 16068 23791 16070 23811
rect 16164 23791 16166 23811
rect 16260 23791 16262 23811
rect 16284 23791 16286 23811
rect 16380 23791 16382 23811
rect 16476 23791 16478 23811
rect 16548 23791 16550 23811
rect 16596 23791 16598 23811
rect 16692 23791 16694 23811
rect 16764 23791 16766 23811
rect 16788 23791 16790 23811
rect 16884 23791 16886 23811
rect 16908 23791 16910 23811
rect 17028 23791 17030 23811
rect 17124 23791 17126 23811
rect 17196 23791 17198 23811
rect 17220 23791 17222 23811
rect 17292 23791 17294 23811
rect 17316 23791 17318 23811
rect 17964 23791 17966 23811
rect 18060 23791 18062 23811
rect 18132 23791 18134 23811
rect 18228 23791 18230 23811
rect 18492 23791 18494 23811
rect 18540 23791 18542 23811
rect 18636 23791 18638 23811
rect 18732 23791 18734 23811
rect 18828 23791 18830 23811
rect 18924 23791 18926 23811
rect 18972 23791 18974 23811
rect 19020 23792 19022 23811
rect 19009 23791 19043 23792
rect 19068 23791 19070 23811
rect 19140 23791 19142 23811
rect 19164 23791 19166 23811
rect 19236 23791 19238 23811
rect 19260 23791 19262 23811
rect 19681 23791 19715 23792
rect -983 23787 -43 23791
rect -1463 23782 -1460 23787
rect -1452 23784 -1450 23787
rect -1356 23784 -1354 23787
rect -1452 23782 -1449 23784
rect -1453 23768 -1449 23782
rect -1356 23768 -1353 23784
rect -1332 23768 -1330 23787
rect -1260 23768 -1258 23787
rect -1247 23782 -1244 23787
rect -1236 23782 -1234 23787
rect -1237 23768 -1234 23782
rect -876 23784 -874 23787
rect -876 23768 -873 23784
rect -780 23768 -778 23787
rect -1439 23767 -1405 23768
rect -1367 23767 -1309 23768
rect -1271 23767 -1237 23768
rect -1439 23763 -1237 23767
rect -887 23767 -853 23768
rect -839 23767 -805 23768
rect -887 23763 -805 23767
rect -791 23767 -757 23768
rect -564 23767 -562 23787
rect -468 23767 -466 23787
rect -321 23784 -307 23787
rect -132 23767 -130 23787
rect -57 23784 -43 23787
rect -33 23787 5765 23791
rect -33 23784 -19 23787
rect -12 23784 -9 23787
rect 84 23767 86 23787
rect 180 23767 182 23787
rect 468 23767 470 23787
rect 492 23767 494 23787
rect 564 23767 566 23787
rect 588 23767 590 23787
rect 660 23767 662 23787
rect 708 23767 710 23787
rect 948 23767 950 23787
rect 1044 23767 1046 23787
rect 1092 23767 1094 23787
rect 1140 23767 1142 23787
rect 1308 23767 1310 23787
rect 1356 23767 1358 23787
rect 1572 23767 1574 23787
rect 1860 23767 1862 23787
rect 1956 23767 1958 23787
rect 2052 23767 2054 23787
rect 2148 23767 2150 23787
rect 2244 23767 2246 23787
rect 2340 23767 2342 23787
rect 2436 23767 2438 23787
rect 2532 23767 2534 23787
rect 2628 23767 2630 23787
rect 2724 23767 2726 23787
rect 2940 23767 2942 23787
rect 2988 23767 2990 23787
rect 3324 23767 3326 23787
rect 3540 23767 3542 23787
rect 3780 23767 3782 23787
rect 4068 23767 4070 23787
rect 4153 23767 4211 23768
rect 4308 23767 4310 23787
rect 4932 23767 4934 23787
rect 4980 23767 4982 23787
rect 5028 23767 5030 23787
rect 5124 23767 5126 23787
rect 5148 23767 5150 23787
rect 5220 23767 5222 23787
rect 5244 23767 5246 23787
rect 5460 23767 5462 23787
rect 5508 23767 5510 23787
rect 5556 23767 5558 23787
rect 5652 23767 5654 23787
rect 5748 23767 5750 23787
rect 5751 23784 5765 23787
rect 5775 23787 11237 23791
rect 5775 23784 5789 23787
rect 5796 23784 5799 23787
rect 5844 23767 5846 23787
rect 5892 23767 5894 23787
rect 6276 23767 6278 23787
rect 6300 23767 6302 23787
rect 6372 23767 6374 23787
rect 6396 23767 6398 23787
rect 6492 23767 6494 23787
rect 6516 23767 6518 23787
rect 6588 23767 6590 23787
rect 6612 23767 6614 23787
rect 6636 23767 6638 23787
rect 6708 23767 6710 23787
rect 6804 23767 6806 23787
rect 6900 23767 6902 23787
rect 7164 23767 7166 23787
rect 7284 23767 7286 23787
rect 7380 23767 7382 23787
rect 7404 23767 7406 23787
rect 7476 23767 7478 23787
rect 7500 23767 7502 23787
rect 7572 23767 7574 23787
rect 7596 23767 7598 23787
rect 7668 23767 7670 23787
rect 7692 23767 7694 23787
rect 7908 23767 7910 23787
rect 8124 23767 8126 23787
rect 8220 23767 8222 23787
rect 8316 23767 8318 23787
rect 8412 23767 8414 23787
rect 8700 23767 8702 23787
rect 8748 23767 8750 23787
rect 8796 23767 8798 23787
rect 8844 23767 8846 23787
rect 8868 23767 8870 23787
rect 9516 23767 9518 23787
rect 9684 23767 9686 23787
rect 9780 23767 9782 23787
rect 9804 23767 9806 23787
rect 9828 23767 9830 23787
rect 10044 23767 10046 23787
rect 10140 23767 10142 23787
rect 10236 23767 10238 23787
rect 10332 23767 10334 23787
rect 10380 23767 10382 23787
rect 10428 23767 10430 23787
rect 10524 23767 10526 23787
rect 10548 23767 10550 23787
rect 10620 23767 10622 23787
rect 10644 23767 10646 23787
rect 10716 23767 10718 23787
rect 10860 23767 10862 23787
rect 10956 23767 10958 23787
rect 11052 23767 11054 23787
rect 11100 23767 11102 23787
rect 11148 23767 11150 23787
rect 11220 23767 11222 23787
rect 11223 23784 11237 23787
rect 11244 23787 19715 23791
rect 11244 23784 11261 23787
rect 11244 23767 11246 23784
rect 11257 23767 11315 23768
rect 11340 23767 11342 23787
rect 11508 23767 11510 23787
rect 11676 23767 11678 23787
rect 11724 23767 11726 23787
rect 11796 23767 11798 23787
rect 12060 23767 12062 23787
rect 12276 23767 12278 23787
rect 12372 23767 12374 23787
rect 12468 23767 12470 23787
rect 12564 23767 12566 23787
rect 12780 23767 12782 23787
rect 12876 23767 12878 23787
rect 13044 23767 13046 23787
rect 13164 23767 13166 23787
rect 13260 23767 13262 23787
rect 13332 23767 13334 23787
rect 13356 23767 13358 23787
rect 13500 23767 13502 23787
rect 13572 23767 13574 23787
rect 13836 23767 13838 23787
rect 13932 23767 13934 23787
rect 14004 23767 14006 23787
rect 14028 23767 14030 23787
rect 14172 23767 14174 23787
rect 14940 23767 14942 23787
rect 15036 23767 15038 23787
rect 15276 23767 15278 23787
rect 15372 23767 15374 23787
rect 15468 23767 15470 23787
rect 15564 23767 15566 23787
rect 15660 23767 15662 23787
rect 15684 23767 15686 23787
rect 15732 23767 15734 23787
rect 15756 23767 15758 23787
rect 15780 23767 15782 23787
rect 15828 23767 15830 23787
rect 15852 23767 15854 23787
rect 15876 23767 15878 23787
rect 15948 23767 15950 23787
rect 15972 23767 15974 23787
rect 16044 23767 16046 23787
rect 16068 23767 16070 23787
rect 16164 23767 16166 23787
rect 16260 23767 16262 23787
rect 16284 23767 16286 23787
rect 16380 23767 16382 23787
rect 16476 23767 16478 23787
rect 16548 23767 16550 23787
rect 16596 23767 16598 23787
rect 16692 23767 16694 23787
rect 16764 23767 16766 23787
rect 16788 23767 16790 23787
rect 16884 23767 16886 23787
rect 16908 23767 16910 23787
rect 17028 23767 17030 23787
rect 17124 23767 17126 23787
rect 17196 23767 17198 23787
rect 17220 23767 17222 23787
rect 17292 23767 17294 23787
rect 17316 23767 17318 23787
rect 17964 23767 17966 23787
rect 18060 23767 18062 23787
rect 18132 23767 18134 23787
rect 18228 23767 18230 23787
rect 18492 23767 18494 23787
rect 18540 23767 18542 23787
rect 18636 23767 18638 23787
rect 18732 23767 18734 23787
rect 18828 23767 18830 23787
rect 18924 23767 18926 23787
rect 18972 23767 18974 23787
rect 19009 23782 19012 23787
rect 19020 23782 19022 23787
rect 19019 23768 19022 23782
rect 19068 23767 19070 23787
rect 19140 23767 19142 23787
rect 19164 23767 19166 23787
rect 19236 23767 19238 23787
rect 19260 23767 19262 23787
rect 19513 23767 19547 23768
rect -791 23763 19547 23767
rect -1377 23760 -1363 23763
rect -1356 23760 -1353 23763
rect -1343 23758 -1340 23763
rect -1332 23760 -1330 23763
rect -1332 23758 -1329 23760
rect -1271 23758 -1268 23763
rect -1260 23760 -1258 23763
rect -887 23760 -883 23763
rect -876 23760 -873 23763
rect -1260 23758 -1257 23760
rect -791 23758 -788 23763
rect -780 23760 -778 23763
rect -780 23758 -777 23760
rect -1343 23750 -1339 23758
rect -1353 23744 -1343 23750
rect -1333 23744 -1329 23758
rect -1261 23750 -1257 23758
rect -1247 23750 -1243 23758
rect -1261 23744 -1247 23750
rect -781 23744 -777 23758
rect -564 23744 -562 23763
rect -671 23743 -637 23744
rect -599 23743 -541 23744
rect -468 23743 -466 23763
rect -132 23743 -130 23763
rect 84 23743 86 23763
rect 180 23743 182 23763
rect 468 23743 470 23763
rect 492 23743 494 23763
rect 564 23743 566 23763
rect 588 23743 590 23763
rect 660 23743 662 23763
rect 708 23743 710 23763
rect 948 23743 950 23763
rect 1044 23743 1046 23763
rect 1092 23743 1094 23763
rect 1140 23743 1142 23763
rect 1308 23743 1310 23763
rect 1356 23743 1358 23763
rect 1572 23743 1574 23763
rect 1860 23743 1862 23763
rect 1956 23743 1958 23763
rect 2052 23743 2054 23763
rect 2148 23743 2150 23763
rect 2244 23743 2246 23763
rect 2340 23743 2342 23763
rect 2436 23743 2438 23763
rect 2532 23743 2534 23763
rect 2628 23743 2630 23763
rect 2724 23743 2726 23763
rect 2940 23743 2942 23763
rect 2988 23743 2990 23763
rect 3324 23743 3326 23763
rect 3540 23743 3542 23763
rect 3780 23743 3782 23763
rect 4068 23743 4070 23763
rect 4153 23758 4156 23763
rect 4163 23744 4166 23758
rect 4164 23743 4166 23744
rect 4308 23743 4310 23763
rect 4932 23743 4934 23763
rect 4980 23743 4982 23763
rect 5028 23743 5030 23763
rect 5124 23743 5126 23763
rect 5148 23743 5150 23763
rect 5220 23743 5222 23763
rect 5244 23743 5246 23763
rect 5460 23743 5462 23763
rect 5508 23743 5510 23763
rect 5556 23743 5558 23763
rect 5617 23743 5651 23744
rect 5652 23743 5654 23763
rect 5748 23743 5750 23763
rect 5761 23743 5819 23744
rect 5844 23743 5846 23763
rect 5892 23743 5894 23763
rect 6276 23743 6278 23763
rect 6300 23743 6302 23763
rect 6372 23743 6374 23763
rect 6396 23743 6398 23763
rect 6492 23743 6494 23763
rect 6516 23743 6518 23763
rect 6588 23743 6590 23763
rect 6612 23743 6614 23763
rect 6636 23743 6638 23763
rect 6708 23743 6710 23763
rect 6804 23743 6806 23763
rect 6900 23743 6902 23763
rect 7164 23743 7166 23763
rect 7284 23743 7286 23763
rect 7380 23743 7382 23763
rect 7404 23743 7406 23763
rect 7476 23743 7478 23763
rect 7500 23743 7502 23763
rect 7572 23743 7574 23763
rect 7596 23743 7598 23763
rect 7668 23743 7670 23763
rect 7692 23743 7694 23763
rect 7908 23743 7910 23763
rect 8124 23743 8126 23763
rect 8220 23743 8222 23763
rect 8316 23743 8318 23763
rect 8412 23743 8414 23763
rect 8700 23743 8702 23763
rect 8748 23743 8750 23763
rect 8796 23743 8798 23763
rect 8844 23743 8846 23763
rect 8868 23743 8870 23763
rect 9516 23743 9518 23763
rect 9684 23743 9686 23763
rect 9780 23743 9782 23763
rect 9804 23743 9806 23763
rect 9828 23743 9830 23763
rect 10044 23743 10046 23763
rect 10140 23743 10142 23763
rect 10236 23743 10238 23763
rect 10332 23743 10334 23763
rect 10380 23744 10382 23763
rect 10345 23743 10403 23744
rect 10428 23743 10430 23763
rect 10524 23743 10526 23763
rect 10548 23743 10550 23763
rect 10620 23743 10622 23763
rect 10644 23743 10646 23763
rect 10716 23743 10718 23763
rect 10860 23743 10862 23763
rect 10956 23743 10958 23763
rect 11052 23743 11054 23763
rect 11100 23743 11102 23763
rect 11148 23743 11150 23763
rect 11220 23743 11222 23763
rect 11244 23743 11246 23763
rect 11340 23743 11342 23763
rect 11364 23743 11367 23760
rect 11508 23743 11510 23763
rect 11676 23743 11678 23763
rect 11724 23743 11726 23763
rect 11796 23743 11798 23763
rect 12060 23743 12062 23763
rect 12276 23743 12278 23763
rect 12372 23743 12374 23763
rect 12468 23743 12470 23763
rect 12564 23743 12566 23763
rect 12780 23743 12782 23763
rect 12876 23743 12878 23763
rect 13044 23743 13046 23763
rect 13164 23743 13166 23763
rect 13260 23743 13262 23763
rect 13332 23743 13334 23763
rect 13356 23743 13358 23763
rect 13500 23743 13502 23763
rect 13572 23743 13574 23763
rect 13836 23743 13838 23763
rect 13932 23743 13934 23763
rect 14004 23743 14006 23763
rect 14028 23743 14030 23763
rect 14172 23743 14174 23763
rect 14559 23760 14573 23763
rect 14940 23743 14942 23763
rect 15036 23743 15038 23763
rect 15276 23743 15278 23763
rect 15372 23743 15374 23763
rect 15468 23743 15470 23763
rect 15564 23743 15566 23763
rect 15660 23743 15662 23763
rect 15684 23743 15686 23763
rect 15732 23743 15734 23763
rect 15756 23743 15758 23763
rect 15780 23743 15782 23763
rect 15828 23743 15830 23763
rect 15852 23743 15854 23763
rect 15876 23743 15878 23763
rect 15948 23743 15950 23763
rect 15972 23743 15974 23763
rect 16044 23743 16046 23763
rect 16068 23743 16070 23763
rect 16164 23743 16166 23763
rect 16260 23743 16262 23763
rect 16284 23743 16286 23763
rect 16380 23743 16382 23763
rect 16476 23743 16478 23763
rect 16548 23743 16550 23763
rect 16596 23743 16598 23763
rect 16692 23743 16694 23763
rect 16764 23743 16766 23763
rect 16788 23743 16790 23763
rect 16884 23743 16886 23763
rect 16908 23743 16910 23763
rect 17028 23743 17030 23763
rect 17124 23743 17126 23763
rect 17196 23743 17198 23763
rect 17220 23743 17222 23763
rect 17292 23743 17294 23763
rect 17316 23743 17318 23763
rect 17964 23743 17966 23763
rect 18060 23744 18062 23763
rect 18132 23744 18134 23763
rect 18228 23744 18230 23763
rect 18492 23744 18494 23763
rect 18540 23744 18542 23763
rect 18025 23743 18083 23744
rect 18121 23743 18155 23744
rect -671 23739 4253 23743
rect -575 23734 -572 23739
rect -564 23736 -562 23739
rect -468 23736 -466 23739
rect -564 23734 -561 23736
rect -575 23726 -571 23734
rect -585 23720 -575 23726
rect -565 23720 -561 23734
rect -468 23720 -465 23736
rect -479 23719 -445 23720
rect -132 23719 -130 23739
rect 84 23719 86 23739
rect 180 23719 182 23739
rect 468 23719 470 23739
rect 492 23719 494 23739
rect 564 23719 566 23739
rect 588 23719 590 23739
rect 660 23719 662 23739
rect 708 23719 710 23739
rect 948 23719 950 23739
rect 1044 23719 1046 23739
rect 1092 23719 1094 23739
rect 1140 23719 1142 23739
rect 1308 23719 1310 23739
rect 1356 23719 1358 23739
rect 1572 23719 1574 23739
rect 1860 23719 1862 23739
rect 1956 23719 1958 23739
rect 2052 23719 2054 23739
rect 2148 23719 2150 23739
rect 2244 23719 2246 23739
rect 2340 23719 2342 23739
rect 2436 23719 2438 23739
rect 2532 23719 2534 23739
rect 2628 23719 2630 23739
rect 2724 23719 2726 23739
rect 2940 23719 2942 23739
rect 2988 23719 2990 23739
rect 3324 23719 3326 23739
rect 3540 23719 3542 23739
rect 3780 23719 3782 23739
rect 4068 23719 4070 23739
rect 4164 23719 4166 23739
rect 4239 23736 4253 23739
rect 4263 23739 11357 23743
rect 4263 23736 4277 23739
rect 4308 23719 4310 23739
rect 4932 23719 4934 23739
rect 4980 23719 4982 23739
rect 5028 23719 5030 23739
rect 5124 23719 5126 23739
rect 5148 23719 5150 23739
rect 5220 23719 5222 23739
rect 5244 23719 5246 23739
rect 5460 23719 5462 23739
rect 5508 23719 5510 23739
rect 5556 23719 5558 23739
rect 5652 23719 5654 23739
rect 5748 23719 5750 23739
rect 5761 23734 5764 23739
rect 5771 23720 5774 23734
rect 5772 23719 5774 23720
rect 5844 23719 5846 23739
rect 5892 23736 5894 23739
rect 5892 23719 5895 23736
rect 6276 23719 6278 23739
rect 6300 23719 6302 23739
rect 6372 23719 6374 23739
rect 6396 23719 6398 23739
rect 6492 23719 6494 23739
rect 6516 23719 6518 23739
rect 6588 23719 6590 23739
rect 6612 23719 6614 23739
rect 6636 23719 6638 23739
rect 6708 23719 6710 23739
rect 6804 23719 6806 23739
rect 6900 23719 6902 23739
rect 7164 23719 7166 23739
rect 7284 23719 7286 23739
rect 7380 23719 7382 23739
rect 7404 23719 7406 23739
rect 7476 23719 7478 23739
rect 7500 23719 7502 23739
rect 7572 23719 7574 23739
rect 7596 23719 7598 23739
rect 7668 23719 7670 23739
rect 7692 23719 7694 23739
rect 7908 23719 7910 23739
rect 8124 23719 8126 23739
rect 8220 23719 8222 23739
rect 8316 23719 8318 23739
rect 8412 23719 8414 23739
rect 8700 23719 8702 23739
rect 8748 23719 8750 23739
rect 8796 23719 8798 23739
rect 8844 23719 8846 23739
rect 8868 23719 8870 23739
rect 9516 23719 9518 23739
rect 9684 23719 9686 23739
rect 9780 23719 9782 23739
rect 9804 23719 9806 23739
rect 9828 23719 9830 23739
rect 10044 23719 10046 23739
rect 10140 23719 10142 23739
rect 10236 23719 10238 23739
rect 10332 23719 10334 23739
rect 10369 23734 10372 23739
rect 10380 23734 10382 23739
rect 10379 23720 10382 23734
rect 10428 23719 10430 23739
rect 10452 23719 10455 23736
rect 10524 23719 10526 23739
rect 10548 23719 10550 23739
rect 10620 23719 10622 23739
rect 10644 23719 10646 23739
rect 10716 23719 10718 23739
rect 10860 23719 10862 23739
rect 10956 23719 10958 23739
rect 11052 23719 11054 23739
rect 11100 23719 11102 23739
rect 11148 23719 11150 23739
rect 11220 23719 11222 23739
rect 11244 23719 11246 23739
rect 11340 23719 11342 23739
rect 11343 23736 11357 23739
rect 11364 23739 18155 23743
rect 18217 23743 18251 23744
rect 18385 23743 18419 23744
rect 18217 23739 18419 23743
rect 18433 23743 18467 23744
rect 18481 23743 18515 23744
rect 18433 23739 18515 23743
rect 18529 23743 18563 23744
rect 18636 23743 18638 23763
rect 18732 23743 18734 23763
rect 18828 23743 18830 23763
rect 18924 23743 18926 23763
rect 18972 23743 18974 23763
rect 19068 23743 19070 23763
rect 19095 23760 19109 23763
rect 19140 23743 19142 23763
rect 19164 23743 19166 23763
rect 19236 23743 19238 23763
rect 19260 23744 19262 23763
rect 19249 23743 19283 23744
rect 18529 23739 19283 23743
rect 19297 23743 19331 23744
rect 19489 23743 19523 23744
rect 19297 23739 19523 23743
rect 11364 23736 11381 23739
rect 11364 23719 11366 23736
rect 11508 23719 11510 23739
rect 11593 23719 11651 23720
rect 11676 23719 11678 23739
rect 11724 23719 11726 23739
rect 11796 23719 11798 23739
rect 12060 23719 12062 23739
rect 12276 23719 12278 23739
rect 12372 23719 12374 23739
rect 12468 23719 12470 23739
rect 12564 23719 12566 23739
rect 12780 23719 12782 23739
rect 12876 23719 12878 23739
rect 13044 23719 13046 23739
rect 13164 23719 13166 23739
rect 13260 23719 13262 23739
rect 13332 23719 13334 23739
rect 13356 23719 13358 23739
rect 13500 23719 13502 23739
rect 13572 23719 13574 23739
rect 13836 23719 13838 23739
rect 13932 23719 13934 23739
rect 14004 23719 14006 23739
rect 14028 23719 14030 23739
rect 14172 23719 14174 23739
rect 14940 23719 14942 23739
rect 15036 23719 15038 23739
rect 15276 23719 15278 23739
rect 15372 23719 15374 23739
rect 15468 23719 15470 23739
rect 15564 23719 15566 23739
rect 15660 23719 15662 23739
rect 15684 23719 15686 23739
rect 15732 23719 15734 23739
rect 15756 23719 15758 23739
rect 15780 23719 15782 23739
rect 15828 23719 15830 23739
rect 15852 23719 15854 23739
rect 15876 23719 15878 23739
rect 15948 23719 15950 23739
rect 15972 23719 15974 23739
rect 16044 23719 16046 23739
rect 16068 23719 16070 23739
rect 16164 23719 16166 23739
rect 16260 23719 16262 23739
rect 16284 23719 16286 23739
rect 16380 23719 16382 23739
rect 16476 23719 16478 23739
rect 16548 23719 16550 23739
rect 16596 23719 16598 23739
rect 16692 23719 16694 23739
rect 16764 23719 16766 23739
rect 16788 23719 16790 23739
rect 16884 23719 16886 23739
rect 16908 23719 16910 23739
rect 17028 23719 17030 23739
rect 17124 23719 17126 23739
rect 17196 23719 17198 23739
rect 17220 23719 17222 23739
rect 17292 23719 17294 23739
rect 17316 23719 17318 23739
rect 17964 23720 17966 23739
rect 18049 23734 18052 23739
rect 18060 23734 18062 23739
rect 18121 23734 18124 23739
rect 18132 23736 18134 23739
rect 18132 23734 18135 23736
rect 18217 23734 18220 23739
rect 18228 23736 18230 23739
rect 18228 23734 18231 23736
rect 18481 23734 18484 23739
rect 18492 23736 18494 23739
rect 18492 23734 18495 23736
rect 18529 23734 18532 23739
rect 18540 23736 18542 23739
rect 18636 23736 18638 23739
rect 18540 23734 18543 23736
rect 18059 23720 18062 23734
rect 18131 23726 18135 23734
rect 18145 23726 18149 23734
rect 18131 23720 18145 23726
rect 18227 23720 18231 23734
rect 18491 23720 18495 23734
rect 18539 23720 18543 23734
rect 18636 23720 18639 23736
rect 17857 23719 17891 23720
rect -479 23715 5861 23719
rect -479 23712 -475 23715
rect -468 23712 -465 23715
rect -359 23695 -325 23696
rect -132 23695 -130 23715
rect 84 23695 86 23715
rect 180 23695 182 23715
rect 468 23695 470 23715
rect 492 23695 494 23715
rect 505 23695 563 23696
rect 564 23695 566 23715
rect 588 23695 590 23715
rect 660 23695 662 23715
rect 708 23695 710 23715
rect 948 23695 950 23715
rect 1044 23695 1046 23715
rect 1092 23695 1094 23715
rect 1140 23695 1142 23715
rect 1308 23695 1310 23715
rect 1356 23695 1358 23715
rect 1572 23695 1574 23715
rect 1860 23695 1862 23715
rect 1956 23695 1958 23715
rect 2052 23695 2054 23715
rect 2148 23695 2150 23715
rect 2244 23695 2246 23715
rect 2340 23695 2342 23715
rect 2436 23695 2438 23715
rect 2532 23695 2534 23715
rect 2628 23695 2630 23715
rect 2724 23695 2726 23715
rect 2940 23695 2942 23715
rect 2988 23695 2990 23715
rect 3324 23695 3326 23715
rect 3540 23695 3542 23715
rect 3780 23695 3782 23715
rect 4068 23695 4070 23715
rect 4164 23695 4166 23715
rect 4308 23695 4310 23715
rect 4932 23695 4934 23715
rect 4980 23695 4982 23715
rect 5028 23695 5030 23715
rect 5124 23695 5126 23715
rect 5148 23695 5150 23715
rect 5220 23696 5222 23715
rect 5185 23695 5243 23696
rect 5244 23695 5246 23715
rect 5460 23695 5462 23715
rect 5508 23695 5510 23715
rect 5556 23695 5558 23715
rect 5652 23695 5654 23715
rect 5703 23712 5717 23715
rect 5748 23695 5750 23715
rect 5772 23695 5774 23715
rect 5844 23695 5846 23715
rect 5847 23712 5861 23715
rect 5871 23715 10445 23719
rect 5871 23712 5885 23715
rect 5892 23712 5895 23715
rect 6276 23695 6278 23715
rect 6300 23695 6302 23715
rect 6372 23695 6374 23715
rect 6396 23695 6398 23715
rect 6492 23695 6494 23715
rect 6516 23695 6518 23715
rect 6588 23695 6590 23715
rect 6612 23695 6614 23715
rect 6636 23695 6638 23715
rect 6708 23695 6710 23715
rect 6804 23695 6806 23715
rect 6900 23695 6902 23715
rect 7164 23695 7166 23715
rect 7284 23695 7286 23715
rect 7380 23695 7382 23715
rect 7404 23695 7406 23715
rect 7476 23695 7478 23715
rect 7500 23695 7502 23715
rect 7572 23695 7574 23715
rect 7596 23695 7598 23715
rect 7668 23695 7670 23715
rect 7692 23695 7694 23715
rect 7908 23695 7910 23715
rect 8124 23695 8126 23715
rect 8220 23695 8222 23715
rect 8316 23695 8318 23715
rect 8412 23695 8414 23715
rect 8700 23695 8702 23715
rect 8748 23695 8750 23715
rect 8796 23695 8798 23715
rect 8844 23695 8846 23715
rect 8868 23695 8870 23715
rect 9516 23695 9518 23715
rect 9684 23695 9686 23715
rect 9780 23695 9782 23715
rect 9804 23695 9806 23715
rect 9828 23695 9830 23715
rect 10044 23695 10046 23715
rect 10140 23695 10142 23715
rect 10236 23695 10238 23715
rect 10332 23695 10334 23715
rect 10428 23695 10430 23715
rect 10431 23712 10445 23715
rect 10452 23715 17891 23719
rect 17953 23719 17987 23720
rect 18001 23719 18035 23720
rect 17953 23715 18035 23719
rect 18625 23719 18659 23720
rect 18732 23719 18734 23739
rect 18828 23719 18830 23739
rect 18924 23720 18926 23739
rect 18972 23720 18974 23739
rect 19068 23720 19070 23739
rect 19140 23720 19142 23739
rect 19164 23720 19166 23739
rect 19236 23720 19238 23739
rect 19249 23734 19252 23739
rect 19260 23734 19262 23739
rect 19259 23720 19262 23734
rect 18913 23719 18947 23720
rect 18625 23715 18947 23719
rect 18961 23719 18995 23720
rect 19033 23719 19091 23720
rect 19129 23719 19187 23720
rect 19225 23719 19259 23720
rect 18961 23715 19259 23719
rect 10452 23712 10469 23715
rect 10452 23695 10454 23712
rect 10524 23695 10526 23715
rect 10548 23695 10550 23715
rect 10620 23695 10622 23715
rect 10644 23695 10646 23715
rect 10716 23695 10718 23715
rect 10860 23695 10862 23715
rect 10956 23695 10958 23715
rect 11052 23695 11054 23715
rect 11100 23695 11102 23715
rect 11148 23695 11150 23715
rect 11220 23695 11222 23715
rect 11244 23695 11246 23715
rect 11340 23695 11342 23715
rect 11364 23695 11366 23715
rect 11508 23695 11510 23715
rect 11593 23710 11596 23715
rect 11603 23696 11606 23710
rect 11569 23695 11603 23696
rect 11604 23695 11606 23696
rect 11676 23695 11678 23715
rect 11724 23712 11726 23715
rect 11700 23695 11703 23712
rect 11724 23695 11727 23712
rect 11796 23695 11798 23715
rect 12060 23695 12062 23715
rect 12276 23695 12278 23715
rect 12372 23695 12374 23715
rect 12468 23695 12470 23715
rect 12564 23695 12566 23715
rect 12780 23695 12782 23715
rect 12876 23695 12878 23715
rect 13044 23695 13046 23715
rect 13164 23695 13166 23715
rect 13260 23695 13262 23715
rect 13332 23695 13334 23715
rect 13356 23695 13358 23715
rect 13500 23695 13502 23715
rect 13572 23695 13574 23715
rect 13836 23695 13838 23715
rect 13932 23695 13934 23715
rect 14004 23695 14006 23715
rect 14028 23695 14030 23715
rect 14172 23695 14174 23715
rect 14940 23695 14942 23715
rect 15036 23695 15038 23715
rect 15276 23695 15278 23715
rect 15372 23695 15374 23715
rect 15468 23695 15470 23715
rect 15564 23695 15566 23715
rect 15660 23695 15662 23715
rect 15684 23695 15686 23715
rect 15732 23695 15734 23715
rect 15756 23695 15758 23715
rect 15780 23695 15782 23715
rect 15828 23695 15830 23715
rect 15852 23695 15854 23715
rect 15876 23695 15878 23715
rect 15948 23695 15950 23715
rect 15972 23695 15974 23715
rect 16044 23695 16046 23715
rect 16068 23695 16070 23715
rect 16164 23695 16166 23715
rect 16260 23695 16262 23715
rect 16284 23695 16286 23715
rect 16380 23695 16382 23715
rect 16476 23695 16478 23715
rect 16548 23695 16550 23715
rect 16596 23695 16598 23715
rect 16692 23695 16694 23715
rect 16764 23695 16766 23715
rect 16788 23695 16790 23715
rect 16884 23695 16886 23715
rect 16908 23695 16910 23715
rect 17028 23695 17030 23715
rect 17124 23695 17126 23715
rect 17196 23695 17198 23715
rect 17220 23695 17222 23715
rect 17292 23695 17294 23715
rect 17316 23695 17318 23715
rect 17953 23710 17956 23715
rect 17964 23712 17966 23715
rect 18625 23712 18629 23715
rect 18636 23712 18639 23715
rect 18732 23712 18734 23715
rect 17964 23710 17967 23712
rect 17963 23696 17967 23710
rect 18732 23696 18735 23712
rect 17449 23695 17483 23696
rect -359 23691 11693 23695
rect -239 23671 -205 23672
rect -132 23671 -130 23691
rect 84 23671 86 23691
rect 180 23671 182 23691
rect 468 23671 470 23691
rect 492 23671 494 23691
rect 564 23671 566 23691
rect 588 23672 590 23691
rect 612 23672 615 23688
rect 660 23672 662 23691
rect 708 23672 710 23691
rect 577 23671 605 23672
rect -239 23667 605 23671
rect -132 23664 -130 23667
rect -132 23648 -129 23664
rect -143 23647 -109 23648
rect -95 23647 -61 23648
rect -143 23643 -61 23647
rect -23 23647 11 23648
rect 84 23647 86 23667
rect 180 23647 182 23667
rect 468 23647 470 23667
rect 492 23648 494 23667
rect 564 23648 566 23667
rect 577 23662 580 23667
rect 588 23662 590 23667
rect 591 23664 605 23667
rect 612 23671 635 23672
rect 649 23671 683 23672
rect 612 23667 683 23671
rect 697 23671 731 23672
rect 769 23671 803 23672
rect 697 23667 803 23671
rect 841 23671 875 23672
rect 948 23671 950 23691
rect 1044 23671 1046 23691
rect 1092 23671 1094 23691
rect 1140 23671 1142 23691
rect 1201 23671 1235 23672
rect 1308 23671 1310 23691
rect 1321 23671 1355 23672
rect 1356 23671 1358 23691
rect 1572 23671 1574 23691
rect 1860 23671 1862 23691
rect 1956 23671 1958 23691
rect 2052 23671 2054 23691
rect 2148 23671 2150 23691
rect 2244 23671 2246 23691
rect 2340 23671 2342 23691
rect 2436 23671 2438 23691
rect 2532 23671 2534 23691
rect 2628 23671 2630 23691
rect 2724 23671 2726 23691
rect 2940 23671 2942 23691
rect 2988 23671 2990 23691
rect 3324 23671 3326 23691
rect 3540 23671 3542 23691
rect 3780 23671 3782 23691
rect 4068 23671 4070 23691
rect 4164 23671 4166 23691
rect 4308 23671 4310 23691
rect 4932 23671 4934 23691
rect 4980 23672 4982 23691
rect 4969 23671 5003 23672
rect 5028 23671 5030 23691
rect 5124 23671 5126 23691
rect 5148 23671 5150 23691
rect 5185 23686 5188 23691
rect 5209 23686 5212 23691
rect 5220 23686 5222 23691
rect 5195 23672 5198 23686
rect 5219 23672 5222 23686
rect 5196 23671 5198 23672
rect 5244 23671 5246 23691
rect 5292 23671 5295 23688
rect 5460 23671 5462 23691
rect 5508 23671 5510 23691
rect 5556 23671 5558 23691
rect 5652 23671 5654 23691
rect 5748 23671 5750 23691
rect 5772 23671 5774 23691
rect 5844 23671 5846 23691
rect 6276 23671 6278 23691
rect 6300 23671 6302 23691
rect 6372 23671 6374 23691
rect 6396 23671 6398 23691
rect 6492 23671 6494 23691
rect 6516 23671 6518 23691
rect 6588 23671 6590 23691
rect 6612 23671 6614 23691
rect 6636 23671 6638 23691
rect 6708 23671 6710 23691
rect 6804 23671 6806 23691
rect 6900 23671 6902 23691
rect 7164 23671 7166 23691
rect 7284 23671 7286 23691
rect 7380 23671 7382 23691
rect 7404 23671 7406 23691
rect 7476 23671 7478 23691
rect 7500 23671 7502 23691
rect 7572 23671 7574 23691
rect 7596 23671 7598 23691
rect 7668 23671 7670 23691
rect 7692 23671 7694 23691
rect 7908 23671 7910 23691
rect 8124 23671 8126 23691
rect 8220 23671 8222 23691
rect 8316 23671 8318 23691
rect 8412 23671 8414 23691
rect 8700 23671 8702 23691
rect 8748 23671 8750 23691
rect 8796 23671 8798 23691
rect 8844 23671 8846 23691
rect 8868 23671 8870 23691
rect 9516 23671 9518 23691
rect 9684 23671 9686 23691
rect 9780 23671 9782 23691
rect 9804 23671 9806 23691
rect 9828 23671 9830 23691
rect 10044 23671 10046 23691
rect 10140 23671 10142 23691
rect 10236 23671 10238 23691
rect 10332 23671 10334 23691
rect 10428 23671 10430 23691
rect 10452 23671 10454 23691
rect 10524 23671 10526 23691
rect 10548 23671 10550 23691
rect 10620 23671 10622 23691
rect 10644 23671 10646 23691
rect 10716 23671 10718 23691
rect 10860 23671 10862 23691
rect 10956 23671 10958 23691
rect 11052 23671 11054 23691
rect 11100 23671 11102 23691
rect 11148 23671 11150 23691
rect 11220 23671 11222 23691
rect 11244 23671 11246 23691
rect 11340 23671 11342 23691
rect 11364 23671 11366 23691
rect 11508 23671 11510 23691
rect 11604 23671 11606 23691
rect 11676 23688 11678 23691
rect 11679 23688 11693 23691
rect 11700 23691 17483 23695
rect 18721 23695 18755 23696
rect 18828 23695 18830 23715
rect 18913 23710 18916 23715
rect 18924 23710 18926 23715
rect 18961 23710 18964 23715
rect 18972 23710 18974 23715
rect 18923 23696 18926 23710
rect 18971 23696 18974 23710
rect 19057 23710 19060 23715
rect 19068 23712 19070 23715
rect 19068 23710 19071 23712
rect 19129 23710 19132 23715
rect 19140 23712 19142 23715
rect 19140 23710 19143 23712
rect 19057 23702 19061 23710
rect 19047 23696 19057 23702
rect 19067 23696 19071 23710
rect 19139 23702 19143 23710
rect 19153 23710 19156 23715
rect 19164 23712 19166 23715
rect 19164 23710 19167 23712
rect 19225 23710 19228 23715
rect 19236 23712 19238 23715
rect 19236 23710 19239 23712
rect 19153 23702 19157 23710
rect 19139 23696 19153 23702
rect 19163 23696 19167 23710
rect 19235 23702 19239 23710
rect 19249 23702 19253 23710
rect 19235 23696 19249 23702
rect 18889 23695 18923 23696
rect 18721 23691 18923 23695
rect 11700 23688 11717 23691
rect 11724 23688 11727 23691
rect 11676 23671 11679 23688
rect 11700 23671 11702 23688
rect 11796 23671 11798 23691
rect 11929 23671 11987 23672
rect 12060 23671 12062 23691
rect 12276 23671 12278 23691
rect 12372 23671 12374 23691
rect 12468 23671 12470 23691
rect 12564 23671 12566 23691
rect 12780 23671 12782 23691
rect 12876 23671 12878 23691
rect 13044 23671 13046 23691
rect 13164 23671 13166 23691
rect 13260 23671 13262 23691
rect 13332 23671 13334 23691
rect 13356 23671 13358 23691
rect 13500 23671 13502 23691
rect 13572 23671 13574 23691
rect 13836 23671 13838 23691
rect 13932 23671 13934 23691
rect 14004 23671 14006 23691
rect 14028 23671 14030 23691
rect 14172 23671 14174 23691
rect 14940 23671 14942 23691
rect 15036 23671 15038 23691
rect 15276 23671 15278 23691
rect 15372 23671 15374 23691
rect 15468 23671 15470 23691
rect 15564 23671 15566 23691
rect 15660 23671 15662 23691
rect 15684 23671 15686 23691
rect 15732 23671 15734 23691
rect 15756 23671 15758 23691
rect 15780 23671 15782 23691
rect 15828 23671 15830 23691
rect 15852 23671 15854 23691
rect 15876 23671 15878 23691
rect 15948 23671 15950 23691
rect 15972 23671 15974 23691
rect 16044 23671 16046 23691
rect 16068 23671 16070 23691
rect 16164 23671 16166 23691
rect 16260 23671 16262 23691
rect 16284 23671 16286 23691
rect 16380 23671 16382 23691
rect 16476 23671 16478 23691
rect 16548 23671 16550 23691
rect 16596 23671 16598 23691
rect 16692 23671 16694 23691
rect 16764 23671 16766 23691
rect 16788 23671 16790 23691
rect 16884 23671 16886 23691
rect 16908 23671 16910 23691
rect 17028 23671 17030 23691
rect 17124 23671 17126 23691
rect 17196 23671 17198 23691
rect 17220 23671 17222 23691
rect 17292 23671 17294 23691
rect 17316 23672 17318 23691
rect 18721 23688 18725 23691
rect 18732 23688 18735 23691
rect 18828 23688 18830 23691
rect 18828 23672 18831 23688
rect 17305 23671 17339 23672
rect 841 23667 5285 23671
rect 612 23664 629 23667
rect 601 23662 604 23664
rect 612 23662 614 23664
rect 649 23662 652 23667
rect 660 23662 662 23667
rect 697 23662 700 23667
rect 708 23664 710 23667
rect 948 23664 950 23667
rect 708 23662 711 23664
rect 587 23648 590 23662
rect 611 23648 614 23662
rect 659 23648 662 23662
rect 673 23654 677 23662
rect 663 23648 673 23654
rect 707 23648 711 23662
rect 793 23654 797 23662
rect 865 23654 869 23662
rect 783 23648 793 23654
rect 855 23648 865 23654
rect 948 23648 951 23664
rect 1044 23648 1046 23667
rect 1092 23648 1094 23667
rect 1140 23648 1142 23667
rect 1308 23664 1310 23667
rect 481 23647 539 23648
rect 553 23647 587 23648
rect -23 23643 587 23647
rect 937 23647 971 23648
rect 985 23647 1019 23648
rect 937 23643 1019 23647
rect 1033 23647 1067 23648
rect 1081 23647 1115 23648
rect 1033 23643 1115 23647
rect 1129 23647 1163 23648
rect 1308 23647 1311 23664
rect 1356 23647 1358 23667
rect 1572 23647 1574 23667
rect 1657 23647 1715 23648
rect 1860 23647 1862 23667
rect 1956 23647 1958 23667
rect 2052 23647 2054 23667
rect 2148 23647 2150 23667
rect 2244 23647 2246 23667
rect 2340 23647 2342 23667
rect 2436 23647 2438 23667
rect 2532 23647 2534 23667
rect 2628 23647 2630 23667
rect 2724 23647 2726 23667
rect 2940 23647 2942 23667
rect 2988 23647 2990 23667
rect 3324 23647 3326 23667
rect 3540 23647 3542 23667
rect 3780 23647 3782 23667
rect 4068 23647 4070 23667
rect 4164 23647 4166 23667
rect 4308 23647 4310 23667
rect 4932 23647 4934 23667
rect 4969 23662 4972 23667
rect 4980 23662 4982 23667
rect 4979 23648 4982 23662
rect 5028 23647 5030 23667
rect 5124 23647 5126 23667
rect 5148 23647 5150 23667
rect 5196 23647 5198 23667
rect 5244 23647 5246 23667
rect 5271 23664 5285 23667
rect 5292 23667 17339 23671
rect 18817 23671 18851 23672
rect 18865 23671 18899 23672
rect 18817 23667 18899 23671
rect 5292 23664 5309 23667
rect 5292 23647 5294 23664
rect 5460 23647 5462 23667
rect 5508 23647 5510 23667
rect 5556 23647 5558 23667
rect 5652 23647 5654 23667
rect 5748 23647 5750 23667
rect 5772 23647 5774 23667
rect 5844 23647 5846 23667
rect 6276 23647 6278 23667
rect 6300 23647 6302 23667
rect 6372 23647 6374 23667
rect 6396 23647 6398 23667
rect 6492 23647 6494 23667
rect 6516 23647 6518 23667
rect 6588 23647 6590 23667
rect 6612 23647 6614 23667
rect 6636 23647 6638 23667
rect 6708 23647 6710 23667
rect 6804 23647 6806 23667
rect 6900 23647 6902 23667
rect 7164 23647 7166 23667
rect 7284 23647 7286 23667
rect 7380 23647 7382 23667
rect 7404 23647 7406 23667
rect 7476 23647 7478 23667
rect 7500 23647 7502 23667
rect 7572 23647 7574 23667
rect 7596 23647 7598 23667
rect 7668 23647 7670 23667
rect 7692 23647 7694 23667
rect 7908 23647 7910 23667
rect 8124 23647 8126 23667
rect 8220 23647 8222 23667
rect 8316 23647 8318 23667
rect 8412 23647 8414 23667
rect 8700 23647 8702 23667
rect 8748 23647 8750 23667
rect 8796 23647 8798 23667
rect 8844 23647 8846 23667
rect 8868 23647 8870 23667
rect 9516 23647 9518 23667
rect 9684 23647 9686 23667
rect 9780 23647 9782 23667
rect 9804 23647 9806 23667
rect 9828 23647 9830 23667
rect 9913 23647 9971 23648
rect 10044 23647 10046 23667
rect 10140 23647 10142 23667
rect 10236 23647 10238 23667
rect 10332 23647 10334 23667
rect 10428 23647 10430 23667
rect 10452 23647 10454 23667
rect 10524 23647 10526 23667
rect 10548 23647 10550 23667
rect 10620 23647 10622 23667
rect 10644 23647 10646 23667
rect 10716 23647 10718 23667
rect 10860 23647 10862 23667
rect 10956 23647 10958 23667
rect 11052 23647 11054 23667
rect 11100 23647 11102 23667
rect 11148 23647 11150 23667
rect 11220 23647 11222 23667
rect 11244 23647 11246 23667
rect 11340 23647 11342 23667
rect 11364 23647 11366 23667
rect 11508 23647 11510 23667
rect 11604 23647 11606 23667
rect 11655 23664 11669 23667
rect 11676 23664 11679 23667
rect 11700 23647 11702 23667
rect 11796 23647 11798 23667
rect 11929 23662 11932 23667
rect 12060 23664 12062 23667
rect 11939 23648 11942 23662
rect 11940 23647 11942 23648
rect 12060 23647 12063 23664
rect 12276 23647 12278 23667
rect 12372 23647 12374 23667
rect 12468 23647 12470 23667
rect 12564 23647 12566 23667
rect 12780 23647 12782 23667
rect 12876 23647 12878 23667
rect 13044 23647 13046 23667
rect 13164 23647 13166 23667
rect 13260 23647 13262 23667
rect 13332 23647 13334 23667
rect 13356 23647 13358 23667
rect 13500 23647 13502 23667
rect 13572 23647 13574 23667
rect 13836 23647 13838 23667
rect 13932 23647 13934 23667
rect 14004 23647 14006 23667
rect 14028 23647 14030 23667
rect 14172 23647 14174 23667
rect 14940 23647 14942 23667
rect 15036 23647 15038 23667
rect 15276 23647 15278 23667
rect 15372 23647 15374 23667
rect 15468 23647 15470 23667
rect 15564 23647 15566 23667
rect 15660 23647 15662 23667
rect 15684 23647 15686 23667
rect 15732 23647 15734 23667
rect 15756 23647 15758 23667
rect 15780 23647 15782 23667
rect 15828 23647 15830 23667
rect 15852 23647 15854 23667
rect 15876 23647 15878 23667
rect 15948 23647 15950 23667
rect 15972 23647 15974 23667
rect 16044 23647 16046 23667
rect 16068 23647 16070 23667
rect 16164 23647 16166 23667
rect 16260 23647 16262 23667
rect 16284 23647 16286 23667
rect 16380 23647 16382 23667
rect 16476 23647 16478 23667
rect 16548 23647 16550 23667
rect 16596 23647 16598 23667
rect 16692 23647 16694 23667
rect 16764 23647 16766 23667
rect 16788 23647 16790 23667
rect 16884 23647 16886 23667
rect 16908 23647 16910 23667
rect 17028 23647 17030 23667
rect 17124 23647 17126 23667
rect 17196 23647 17198 23667
rect 17220 23647 17222 23667
rect 17292 23648 17294 23667
rect 17305 23662 17308 23667
rect 17316 23662 17318 23667
rect 18817 23664 18821 23667
rect 18828 23664 18831 23667
rect 17315 23648 17318 23662
rect 17281 23647 17315 23648
rect 1129 23643 12029 23647
rect -143 23640 -139 23643
rect -132 23640 -129 23643
rect 84 23640 86 23643
rect 1 23630 5 23638
rect -9 23624 1 23630
rect 84 23624 87 23640
rect 73 23623 107 23624
rect 180 23623 182 23643
rect 468 23624 470 23643
rect 481 23638 484 23643
rect 492 23638 494 23643
rect 553 23638 556 23643
rect 564 23638 566 23643
rect 937 23640 941 23643
rect 948 23640 951 23643
rect 1033 23638 1036 23643
rect 1044 23640 1046 23643
rect 1044 23638 1047 23640
rect 1081 23638 1084 23643
rect 1092 23640 1094 23643
rect 1092 23638 1095 23640
rect 1129 23638 1132 23643
rect 1140 23640 1142 23643
rect 1287 23640 1301 23643
rect 1308 23640 1311 23643
rect 1140 23638 1143 23640
rect 491 23624 494 23638
rect 563 23624 566 23638
rect 577 23630 581 23638
rect 567 23624 577 23630
rect 1043 23624 1047 23638
rect 1091 23624 1095 23638
rect 1139 23624 1143 23638
rect 1356 23624 1358 23643
rect 1407 23640 1421 23643
rect 361 23623 419 23624
rect 457 23623 491 23624
rect 73 23619 491 23623
rect 1249 23623 1283 23624
rect 1297 23623 1331 23624
rect 1249 23619 1331 23623
rect 1345 23623 1379 23624
rect 1572 23623 1574 23643
rect 1657 23638 1660 23643
rect 1667 23624 1670 23638
rect 1668 23623 1670 23624
rect 1764 23623 1767 23640
rect 1860 23623 1862 23643
rect 1956 23623 1958 23643
rect 2052 23623 2054 23643
rect 2148 23623 2150 23643
rect 2244 23623 2246 23643
rect 2340 23623 2342 23643
rect 2436 23623 2438 23643
rect 2532 23623 2534 23643
rect 2628 23623 2630 23643
rect 2724 23623 2726 23643
rect 2809 23623 2867 23624
rect 2940 23623 2942 23643
rect 2988 23623 2990 23643
rect 3073 23623 3131 23624
rect 3324 23623 3326 23643
rect 3540 23623 3542 23643
rect 3780 23623 3782 23643
rect 4068 23623 4070 23643
rect 4164 23623 4166 23643
rect 4308 23623 4310 23643
rect 4932 23623 4934 23643
rect 5028 23623 5030 23643
rect 5055 23640 5069 23643
rect 5124 23623 5126 23643
rect 5148 23623 5150 23643
rect 5196 23623 5198 23643
rect 5244 23623 5246 23643
rect 5292 23623 5294 23643
rect 5460 23623 5462 23643
rect 5508 23623 5510 23643
rect 5556 23623 5558 23643
rect 5652 23623 5654 23643
rect 5748 23623 5750 23643
rect 5772 23623 5774 23643
rect 5844 23623 5846 23643
rect 6276 23623 6278 23643
rect 6300 23623 6302 23643
rect 6372 23623 6374 23643
rect 6396 23623 6398 23643
rect 6492 23623 6494 23643
rect 6516 23623 6518 23643
rect 6588 23623 6590 23643
rect 6612 23623 6614 23643
rect 6636 23623 6638 23643
rect 6708 23623 6710 23643
rect 6804 23623 6806 23643
rect 6900 23623 6902 23643
rect 7164 23623 7166 23643
rect 7284 23623 7286 23643
rect 7380 23623 7382 23643
rect 7404 23623 7406 23643
rect 7476 23623 7478 23643
rect 7500 23623 7502 23643
rect 7572 23623 7574 23643
rect 7596 23623 7598 23643
rect 7668 23623 7670 23643
rect 7692 23623 7694 23643
rect 7908 23623 7910 23643
rect 8124 23623 8126 23643
rect 8220 23623 8222 23643
rect 8316 23623 8318 23643
rect 8412 23623 8414 23643
rect 8700 23623 8702 23643
rect 8748 23623 8750 23643
rect 8796 23623 8798 23643
rect 8844 23623 8846 23643
rect 8868 23623 8870 23643
rect 9516 23623 9518 23643
rect 9684 23623 9686 23643
rect 9780 23623 9782 23643
rect 9804 23623 9806 23643
rect 9828 23623 9830 23643
rect 9913 23638 9916 23643
rect 10044 23640 10046 23643
rect 9923 23624 9926 23638
rect 9924 23623 9926 23624
rect 10020 23623 10023 23640
rect 10044 23623 10047 23640
rect 10140 23623 10142 23643
rect 10236 23623 10238 23643
rect 10332 23623 10334 23643
rect 10428 23623 10430 23643
rect 10452 23623 10454 23643
rect 10524 23623 10526 23643
rect 10548 23623 10550 23643
rect 10620 23623 10622 23643
rect 10644 23623 10646 23643
rect 10716 23623 10718 23643
rect 10860 23623 10862 23643
rect 10956 23623 10958 23643
rect 11052 23623 11054 23643
rect 11100 23623 11102 23643
rect 11148 23623 11150 23643
rect 11220 23623 11222 23643
rect 11244 23623 11246 23643
rect 11340 23623 11342 23643
rect 11364 23623 11366 23643
rect 11508 23623 11510 23643
rect 11604 23623 11606 23643
rect 11700 23623 11702 23643
rect 11796 23623 11798 23643
rect 11940 23623 11942 23643
rect 12015 23640 12029 23643
rect 12039 23643 17315 23647
rect 12039 23640 12053 23643
rect 12060 23640 12063 23643
rect 12276 23623 12278 23643
rect 12372 23623 12374 23643
rect 12468 23623 12470 23643
rect 12564 23623 12566 23643
rect 12780 23623 12782 23643
rect 12876 23623 12878 23643
rect 13044 23623 13046 23643
rect 13164 23623 13166 23643
rect 13260 23623 13262 23643
rect 13332 23623 13334 23643
rect 13356 23623 13358 23643
rect 13500 23623 13502 23643
rect 13572 23623 13574 23643
rect 13836 23623 13838 23643
rect 13932 23623 13934 23643
rect 14004 23623 14006 23643
rect 14028 23623 14030 23643
rect 14172 23623 14174 23643
rect 14940 23623 14942 23643
rect 15036 23623 15038 23643
rect 15276 23623 15278 23643
rect 15372 23623 15374 23643
rect 15468 23623 15470 23643
rect 15564 23623 15566 23643
rect 15660 23623 15662 23643
rect 15684 23623 15686 23643
rect 15732 23623 15734 23643
rect 15756 23623 15758 23643
rect 15780 23623 15782 23643
rect 15828 23623 15830 23643
rect 15852 23623 15854 23643
rect 15876 23623 15878 23643
rect 15948 23623 15950 23643
rect 15972 23623 15974 23643
rect 16044 23623 16046 23643
rect 16068 23623 16070 23643
rect 16164 23623 16166 23643
rect 16260 23623 16262 23643
rect 16284 23623 16286 23643
rect 16380 23623 16382 23643
rect 16476 23623 16478 23643
rect 16548 23623 16550 23643
rect 16596 23623 16598 23643
rect 16692 23623 16694 23643
rect 16764 23623 16766 23643
rect 16788 23623 16790 23643
rect 16884 23623 16886 23643
rect 16908 23623 16910 23643
rect 17028 23623 17030 23643
rect 17124 23623 17126 23643
rect 17196 23623 17198 23643
rect 17220 23624 17222 23643
rect 17281 23638 17284 23643
rect 17292 23638 17294 23643
rect 17291 23624 17294 23638
rect 17209 23623 17243 23624
rect 1345 23619 1757 23623
rect 73 23616 77 23619
rect 84 23616 87 23619
rect 180 23616 182 23619
rect 180 23600 183 23616
rect 457 23614 460 23619
rect 468 23616 470 23619
rect 468 23614 471 23616
rect 1345 23614 1348 23619
rect 1356 23616 1358 23619
rect 1356 23614 1359 23616
rect 467 23606 471 23614
rect 481 23606 485 23614
rect 467 23600 481 23606
rect 1355 23600 1359 23614
rect 169 23599 203 23600
rect 337 23599 371 23600
rect 169 23595 371 23599
rect 1465 23599 1499 23600
rect 1572 23599 1574 23619
rect 1668 23599 1670 23619
rect 1743 23616 1757 23619
rect 1764 23619 10013 23623
rect 1764 23616 1781 23619
rect 1764 23599 1766 23616
rect 1860 23599 1862 23619
rect 1956 23599 1958 23619
rect 2052 23599 2054 23619
rect 2148 23599 2150 23619
rect 2244 23599 2246 23619
rect 2340 23599 2342 23619
rect 2436 23599 2438 23619
rect 2532 23599 2534 23619
rect 2628 23599 2630 23619
rect 2724 23599 2726 23619
rect 2809 23614 2812 23619
rect 2940 23616 2942 23619
rect 2819 23600 2822 23614
rect 2820 23599 2822 23600
rect 2916 23599 2919 23616
rect 2940 23599 2943 23616
rect 2988 23599 2990 23619
rect 3073 23614 3076 23619
rect 3083 23600 3086 23614
rect 3084 23599 3086 23600
rect 3324 23599 3326 23619
rect 3540 23599 3542 23619
rect 3780 23599 3782 23619
rect 4068 23599 4070 23619
rect 4164 23599 4166 23619
rect 4308 23599 4310 23619
rect 4932 23599 4934 23619
rect 5028 23599 5030 23619
rect 5124 23599 5126 23619
rect 5148 23599 5150 23619
rect 5196 23599 5198 23619
rect 5244 23599 5246 23619
rect 5292 23599 5294 23619
rect 5460 23599 5462 23619
rect 5508 23599 5510 23619
rect 5556 23599 5558 23619
rect 5652 23599 5654 23619
rect 5748 23599 5750 23619
rect 5772 23599 5774 23619
rect 5844 23599 5846 23619
rect 6276 23599 6278 23619
rect 6300 23599 6302 23619
rect 6372 23599 6374 23619
rect 6396 23599 6398 23619
rect 6492 23599 6494 23619
rect 6516 23599 6518 23619
rect 6588 23599 6590 23619
rect 6612 23599 6614 23619
rect 6636 23599 6638 23619
rect 6708 23599 6710 23619
rect 6804 23599 6806 23619
rect 6900 23599 6902 23619
rect 7164 23599 7166 23619
rect 7284 23599 7286 23619
rect 7380 23600 7382 23619
rect 7369 23599 7403 23600
rect 7404 23599 7406 23619
rect 7476 23599 7478 23619
rect 7500 23599 7502 23619
rect 7572 23600 7574 23619
rect 7561 23599 7595 23600
rect 7596 23599 7598 23619
rect 7668 23599 7670 23619
rect 7692 23599 7694 23619
rect 7908 23599 7910 23619
rect 8124 23599 8126 23619
rect 8220 23599 8222 23619
rect 8316 23599 8318 23619
rect 8412 23599 8414 23619
rect 8700 23599 8702 23619
rect 8748 23599 8750 23619
rect 8796 23599 8798 23619
rect 8844 23599 8846 23619
rect 8868 23599 8870 23619
rect 9516 23599 9518 23619
rect 9684 23599 9686 23619
rect 9780 23599 9782 23619
rect 9804 23599 9806 23619
rect 9828 23599 9830 23619
rect 9924 23599 9926 23619
rect 9999 23616 10013 23619
rect 10020 23619 17243 23623
rect 10020 23616 10037 23619
rect 10044 23616 10047 23619
rect 10020 23599 10022 23616
rect 10140 23599 10142 23619
rect 10236 23599 10238 23619
rect 10332 23599 10334 23619
rect 10428 23599 10430 23619
rect 10452 23599 10454 23619
rect 10524 23599 10526 23619
rect 10548 23599 10550 23619
rect 10620 23599 10622 23619
rect 10644 23599 10646 23619
rect 10716 23599 10718 23619
rect 10860 23599 10862 23619
rect 10956 23599 10958 23619
rect 11052 23599 11054 23619
rect 11100 23599 11102 23619
rect 11148 23599 11150 23619
rect 11220 23599 11222 23619
rect 11244 23599 11246 23619
rect 11340 23599 11342 23619
rect 11364 23599 11366 23619
rect 11508 23599 11510 23619
rect 11604 23599 11606 23619
rect 11700 23599 11702 23619
rect 11796 23600 11798 23619
rect 11785 23599 11867 23600
rect 11940 23599 11942 23619
rect 12276 23599 12278 23619
rect 12372 23599 12374 23619
rect 12468 23599 12470 23619
rect 12564 23599 12566 23619
rect 12780 23599 12782 23619
rect 12876 23599 12878 23619
rect 13044 23599 13046 23619
rect 13164 23599 13166 23619
rect 13260 23599 13262 23619
rect 13332 23599 13334 23619
rect 13356 23599 13358 23619
rect 13500 23599 13502 23619
rect 13572 23599 13574 23619
rect 13836 23599 13838 23619
rect 13932 23599 13934 23619
rect 14004 23599 14006 23619
rect 14028 23599 14030 23619
rect 14172 23599 14174 23619
rect 14940 23599 14942 23619
rect 15036 23599 15038 23619
rect 15276 23599 15278 23619
rect 15372 23599 15374 23619
rect 15468 23599 15470 23619
rect 15564 23599 15566 23619
rect 15660 23599 15662 23619
rect 15684 23599 15686 23619
rect 15732 23599 15734 23619
rect 15756 23599 15758 23619
rect 15780 23599 15782 23619
rect 15828 23599 15830 23619
rect 15852 23599 15854 23619
rect 15876 23599 15878 23619
rect 15948 23599 15950 23619
rect 15972 23599 15974 23619
rect 16044 23599 16046 23619
rect 16068 23599 16070 23619
rect 16164 23599 16166 23619
rect 16260 23599 16262 23619
rect 16284 23599 16286 23619
rect 16380 23599 16382 23619
rect 16476 23599 16478 23619
rect 16548 23599 16550 23619
rect 16596 23599 16598 23619
rect 16692 23599 16694 23619
rect 16764 23599 16766 23619
rect 16788 23599 16790 23619
rect 16884 23599 16886 23619
rect 16908 23600 16910 23619
rect 16897 23599 16955 23600
rect 17028 23599 17030 23619
rect 17124 23600 17126 23619
rect 17196 23600 17198 23619
rect 17209 23614 17212 23619
rect 17220 23614 17222 23619
rect 17219 23600 17222 23614
rect 17113 23599 17171 23600
rect 17185 23599 17219 23600
rect 1465 23595 2909 23599
rect 169 23592 173 23595
rect 180 23592 183 23595
rect 1572 23592 1574 23595
rect 1572 23576 1575 23592
rect 1561 23575 1595 23576
rect 1668 23575 1670 23595
rect 1764 23575 1766 23595
rect 1860 23575 1862 23595
rect 1956 23575 1958 23595
rect 2052 23575 2054 23595
rect 2089 23575 2123 23576
rect 2148 23575 2150 23595
rect 2244 23575 2246 23595
rect 2340 23575 2342 23595
rect 2436 23575 2438 23595
rect 2532 23575 2534 23595
rect 2628 23575 2630 23595
rect 2724 23575 2726 23595
rect 2820 23575 2822 23595
rect 2895 23592 2909 23595
rect 2916 23595 3173 23599
rect 2916 23592 2933 23595
rect 2940 23592 2943 23595
rect 2916 23575 2918 23592
rect 2988 23575 2990 23595
rect 3084 23575 3086 23595
rect 3159 23592 3173 23595
rect 3183 23595 17219 23599
rect 3183 23592 3197 23595
rect 3324 23575 3326 23595
rect 3540 23575 3542 23595
rect 3780 23575 3782 23595
rect 4009 23575 4043 23576
rect 4068 23575 4070 23595
rect 4164 23575 4166 23595
rect 4308 23575 4310 23595
rect 4932 23575 4934 23595
rect 5028 23575 5030 23595
rect 5124 23575 5126 23595
rect 5148 23575 5150 23595
rect 5196 23575 5198 23595
rect 5244 23575 5246 23595
rect 5292 23575 5294 23595
rect 5460 23575 5462 23595
rect 5508 23575 5510 23595
rect 5556 23575 5558 23595
rect 5652 23575 5654 23595
rect 5748 23575 5750 23595
rect 5772 23575 5774 23595
rect 5844 23575 5846 23595
rect 6145 23575 6179 23576
rect 6276 23575 6278 23595
rect 6300 23575 6302 23595
rect 6372 23575 6374 23595
rect 6396 23575 6398 23595
rect 6492 23575 6494 23595
rect 6516 23575 6518 23595
rect 6588 23575 6590 23595
rect 6612 23575 6614 23595
rect 6636 23575 6638 23595
rect 6708 23575 6710 23595
rect 6804 23575 6806 23595
rect 6900 23575 6902 23595
rect 7164 23575 7166 23595
rect 7284 23576 7286 23595
rect 7369 23590 7372 23595
rect 7380 23590 7382 23595
rect 7379 23576 7382 23590
rect 7273 23575 7307 23576
rect 7404 23575 7406 23595
rect 7476 23592 7478 23595
rect 7476 23575 7479 23592
rect 7500 23575 7502 23595
rect 7561 23590 7564 23595
rect 7572 23590 7574 23595
rect 7571 23576 7574 23590
rect 7596 23575 7598 23595
rect 7668 23592 7670 23595
rect 7668 23575 7671 23592
rect 7692 23575 7694 23595
rect 7908 23575 7910 23595
rect 8124 23575 8126 23595
rect 8220 23575 8222 23595
rect 8316 23575 8318 23595
rect 8412 23575 8414 23595
rect 8700 23575 8702 23595
rect 8748 23575 8750 23595
rect 8796 23575 8798 23595
rect 8844 23575 8846 23595
rect 8868 23575 8870 23595
rect 9516 23575 9518 23595
rect 9684 23575 9686 23595
rect 9780 23575 9782 23595
rect 9804 23575 9806 23595
rect 9828 23575 9830 23595
rect 9924 23575 9926 23595
rect 10020 23576 10022 23595
rect 10009 23575 10043 23576
rect 10140 23575 10142 23595
rect 10236 23575 10238 23595
rect 10332 23575 10334 23595
rect 10428 23575 10430 23595
rect 10452 23575 10454 23595
rect 10524 23575 10526 23595
rect 10548 23575 10550 23595
rect 10620 23575 10622 23595
rect 10644 23575 10646 23595
rect 10716 23575 10718 23595
rect 10860 23575 10862 23595
rect 10956 23575 10958 23595
rect 11052 23575 11054 23595
rect 11100 23575 11102 23595
rect 11148 23575 11150 23595
rect 11220 23575 11222 23595
rect 11244 23575 11246 23595
rect 11340 23575 11342 23595
rect 11364 23575 11366 23595
rect 11508 23575 11510 23595
rect 11604 23575 11606 23595
rect 11700 23575 11702 23595
rect 11785 23590 11788 23595
rect 11796 23590 11798 23595
rect 11809 23590 11812 23595
rect 11940 23592 11942 23595
rect 11795 23576 11798 23590
rect 11819 23576 11822 23590
rect 11820 23575 11822 23576
rect 11940 23575 11943 23592
rect 12276 23575 12278 23595
rect 12372 23575 12374 23595
rect 12468 23575 12470 23595
rect 12564 23575 12566 23595
rect 12780 23575 12782 23595
rect 12876 23575 12878 23595
rect 13044 23575 13046 23595
rect 13164 23575 13166 23595
rect 13260 23575 13262 23595
rect 13332 23575 13334 23595
rect 13356 23575 13358 23595
rect 13500 23575 13502 23595
rect 13572 23575 13574 23595
rect 13836 23575 13838 23595
rect 13932 23575 13934 23595
rect 14004 23575 14006 23595
rect 14028 23575 14030 23595
rect 14172 23575 14174 23595
rect 14940 23575 14942 23595
rect 15036 23575 15038 23595
rect 15276 23575 15278 23595
rect 15372 23575 15374 23595
rect 15468 23575 15470 23595
rect 15564 23575 15566 23595
rect 15660 23575 15662 23595
rect 15684 23575 15686 23595
rect 15732 23575 15734 23595
rect 15756 23575 15758 23595
rect 15780 23575 15782 23595
rect 15828 23575 15830 23595
rect 15852 23575 15854 23595
rect 15876 23575 15878 23595
rect 15948 23575 15950 23595
rect 15972 23575 15974 23595
rect 16044 23575 16046 23595
rect 16068 23575 16070 23595
rect 16164 23575 16166 23595
rect 16260 23575 16262 23595
rect 16284 23575 16286 23595
rect 16380 23575 16382 23595
rect 16476 23575 16478 23595
rect 16548 23575 16550 23595
rect 16596 23575 16598 23595
rect 16692 23575 16694 23595
rect 16764 23575 16766 23595
rect 16788 23576 16790 23595
rect 16884 23576 16886 23595
rect 16897 23590 16900 23595
rect 16908 23590 16910 23595
rect 16907 23576 16910 23590
rect 17028 23592 17030 23595
rect 17028 23576 17031 23592
rect 17113 23590 17116 23595
rect 17124 23590 17126 23595
rect 17185 23590 17188 23595
rect 17196 23590 17198 23595
rect 17123 23576 17126 23590
rect 17195 23576 17198 23590
rect 17209 23582 17213 23590
rect 17199 23576 17209 23582
rect 16777 23575 16835 23576
rect 16873 23575 16907 23576
rect 1561 23571 11909 23575
rect 1561 23568 1565 23571
rect 1572 23568 1575 23571
rect 1668 23568 1670 23571
rect 1668 23552 1671 23568
rect 1764 23552 1766 23571
rect 1657 23551 1691 23552
rect 1705 23551 1739 23552
rect 1657 23547 1739 23551
rect 1753 23551 1787 23552
rect 1860 23551 1862 23571
rect 1956 23551 1958 23571
rect 2052 23551 2054 23571
rect 2148 23551 2150 23571
rect 2244 23551 2246 23571
rect 2340 23551 2342 23571
rect 2436 23551 2438 23571
rect 2532 23551 2534 23571
rect 2628 23551 2630 23571
rect 2724 23551 2726 23571
rect 2820 23551 2822 23571
rect 2916 23551 2918 23571
rect 2988 23551 2990 23571
rect 3084 23551 3086 23571
rect 3324 23551 3326 23571
rect 3540 23551 3542 23571
rect 3780 23551 3782 23571
rect 4068 23551 4070 23571
rect 4164 23551 4166 23571
rect 4308 23551 4310 23571
rect 4932 23551 4934 23571
rect 5028 23551 5030 23571
rect 5124 23551 5126 23571
rect 5148 23551 5150 23571
rect 5196 23551 5198 23571
rect 5244 23551 5246 23571
rect 5292 23551 5294 23571
rect 5460 23551 5462 23571
rect 5508 23551 5510 23571
rect 5556 23551 5558 23571
rect 5652 23551 5654 23571
rect 5748 23551 5750 23571
rect 5772 23551 5774 23571
rect 5844 23551 5846 23571
rect 6276 23551 6278 23571
rect 6300 23551 6302 23571
rect 6372 23551 6374 23571
rect 6396 23551 6398 23571
rect 6492 23551 6494 23571
rect 6516 23551 6518 23571
rect 6588 23551 6590 23571
rect 6612 23551 6614 23571
rect 6636 23551 6638 23571
rect 6708 23551 6710 23571
rect 6804 23551 6806 23571
rect 6900 23551 6902 23571
rect 7164 23551 7166 23571
rect 7273 23566 7276 23571
rect 7284 23566 7286 23571
rect 7283 23552 7286 23566
rect 7404 23551 7406 23571
rect 7455 23568 7469 23571
rect 7476 23568 7479 23571
rect 7500 23551 7502 23571
rect 7596 23551 7598 23571
rect 7647 23568 7661 23571
rect 7668 23568 7671 23571
rect 7692 23551 7694 23571
rect 7908 23551 7910 23571
rect 8124 23551 8126 23571
rect 8220 23551 8222 23571
rect 8316 23551 8318 23571
rect 8412 23551 8414 23571
rect 8700 23551 8702 23571
rect 8748 23551 8750 23571
rect 8796 23551 8798 23571
rect 8844 23551 8846 23571
rect 8868 23551 8870 23571
rect 9516 23551 9518 23571
rect 9684 23551 9686 23571
rect 9780 23551 9782 23571
rect 9804 23551 9806 23571
rect 9828 23551 9830 23571
rect 9924 23551 9926 23571
rect 10009 23566 10012 23571
rect 10020 23566 10022 23571
rect 10019 23552 10022 23566
rect 10140 23551 10142 23571
rect 10236 23551 10238 23571
rect 10332 23551 10334 23571
rect 10428 23551 10430 23571
rect 10452 23551 10454 23571
rect 10524 23551 10526 23571
rect 10548 23551 10550 23571
rect 10620 23551 10622 23571
rect 10644 23551 10646 23571
rect 10716 23551 10718 23571
rect 10860 23551 10862 23571
rect 10956 23551 10958 23571
rect 11052 23551 11054 23571
rect 11100 23551 11102 23571
rect 11148 23551 11150 23571
rect 11220 23551 11222 23571
rect 11244 23551 11246 23571
rect 11340 23551 11342 23571
rect 11364 23551 11366 23571
rect 11508 23551 11510 23571
rect 11604 23551 11606 23571
rect 11700 23551 11702 23571
rect 11820 23551 11822 23571
rect 11871 23568 11885 23571
rect 11895 23568 11909 23571
rect 11919 23571 16907 23575
rect 17017 23575 17051 23576
rect 17089 23575 17123 23576
rect 17017 23571 17123 23575
rect 11919 23568 11933 23571
rect 11940 23568 11943 23571
rect 12276 23551 12278 23571
rect 12372 23551 12374 23571
rect 12468 23551 12470 23571
rect 12564 23551 12566 23571
rect 12780 23551 12782 23571
rect 12876 23551 12878 23571
rect 13044 23551 13046 23571
rect 13164 23551 13166 23571
rect 13260 23551 13262 23571
rect 13332 23551 13334 23571
rect 13356 23551 13358 23571
rect 13500 23551 13502 23571
rect 13572 23551 13574 23571
rect 13836 23551 13838 23571
rect 13932 23551 13934 23571
rect 14004 23551 14006 23571
rect 14028 23551 14030 23571
rect 14172 23551 14174 23571
rect 14940 23551 14942 23571
rect 15036 23551 15038 23571
rect 15276 23551 15278 23571
rect 15372 23551 15374 23571
rect 15468 23551 15470 23571
rect 15564 23551 15566 23571
rect 15660 23551 15662 23571
rect 15684 23551 15686 23571
rect 15732 23551 15734 23571
rect 15756 23551 15758 23571
rect 15780 23551 15782 23571
rect 15828 23551 15830 23571
rect 15852 23551 15854 23571
rect 15876 23551 15878 23571
rect 15948 23551 15950 23571
rect 15972 23551 15974 23571
rect 16044 23551 16046 23571
rect 16068 23551 16070 23571
rect 16164 23551 16166 23571
rect 16260 23551 16262 23571
rect 16284 23551 16286 23571
rect 16380 23551 16382 23571
rect 16476 23551 16478 23571
rect 16548 23551 16550 23571
rect 16596 23551 16598 23571
rect 16692 23551 16694 23571
rect 16764 23552 16766 23571
rect 16777 23566 16780 23571
rect 16788 23566 16790 23571
rect 16873 23566 16876 23571
rect 16884 23568 16886 23571
rect 17017 23568 17021 23571
rect 17028 23568 17031 23571
rect 16884 23566 16887 23568
rect 16787 23552 16790 23566
rect 16883 23558 16887 23566
rect 16897 23558 16901 23566
rect 17113 23558 17117 23566
rect 16883 23552 16897 23558
rect 17103 23552 17113 23558
rect 16753 23551 16787 23552
rect 1753 23547 16787 23551
rect 1657 23544 1661 23547
rect 1668 23544 1671 23547
rect 1753 23542 1756 23547
rect 1764 23544 1766 23547
rect 1860 23544 1862 23547
rect 1764 23542 1767 23544
rect 1763 23528 1767 23542
rect 1860 23528 1863 23544
rect 1849 23527 1883 23528
rect 1956 23527 1958 23547
rect 2052 23527 2054 23547
rect 2148 23527 2150 23547
rect 2175 23544 2189 23547
rect 2244 23527 2246 23547
rect 2340 23527 2342 23547
rect 2436 23527 2438 23547
rect 2532 23527 2534 23547
rect 2628 23527 2630 23547
rect 2724 23527 2726 23547
rect 2820 23527 2822 23547
rect 2916 23527 2918 23547
rect 2988 23527 2990 23547
rect 3084 23527 3086 23547
rect 3324 23527 3326 23547
rect 3540 23527 3542 23547
rect 3780 23527 3782 23547
rect 4068 23527 4070 23547
rect 4095 23544 4109 23547
rect 4164 23527 4166 23547
rect 4308 23527 4310 23547
rect 4932 23527 4934 23547
rect 5028 23527 5030 23547
rect 5124 23527 5126 23547
rect 5148 23527 5150 23547
rect 5196 23527 5198 23547
rect 5244 23527 5246 23547
rect 5292 23527 5294 23547
rect 5460 23527 5462 23547
rect 5508 23527 5510 23547
rect 5556 23527 5558 23547
rect 5652 23527 5654 23547
rect 5748 23527 5750 23547
rect 5772 23527 5774 23547
rect 5844 23527 5846 23547
rect 6231 23544 6245 23547
rect 6276 23527 6278 23547
rect 6300 23527 6302 23547
rect 6372 23527 6374 23547
rect 6396 23527 6398 23547
rect 6492 23527 6494 23547
rect 6516 23527 6518 23547
rect 6588 23527 6590 23547
rect 6612 23527 6614 23547
rect 6636 23527 6638 23547
rect 6708 23527 6710 23547
rect 6804 23527 6806 23547
rect 6900 23527 6902 23547
rect 7164 23527 7166 23547
rect 7359 23544 7373 23547
rect 7404 23527 7406 23547
rect 7500 23527 7502 23547
rect 7596 23527 7598 23547
rect 7692 23527 7694 23547
rect 7908 23527 7910 23547
rect 8124 23527 8126 23547
rect 8220 23527 8222 23547
rect 8316 23527 8318 23547
rect 8412 23527 8414 23547
rect 8700 23527 8702 23547
rect 8748 23527 8750 23547
rect 8796 23527 8798 23547
rect 8844 23527 8846 23547
rect 8868 23527 8870 23547
rect 9516 23527 9518 23547
rect 9684 23527 9686 23547
rect 9780 23527 9782 23547
rect 9804 23527 9806 23547
rect 9828 23527 9830 23547
rect 9924 23527 9926 23547
rect 10095 23544 10109 23547
rect 10140 23527 10142 23547
rect 10236 23527 10238 23547
rect 10332 23527 10334 23547
rect 10428 23527 10430 23547
rect 10452 23527 10454 23547
rect 10524 23527 10526 23547
rect 10548 23527 10550 23547
rect 10620 23527 10622 23547
rect 10644 23527 10646 23547
rect 10716 23527 10718 23547
rect 10860 23527 10862 23547
rect 10956 23527 10958 23547
rect 11052 23527 11054 23547
rect 11100 23527 11102 23547
rect 11148 23527 11150 23547
rect 11220 23527 11222 23547
rect 11244 23527 11246 23547
rect 11340 23527 11342 23547
rect 11364 23527 11366 23547
rect 11508 23527 11510 23547
rect 11604 23527 11606 23547
rect 11700 23527 11702 23547
rect 11820 23527 11822 23547
rect 12276 23527 12278 23547
rect 12372 23527 12374 23547
rect 12468 23527 12470 23547
rect 12564 23527 12566 23547
rect 12780 23527 12782 23547
rect 12876 23527 12878 23547
rect 13044 23527 13046 23547
rect 13164 23527 13166 23547
rect 13260 23527 13262 23547
rect 13332 23527 13334 23547
rect 13356 23527 13358 23547
rect 13500 23527 13502 23547
rect 13572 23527 13574 23547
rect 13836 23527 13838 23547
rect 13932 23527 13934 23547
rect 14004 23527 14006 23547
rect 14028 23527 14030 23547
rect 14172 23527 14174 23547
rect 14940 23527 14942 23547
rect 15036 23527 15038 23547
rect 15276 23527 15278 23547
rect 15372 23527 15374 23547
rect 15468 23527 15470 23547
rect 15564 23527 15566 23547
rect 15660 23527 15662 23547
rect 15684 23527 15686 23547
rect 15732 23527 15734 23547
rect 15756 23527 15758 23547
rect 15780 23527 15782 23547
rect 15828 23527 15830 23547
rect 15852 23527 15854 23547
rect 15876 23527 15878 23547
rect 15948 23527 15950 23547
rect 15972 23527 15974 23547
rect 16044 23527 16046 23547
rect 16068 23527 16070 23547
rect 16164 23527 16166 23547
rect 16260 23527 16262 23547
rect 16284 23527 16286 23547
rect 16380 23527 16382 23547
rect 16476 23528 16478 23547
rect 16548 23528 16550 23547
rect 16596 23528 16598 23547
rect 16692 23528 16694 23547
rect 16753 23542 16756 23547
rect 16764 23542 16766 23547
rect 16763 23528 16766 23542
rect 16465 23527 16523 23528
rect 16537 23527 16571 23528
rect 1849 23523 16571 23527
rect 16585 23527 16619 23528
rect 16657 23527 16715 23528
rect 16729 23527 16763 23528
rect 16585 23523 16763 23527
rect 1849 23520 1853 23523
rect 1860 23520 1863 23523
rect 1956 23520 1958 23523
rect 1956 23504 1959 23520
rect 1945 23503 1979 23504
rect 2052 23503 2054 23523
rect 2148 23503 2150 23523
rect 2244 23503 2246 23523
rect 2340 23503 2342 23523
rect 2436 23503 2438 23523
rect 2532 23503 2534 23523
rect 2628 23503 2630 23523
rect 2724 23503 2726 23523
rect 2820 23503 2822 23523
rect 2916 23503 2918 23523
rect 2988 23503 2990 23523
rect 3084 23503 3086 23523
rect 3324 23503 3326 23523
rect 3540 23503 3542 23523
rect 3780 23503 3782 23523
rect 4068 23503 4070 23523
rect 4164 23503 4166 23523
rect 4308 23503 4310 23523
rect 4932 23503 4934 23523
rect 5028 23503 5030 23523
rect 5124 23503 5126 23523
rect 5148 23503 5150 23523
rect 5196 23503 5198 23523
rect 5244 23503 5246 23523
rect 5292 23503 5294 23523
rect 5460 23503 5462 23523
rect 5508 23503 5510 23523
rect 5556 23503 5558 23523
rect 5652 23503 5654 23523
rect 5748 23503 5750 23523
rect 5772 23503 5774 23523
rect 5844 23503 5846 23523
rect 6276 23503 6278 23523
rect 6300 23503 6302 23523
rect 6372 23503 6374 23523
rect 6396 23503 6398 23523
rect 6492 23503 6494 23523
rect 6516 23503 6518 23523
rect 6588 23503 6590 23523
rect 6612 23503 6614 23523
rect 6636 23503 6638 23523
rect 6708 23503 6710 23523
rect 6804 23503 6806 23523
rect 6900 23503 6902 23523
rect 7164 23503 7166 23523
rect 7404 23503 7406 23523
rect 7500 23503 7502 23523
rect 7596 23503 7598 23523
rect 7692 23503 7694 23523
rect 7908 23503 7910 23523
rect 8124 23503 8126 23523
rect 8220 23503 8222 23523
rect 8316 23503 8318 23523
rect 8412 23503 8414 23523
rect 8700 23503 8702 23523
rect 8748 23503 8750 23523
rect 8796 23503 8798 23523
rect 8844 23503 8846 23523
rect 8868 23503 8870 23523
rect 9516 23503 9518 23523
rect 9625 23503 9683 23504
rect 9684 23503 9686 23523
rect 9780 23503 9782 23523
rect 9804 23503 9806 23523
rect 9828 23503 9830 23523
rect 9924 23503 9926 23523
rect 10140 23503 10142 23523
rect 10236 23503 10238 23523
rect 10332 23503 10334 23523
rect 10428 23503 10430 23523
rect 10452 23503 10454 23523
rect 10524 23503 10526 23523
rect 10548 23503 10550 23523
rect 10620 23503 10622 23523
rect 10644 23503 10646 23523
rect 10716 23503 10718 23523
rect 10860 23503 10862 23523
rect 10956 23503 10958 23523
rect 11052 23503 11054 23523
rect 11100 23503 11102 23523
rect 11148 23503 11150 23523
rect 11220 23503 11222 23523
rect 11244 23503 11246 23523
rect 11340 23503 11342 23523
rect 11364 23503 11366 23523
rect 11508 23503 11510 23523
rect 11604 23503 11606 23523
rect 11700 23503 11702 23523
rect 11820 23503 11822 23523
rect 12276 23503 12278 23523
rect 12372 23503 12374 23523
rect 12468 23503 12470 23523
rect 12564 23503 12566 23523
rect 12780 23503 12782 23523
rect 12876 23503 12878 23523
rect 13044 23503 13046 23523
rect 13164 23503 13166 23523
rect 13260 23503 13262 23523
rect 13332 23503 13334 23523
rect 13356 23503 13358 23523
rect 13500 23503 13502 23523
rect 13572 23503 13574 23523
rect 13836 23503 13838 23523
rect 13932 23503 13934 23523
rect 14004 23503 14006 23523
rect 14028 23503 14030 23523
rect 14172 23503 14174 23523
rect 14940 23504 14942 23523
rect 15036 23504 15038 23523
rect 14833 23503 14867 23504
rect 1945 23499 14867 23503
rect 14929 23503 14963 23504
rect 15025 23503 15083 23504
rect 15276 23503 15278 23523
rect 15372 23503 15374 23523
rect 15468 23503 15470 23523
rect 15564 23503 15566 23523
rect 15660 23503 15662 23523
rect 15684 23503 15686 23523
rect 15732 23503 15734 23523
rect 15756 23504 15758 23523
rect 15745 23503 15779 23504
rect 15780 23503 15782 23523
rect 15828 23503 15830 23523
rect 15852 23504 15854 23523
rect 15876 23504 15878 23523
rect 15948 23504 15950 23523
rect 15972 23504 15974 23523
rect 16044 23504 16046 23523
rect 16068 23504 16070 23523
rect 16164 23504 16166 23523
rect 16260 23504 16262 23523
rect 16284 23504 16286 23523
rect 16380 23504 16382 23523
rect 16465 23518 16468 23523
rect 16476 23518 16478 23523
rect 16537 23518 16540 23523
rect 16548 23518 16550 23523
rect 16585 23518 16588 23523
rect 16596 23520 16598 23523
rect 16596 23518 16599 23520
rect 16475 23504 16478 23518
rect 16547 23504 16550 23518
rect 16561 23510 16565 23518
rect 16551 23504 16561 23510
rect 16595 23504 16599 23518
rect 16681 23518 16684 23523
rect 16692 23520 16694 23523
rect 16692 23518 16695 23520
rect 16681 23510 16685 23518
rect 16671 23504 16681 23510
rect 16691 23504 16695 23518
rect 16753 23510 16757 23518
rect 16743 23504 16753 23510
rect 15841 23503 15899 23504
rect 15937 23503 15995 23504
rect 16033 23503 16091 23504
rect 16153 23503 16211 23504
rect 16249 23503 16307 23504
rect 16321 23503 16355 23504
rect 14929 23499 16355 23503
rect 16369 23503 16403 23504
rect 16441 23503 16475 23504
rect 16369 23499 16475 23503
rect 1945 23496 1949 23499
rect 1956 23496 1959 23499
rect 2052 23496 2054 23499
rect 2052 23480 2055 23496
rect 2148 23480 2150 23499
rect 2041 23479 2075 23480
rect 2113 23479 2171 23480
rect 2244 23479 2246 23499
rect 2340 23479 2342 23499
rect 2436 23479 2438 23499
rect 2532 23479 2534 23499
rect 2628 23479 2630 23499
rect 2724 23479 2726 23499
rect 2820 23479 2822 23499
rect 2916 23479 2918 23499
rect 2988 23479 2990 23499
rect 3084 23479 3086 23499
rect 3324 23479 3326 23499
rect 3540 23479 3542 23499
rect 3780 23479 3782 23499
rect 4068 23479 4070 23499
rect 4164 23479 4166 23499
rect 4308 23479 4310 23499
rect 4932 23479 4934 23499
rect 5028 23479 5030 23499
rect 5124 23479 5126 23499
rect 5148 23479 5150 23499
rect 5196 23479 5198 23499
rect 5244 23479 5246 23499
rect 5292 23479 5294 23499
rect 5460 23479 5462 23499
rect 5508 23479 5510 23499
rect 5556 23479 5558 23499
rect 5652 23479 5654 23499
rect 5748 23479 5750 23499
rect 5772 23479 5774 23499
rect 5844 23479 5846 23499
rect 6276 23479 6278 23499
rect 6300 23479 6302 23499
rect 6372 23479 6374 23499
rect 6396 23479 6398 23499
rect 6492 23479 6494 23499
rect 6516 23479 6518 23499
rect 6588 23479 6590 23499
rect 6612 23479 6614 23499
rect 6636 23479 6638 23499
rect 6708 23479 6710 23499
rect 6804 23479 6806 23499
rect 6900 23479 6902 23499
rect 7164 23479 7166 23499
rect 7404 23479 7406 23499
rect 7500 23479 7502 23499
rect 7596 23479 7598 23499
rect 7692 23479 7694 23499
rect 7908 23479 7910 23499
rect 8124 23479 8126 23499
rect 8220 23479 8222 23499
rect 8316 23479 8318 23499
rect 8412 23479 8414 23499
rect 8700 23479 8702 23499
rect 8748 23479 8750 23499
rect 8796 23479 8798 23499
rect 8844 23479 8846 23499
rect 8868 23479 8870 23499
rect 9516 23479 9518 23499
rect 9684 23479 9686 23499
rect 9732 23479 9735 23496
rect 9780 23479 9782 23499
rect 9804 23479 9806 23499
rect 9828 23479 9830 23499
rect 9924 23479 9926 23499
rect 10140 23479 10142 23499
rect 10236 23479 10238 23499
rect 10332 23479 10334 23499
rect 10428 23479 10430 23499
rect 10452 23479 10454 23499
rect 10524 23479 10526 23499
rect 10548 23479 10550 23499
rect 10620 23479 10622 23499
rect 10644 23479 10646 23499
rect 10716 23479 10718 23499
rect 10860 23479 10862 23499
rect 10956 23479 10958 23499
rect 11052 23479 11054 23499
rect 11100 23479 11102 23499
rect 11148 23479 11150 23499
rect 11220 23479 11222 23499
rect 11244 23479 11246 23499
rect 11340 23479 11342 23499
rect 11364 23480 11366 23499
rect 11353 23479 11387 23480
rect 2041 23475 9725 23479
rect 2041 23472 2045 23475
rect 2052 23472 2055 23475
rect 2137 23470 2140 23475
rect 2148 23472 2150 23475
rect 2244 23472 2246 23475
rect 2148 23470 2151 23472
rect 2137 23462 2141 23470
rect 2127 23456 2137 23462
rect 2147 23456 2151 23470
rect 2244 23456 2247 23472
rect 2233 23455 2267 23456
rect 2340 23455 2342 23475
rect 2436 23455 2438 23475
rect 2532 23455 2534 23475
rect 2628 23455 2630 23475
rect 2724 23455 2726 23475
rect 2820 23455 2822 23475
rect 2916 23455 2918 23475
rect 2988 23455 2990 23475
rect 3084 23455 3086 23475
rect 3324 23455 3326 23475
rect 3540 23455 3542 23475
rect 3780 23455 3782 23475
rect 4068 23455 4070 23475
rect 4164 23455 4166 23475
rect 4308 23455 4310 23475
rect 4932 23455 4934 23475
rect 5028 23455 5030 23475
rect 5124 23455 5126 23475
rect 5148 23455 5150 23475
rect 5196 23455 5198 23475
rect 5244 23455 5246 23475
rect 5292 23455 5294 23475
rect 5460 23455 5462 23475
rect 5508 23455 5510 23475
rect 5556 23455 5558 23475
rect 5652 23455 5654 23475
rect 5748 23455 5750 23475
rect 5772 23455 5774 23475
rect 5844 23455 5846 23475
rect 6097 23455 6155 23456
rect 6276 23455 6278 23475
rect 6300 23455 6302 23475
rect 6372 23455 6374 23475
rect 6396 23455 6398 23475
rect 6492 23455 6494 23475
rect 6516 23455 6518 23475
rect 6588 23455 6590 23475
rect 6612 23455 6614 23475
rect 6636 23455 6638 23475
rect 6708 23455 6710 23475
rect 6804 23455 6806 23475
rect 6900 23455 6902 23475
rect 7164 23455 7166 23475
rect 7404 23455 7406 23475
rect 7500 23455 7502 23475
rect 7596 23455 7598 23475
rect 7692 23455 7694 23475
rect 7908 23455 7910 23475
rect 8124 23455 8126 23475
rect 8220 23455 8222 23475
rect 8316 23455 8318 23475
rect 8412 23455 8414 23475
rect 8700 23455 8702 23475
rect 8748 23455 8750 23475
rect 8796 23455 8798 23475
rect 8844 23455 8846 23475
rect 8868 23455 8870 23475
rect 9516 23455 9518 23475
rect 9684 23455 9686 23475
rect 9711 23472 9725 23475
rect 9732 23475 11387 23479
rect 11401 23479 11435 23480
rect 11508 23479 11510 23499
rect 11604 23479 11606 23499
rect 11700 23480 11702 23499
rect 11689 23479 11747 23480
rect 11820 23479 11822 23499
rect 12276 23479 12278 23499
rect 12372 23479 12374 23499
rect 12468 23479 12470 23499
rect 12564 23479 12566 23499
rect 12780 23479 12782 23499
rect 12876 23479 12878 23499
rect 13044 23479 13046 23499
rect 13164 23479 13166 23499
rect 13260 23479 13262 23499
rect 13332 23479 13334 23499
rect 13356 23479 13358 23499
rect 13500 23479 13502 23499
rect 13572 23479 13574 23499
rect 13836 23479 13838 23499
rect 13932 23479 13934 23499
rect 14004 23479 14006 23499
rect 14028 23479 14030 23499
rect 14172 23479 14174 23499
rect 14929 23494 14932 23499
rect 14940 23496 14942 23499
rect 14940 23494 14943 23496
rect 15025 23494 15028 23499
rect 15036 23496 15038 23499
rect 15036 23494 15039 23496
rect 14939 23480 14943 23494
rect 15035 23480 15039 23494
rect 14425 23479 14459 23480
rect 11401 23475 14459 23479
rect 15169 23479 15203 23480
rect 15276 23479 15278 23499
rect 15372 23479 15374 23499
rect 15468 23479 15470 23499
rect 15564 23479 15566 23499
rect 15660 23480 15662 23499
rect 15684 23480 15686 23499
rect 15732 23480 15734 23499
rect 15745 23494 15748 23499
rect 15756 23494 15758 23499
rect 15755 23480 15758 23494
rect 15780 23480 15782 23499
rect 15828 23480 15830 23499
rect 15841 23494 15844 23499
rect 15852 23496 15854 23499
rect 15852 23494 15855 23496
rect 15865 23494 15868 23499
rect 15876 23494 15878 23499
rect 15937 23494 15940 23499
rect 15948 23496 15950 23499
rect 15948 23494 15951 23496
rect 15851 23480 15855 23494
rect 15875 23480 15878 23494
rect 15947 23486 15951 23494
rect 15961 23494 15964 23499
rect 15972 23496 15974 23499
rect 15972 23494 15975 23496
rect 16033 23494 16036 23499
rect 16044 23496 16046 23499
rect 16044 23494 16047 23496
rect 15961 23486 15965 23494
rect 15947 23480 15961 23486
rect 15971 23480 15975 23494
rect 16043 23486 16047 23494
rect 16057 23494 16060 23499
rect 16068 23496 16070 23499
rect 16068 23494 16071 23496
rect 16153 23494 16156 23499
rect 16164 23496 16166 23499
rect 16164 23494 16167 23496
rect 16249 23494 16252 23499
rect 16260 23496 16262 23499
rect 16260 23494 16263 23496
rect 16057 23486 16061 23494
rect 16043 23480 16057 23486
rect 16067 23480 16071 23494
rect 16163 23480 16167 23494
rect 16259 23486 16263 23494
rect 16273 23494 16276 23499
rect 16284 23496 16286 23499
rect 16284 23494 16287 23496
rect 16369 23494 16372 23499
rect 16380 23496 16382 23499
rect 16380 23494 16383 23496
rect 16273 23486 16277 23494
rect 16259 23480 16273 23486
rect 16283 23480 16287 23494
rect 16345 23486 16349 23494
rect 16335 23480 16345 23486
rect 16379 23480 16383 23494
rect 16465 23486 16469 23494
rect 16455 23480 16465 23486
rect 15649 23479 15707 23480
rect 15721 23479 15755 23480
rect 15169 23475 15755 23479
rect 15769 23479 15803 23480
rect 15817 23479 15851 23480
rect 15769 23475 15851 23479
rect 9732 23472 9749 23475
rect 9732 23455 9734 23472
rect 9780 23455 9782 23475
rect 9804 23455 9806 23475
rect 9828 23455 9830 23475
rect 9924 23455 9926 23475
rect 10140 23455 10142 23475
rect 10236 23455 10238 23475
rect 10332 23455 10334 23475
rect 10428 23455 10430 23475
rect 10452 23455 10454 23475
rect 10524 23455 10526 23475
rect 10548 23455 10550 23475
rect 10620 23455 10622 23475
rect 10644 23455 10646 23475
rect 10716 23455 10718 23475
rect 10860 23455 10862 23475
rect 10956 23455 10958 23475
rect 11052 23455 11054 23475
rect 11100 23455 11102 23475
rect 11148 23455 11150 23475
rect 11220 23455 11222 23475
rect 11244 23456 11246 23475
rect 11340 23456 11342 23475
rect 11353 23470 11356 23475
rect 11364 23470 11366 23475
rect 11363 23456 11366 23470
rect 11508 23472 11510 23475
rect 11508 23456 11511 23472
rect 11604 23456 11606 23475
rect 11689 23470 11692 23475
rect 11700 23470 11702 23475
rect 11699 23456 11702 23470
rect 11820 23472 11822 23475
rect 11820 23456 11823 23472
rect 11233 23455 11291 23456
rect 11329 23455 11363 23456
rect 2233 23451 11363 23455
rect 11497 23455 11531 23456
rect 11545 23455 11579 23456
rect 11497 23451 11579 23455
rect 11593 23455 11627 23456
rect 11665 23455 11699 23456
rect 11593 23451 11699 23455
rect 11809 23455 11843 23456
rect 12001 23455 12035 23456
rect 11809 23451 12035 23455
rect 12049 23455 12083 23456
rect 12276 23455 12278 23475
rect 12372 23455 12374 23475
rect 12468 23455 12470 23475
rect 12564 23455 12566 23475
rect 12780 23455 12782 23475
rect 12876 23455 12878 23475
rect 13044 23455 13046 23475
rect 13164 23455 13166 23475
rect 13260 23455 13262 23475
rect 13332 23455 13334 23475
rect 13356 23455 13358 23475
rect 13500 23455 13502 23475
rect 13572 23455 13574 23475
rect 13836 23455 13838 23475
rect 13932 23455 13934 23475
rect 14004 23455 14006 23475
rect 14028 23456 14030 23475
rect 14017 23455 14051 23456
rect 12049 23451 14051 23455
rect 14065 23455 14099 23456
rect 14172 23455 14174 23475
rect 15276 23472 15278 23475
rect 15276 23456 15279 23472
rect 15372 23456 15374 23475
rect 15468 23456 15470 23475
rect 15564 23456 15566 23475
rect 15649 23470 15652 23475
rect 15660 23470 15662 23475
rect 15673 23470 15676 23475
rect 15684 23470 15686 23475
rect 15721 23470 15724 23475
rect 15732 23470 15734 23475
rect 15769 23470 15772 23475
rect 15780 23472 15782 23475
rect 15780 23470 15783 23472
rect 15817 23470 15820 23475
rect 15828 23472 15830 23475
rect 15831 23472 15845 23475
rect 15828 23470 15831 23472
rect 15659 23456 15662 23470
rect 15683 23456 15686 23470
rect 15731 23456 15734 23470
rect 15745 23462 15749 23470
rect 15735 23456 15745 23462
rect 15779 23456 15783 23470
rect 15827 23456 15831 23470
rect 14281 23455 14315 23456
rect 14065 23451 14315 23455
rect 15265 23455 15299 23456
rect 15313 23455 15347 23456
rect 15265 23451 15347 23455
rect 15361 23455 15395 23456
rect 15433 23455 15491 23456
rect 15553 23455 15611 23456
rect 15625 23455 15659 23456
rect 15361 23451 15659 23455
rect 2233 23448 2237 23451
rect 2244 23448 2247 23451
rect 2340 23448 2342 23451
rect 2340 23432 2343 23448
rect 2329 23431 2363 23432
rect 2436 23431 2438 23451
rect 2532 23431 2534 23451
rect 2628 23431 2630 23451
rect 2724 23431 2726 23451
rect 2820 23431 2822 23451
rect 2916 23431 2918 23451
rect 2988 23431 2990 23451
rect 3084 23431 3086 23451
rect 3324 23431 3326 23451
rect 3540 23431 3542 23451
rect 3780 23431 3782 23451
rect 4068 23431 4070 23451
rect 4164 23431 4166 23451
rect 4308 23431 4310 23451
rect 4932 23431 4934 23451
rect 5028 23431 5030 23451
rect 5124 23431 5126 23451
rect 5148 23431 5150 23451
rect 5196 23431 5198 23451
rect 5244 23431 5246 23451
rect 5292 23431 5294 23451
rect 5460 23431 5462 23451
rect 5508 23431 5510 23451
rect 5556 23431 5558 23451
rect 5652 23431 5654 23451
rect 5748 23431 5750 23451
rect 5772 23431 5774 23451
rect 5844 23431 5846 23451
rect 6097 23446 6100 23451
rect 6107 23432 6110 23446
rect 6108 23431 6110 23432
rect 6204 23431 6207 23448
rect 6276 23431 6278 23451
rect 6300 23431 6302 23451
rect 6372 23431 6374 23451
rect 6396 23431 6398 23451
rect 6492 23431 6494 23451
rect 6516 23431 6518 23451
rect 6588 23431 6590 23451
rect 6612 23431 6614 23451
rect 6636 23431 6638 23451
rect 6708 23431 6710 23451
rect 6804 23431 6806 23451
rect 6900 23431 6902 23451
rect 7164 23431 7166 23451
rect 7404 23431 7406 23451
rect 7500 23431 7502 23451
rect 7596 23431 7598 23451
rect 7692 23431 7694 23451
rect 7908 23431 7910 23451
rect 8124 23431 8126 23451
rect 8220 23431 8222 23451
rect 8316 23431 8318 23451
rect 8412 23431 8414 23451
rect 8700 23431 8702 23451
rect 8748 23431 8750 23451
rect 8796 23431 8798 23451
rect 8844 23431 8846 23451
rect 8868 23431 8870 23451
rect 9516 23431 9518 23451
rect 9684 23431 9686 23451
rect 9732 23431 9734 23451
rect 9780 23431 9782 23451
rect 9804 23431 9806 23451
rect 9828 23431 9830 23451
rect 9924 23431 9926 23451
rect 10140 23431 10142 23451
rect 10236 23431 10238 23451
rect 10332 23431 10334 23451
rect 10428 23431 10430 23451
rect 10452 23431 10454 23451
rect 10524 23431 10526 23451
rect 10548 23431 10550 23451
rect 10620 23431 10622 23451
rect 10644 23431 10646 23451
rect 10716 23431 10718 23451
rect 10860 23431 10862 23451
rect 10956 23431 10958 23451
rect 11052 23431 11054 23451
rect 11100 23431 11102 23451
rect 11148 23432 11150 23451
rect 11220 23432 11222 23451
rect 11233 23446 11236 23451
rect 11244 23446 11246 23451
rect 11329 23446 11332 23451
rect 11340 23448 11342 23451
rect 11497 23448 11501 23451
rect 11508 23448 11511 23451
rect 11340 23446 11343 23448
rect 11593 23446 11596 23451
rect 11604 23448 11606 23451
rect 11809 23448 11813 23451
rect 11820 23448 11823 23451
rect 11604 23446 11607 23448
rect 11243 23432 11246 23446
rect 11339 23438 11343 23446
rect 11353 23438 11357 23446
rect 11339 23432 11353 23438
rect 11603 23432 11607 23446
rect 11689 23438 11693 23446
rect 11679 23432 11689 23438
rect 12276 23432 12278 23451
rect 12372 23432 12374 23451
rect 11113 23431 11171 23432
rect 11209 23431 11243 23432
rect 2329 23427 6197 23431
rect 2329 23424 2333 23427
rect 2340 23424 2343 23427
rect 2436 23424 2438 23427
rect 2436 23408 2439 23424
rect 2425 23407 2459 23408
rect 2532 23407 2534 23427
rect 2628 23407 2630 23427
rect 2724 23407 2726 23427
rect 2820 23407 2822 23427
rect 2916 23407 2918 23427
rect 2988 23407 2990 23427
rect 3084 23407 3086 23427
rect 3289 23407 3323 23408
rect 3324 23407 3326 23427
rect 3540 23407 3542 23427
rect 3780 23407 3782 23427
rect 4068 23407 4070 23427
rect 4164 23407 4166 23427
rect 4308 23407 4310 23427
rect 4932 23407 4934 23427
rect 5028 23407 5030 23427
rect 5124 23407 5126 23427
rect 5148 23407 5150 23427
rect 5196 23407 5198 23427
rect 5244 23407 5246 23427
rect 5292 23407 5294 23427
rect 5460 23407 5462 23427
rect 5508 23407 5510 23427
rect 5556 23407 5558 23427
rect 5652 23407 5654 23427
rect 5748 23407 5750 23427
rect 5772 23407 5774 23427
rect 5844 23407 5846 23427
rect 6108 23407 6110 23427
rect 6183 23424 6197 23427
rect 6204 23427 11243 23431
rect 11929 23431 11963 23432
rect 11977 23431 12011 23432
rect 11929 23427 12011 23431
rect 12169 23431 12203 23432
rect 12217 23431 12251 23432
rect 12169 23427 12251 23431
rect 12265 23431 12299 23432
rect 12337 23431 12395 23432
rect 12468 23431 12470 23451
rect 12529 23431 12563 23432
rect 12564 23431 12566 23451
rect 12780 23431 12782 23451
rect 12876 23431 12878 23451
rect 12937 23431 12971 23432
rect 13044 23431 13046 23451
rect 13164 23431 13166 23451
rect 13260 23431 13262 23451
rect 13332 23431 13334 23451
rect 13356 23431 13358 23451
rect 13500 23431 13502 23451
rect 13572 23432 13574 23451
rect 13561 23431 13595 23432
rect 12265 23427 13595 23431
rect 13609 23431 13643 23432
rect 13681 23431 13715 23432
rect 13609 23427 13715 23431
rect 13729 23431 13763 23432
rect 13836 23431 13838 23451
rect 13932 23432 13934 23451
rect 14004 23432 14006 23451
rect 14017 23446 14020 23451
rect 14028 23446 14030 23451
rect 14027 23432 14030 23446
rect 14172 23448 14174 23451
rect 15265 23448 15269 23451
rect 15276 23448 15279 23451
rect 14172 23432 14175 23448
rect 15361 23446 15364 23451
rect 15372 23448 15374 23451
rect 15372 23446 15375 23448
rect 15371 23432 15375 23446
rect 15457 23446 15460 23451
rect 15468 23448 15470 23451
rect 15468 23446 15471 23448
rect 15553 23446 15556 23451
rect 15564 23448 15566 23451
rect 15564 23446 15567 23448
rect 15457 23438 15461 23446
rect 15447 23432 15457 23438
rect 15467 23432 15471 23446
rect 15563 23432 15567 23446
rect 15649 23438 15653 23446
rect 15639 23432 15649 23438
rect 13897 23431 13955 23432
rect 13993 23431 14027 23432
rect 13729 23427 14027 23431
rect 14161 23431 14195 23432
rect 14233 23431 14267 23432
rect 14161 23427 14267 23431
rect 6204 23424 6221 23427
rect 6204 23407 6206 23424
rect 6276 23407 6278 23427
rect 6300 23407 6302 23427
rect 6372 23407 6374 23427
rect 6396 23407 6398 23427
rect 6492 23407 6494 23427
rect 6516 23407 6518 23427
rect 6588 23407 6590 23427
rect 6612 23407 6614 23427
rect 6636 23407 6638 23427
rect 6708 23407 6710 23427
rect 6804 23407 6806 23427
rect 6900 23407 6902 23427
rect 7164 23407 7166 23427
rect 7404 23407 7406 23427
rect 7500 23407 7502 23427
rect 7596 23407 7598 23427
rect 7692 23407 7694 23427
rect 7908 23407 7910 23427
rect 8124 23407 8126 23427
rect 8220 23407 8222 23427
rect 8316 23407 8318 23427
rect 8412 23407 8414 23427
rect 8700 23407 8702 23427
rect 8748 23407 8750 23427
rect 8796 23407 8798 23427
rect 8844 23407 8846 23427
rect 8868 23407 8870 23427
rect 9516 23407 9518 23427
rect 9684 23407 9686 23427
rect 9732 23407 9734 23427
rect 9780 23407 9782 23427
rect 9804 23408 9806 23427
rect 9828 23408 9830 23427
rect 9793 23407 9851 23408
rect 9924 23407 9926 23427
rect 10140 23407 10142 23427
rect 10236 23407 10238 23427
rect 10332 23407 10334 23427
rect 10428 23407 10430 23427
rect 10452 23407 10454 23427
rect 10524 23407 10526 23427
rect 10548 23407 10550 23427
rect 10620 23407 10622 23427
rect 10644 23407 10646 23427
rect 10716 23407 10718 23427
rect 10860 23407 10862 23427
rect 10956 23407 10958 23427
rect 11052 23407 11054 23427
rect 11100 23408 11102 23427
rect 11137 23422 11140 23427
rect 11148 23422 11150 23427
rect 11209 23422 11212 23427
rect 11220 23424 11222 23427
rect 11220 23422 11223 23424
rect 12265 23422 12268 23427
rect 12276 23424 12278 23427
rect 12276 23422 12279 23424
rect 11147 23408 11150 23422
rect 11219 23414 11223 23422
rect 11233 23414 11237 23422
rect 11219 23408 11233 23414
rect 12275 23408 12279 23422
rect 12361 23422 12364 23427
rect 12372 23424 12374 23427
rect 12468 23424 12470 23427
rect 12372 23422 12375 23424
rect 12361 23414 12365 23422
rect 12351 23408 12361 23414
rect 12371 23408 12375 23422
rect 12468 23408 12471 23424
rect 11089 23407 11123 23408
rect 2425 23403 11123 23407
rect 12457 23407 12491 23408
rect 12564 23407 12566 23427
rect 12780 23407 12782 23427
rect 12876 23407 12878 23427
rect 13044 23424 13046 23427
rect 13044 23407 13047 23424
rect 13164 23407 13166 23427
rect 13260 23407 13262 23427
rect 13332 23407 13334 23427
rect 13356 23408 13358 23427
rect 13500 23408 13502 23427
rect 13561 23422 13564 23427
rect 13572 23422 13574 23427
rect 13836 23424 13838 23427
rect 13571 23408 13574 23422
rect 13705 23414 13709 23422
rect 13695 23408 13705 23414
rect 13836 23408 13839 23424
rect 13921 23422 13924 23427
rect 13932 23422 13934 23427
rect 13993 23422 13996 23427
rect 14004 23424 14006 23427
rect 14161 23424 14165 23427
rect 14172 23424 14175 23427
rect 14004 23422 14007 23424
rect 13931 23408 13934 23422
rect 14003 23414 14007 23422
rect 14017 23414 14021 23422
rect 14257 23414 14261 23422
rect 14003 23408 14017 23414
rect 14247 23408 14257 23414
rect 13345 23407 13379 23408
rect 12457 23403 13379 23407
rect 13393 23407 13427 23408
rect 13465 23407 13523 23408
rect 13537 23407 13571 23408
rect 13393 23403 13571 23407
rect 13825 23407 13859 23408
rect 13873 23407 13907 23408
rect 13825 23403 13907 23407
rect 2425 23400 2429 23403
rect 2436 23400 2439 23403
rect 2532 23400 2534 23403
rect 2532 23384 2535 23400
rect 2521 23383 2555 23384
rect 2628 23383 2630 23403
rect 2724 23383 2726 23403
rect 2820 23383 2822 23403
rect 2916 23383 2918 23403
rect 2988 23384 2990 23403
rect 2929 23383 2963 23384
rect 2521 23379 2963 23383
rect 2977 23383 3011 23384
rect 3084 23383 3086 23403
rect 3324 23383 3326 23403
rect 3540 23383 3542 23403
rect 3780 23383 3782 23403
rect 4068 23383 4070 23403
rect 4164 23383 4166 23403
rect 4308 23383 4310 23403
rect 4932 23383 4934 23403
rect 5028 23383 5030 23403
rect 5124 23383 5126 23403
rect 5148 23383 5150 23403
rect 5196 23383 5198 23403
rect 5244 23383 5246 23403
rect 5292 23383 5294 23403
rect 5460 23383 5462 23403
rect 5508 23383 5510 23403
rect 5556 23383 5558 23403
rect 5652 23383 5654 23403
rect 5748 23383 5750 23403
rect 5772 23383 5774 23403
rect 5844 23383 5846 23403
rect 6108 23383 6110 23403
rect 6204 23383 6206 23403
rect 6276 23383 6278 23403
rect 6300 23383 6302 23403
rect 6372 23383 6374 23403
rect 6396 23383 6398 23403
rect 6492 23383 6494 23403
rect 6516 23383 6518 23403
rect 6588 23383 6590 23403
rect 6612 23383 6614 23403
rect 6636 23383 6638 23403
rect 6708 23383 6710 23403
rect 6804 23383 6806 23403
rect 6900 23383 6902 23403
rect 7164 23383 7166 23403
rect 7404 23383 7406 23403
rect 7500 23383 7502 23403
rect 7596 23383 7598 23403
rect 7692 23383 7694 23403
rect 7908 23383 7910 23403
rect 8124 23383 8126 23403
rect 8220 23383 8222 23403
rect 8316 23383 8318 23403
rect 8412 23383 8414 23403
rect 8700 23383 8702 23403
rect 8748 23383 8750 23403
rect 8796 23383 8798 23403
rect 8844 23383 8846 23403
rect 8868 23383 8870 23403
rect 9516 23383 9518 23403
rect 9684 23383 9686 23403
rect 9732 23384 9734 23403
rect 9780 23384 9782 23403
rect 9793 23398 9796 23403
rect 9804 23398 9806 23403
rect 9817 23398 9820 23403
rect 9828 23398 9830 23403
rect 9803 23384 9806 23398
rect 9827 23384 9830 23398
rect 9924 23400 9926 23403
rect 9924 23384 9927 23400
rect 9697 23383 9755 23384
rect 9769 23383 9803 23384
rect 2977 23379 9803 23383
rect 9913 23383 9947 23384
rect 10140 23383 10142 23403
rect 10236 23383 10238 23403
rect 10332 23383 10334 23403
rect 10428 23383 10430 23403
rect 10452 23383 10454 23403
rect 10524 23383 10526 23403
rect 10548 23383 10550 23403
rect 10620 23383 10622 23403
rect 10644 23383 10646 23403
rect 10716 23383 10718 23403
rect 10860 23383 10862 23403
rect 10956 23383 10958 23403
rect 11052 23383 11054 23403
rect 11089 23398 11092 23403
rect 11100 23398 11102 23403
rect 12457 23400 12461 23403
rect 12468 23400 12471 23403
rect 12564 23400 12566 23403
rect 12615 23400 12629 23403
rect 11099 23384 11102 23398
rect 12564 23384 12567 23400
rect 11065 23383 11099 23384
rect 9913 23379 11099 23383
rect 12553 23383 12587 23384
rect 12780 23383 12782 23403
rect 12876 23383 12878 23403
rect 13023 23400 13037 23403
rect 13044 23400 13047 23403
rect 13164 23384 13166 23403
rect 13260 23384 13262 23403
rect 13332 23384 13334 23403
rect 13345 23398 13348 23403
rect 13356 23398 13358 23403
rect 13355 23384 13358 23398
rect 13489 23398 13492 23403
rect 13500 23400 13502 23403
rect 13825 23400 13829 23403
rect 13836 23400 13839 23403
rect 13500 23398 13503 23400
rect 13489 23390 13493 23398
rect 13479 23384 13489 23390
rect 13499 23384 13503 23398
rect 13561 23390 13565 23398
rect 13551 23384 13561 23390
rect 13105 23383 13139 23384
rect 12553 23379 13139 23383
rect 13153 23383 13187 23384
rect 13225 23383 13283 23384
rect 13321 23383 13355 23384
rect 13153 23379 13355 23383
rect 2521 23376 2525 23379
rect 2532 23376 2535 23379
rect 2628 23376 2630 23379
rect 2628 23360 2631 23376
rect 2617 23359 2651 23360
rect 2724 23359 2726 23379
rect 2820 23359 2822 23379
rect 2916 23360 2918 23379
rect 2977 23374 2980 23379
rect 2988 23374 2990 23379
rect 2987 23360 2990 23374
rect 3084 23376 3086 23379
rect 3084 23360 3087 23376
rect 2905 23359 2939 23360
rect 2617 23355 2939 23359
rect 3073 23359 3107 23360
rect 3324 23359 3326 23379
rect 3375 23376 3389 23379
rect 3540 23359 3542 23379
rect 3780 23359 3782 23379
rect 4068 23359 4070 23379
rect 4164 23359 4166 23379
rect 4308 23359 4310 23379
rect 4932 23359 4934 23379
rect 5028 23359 5030 23379
rect 5124 23359 5126 23379
rect 5148 23359 5150 23379
rect 5196 23359 5198 23379
rect 5244 23359 5246 23379
rect 5292 23359 5294 23379
rect 5460 23359 5462 23379
rect 5508 23359 5510 23379
rect 5556 23359 5558 23379
rect 5652 23359 5654 23379
rect 5748 23359 5750 23379
rect 5772 23359 5774 23379
rect 5844 23359 5846 23379
rect 6108 23359 6110 23379
rect 6204 23359 6206 23379
rect 6276 23359 6278 23379
rect 6300 23359 6302 23379
rect 6372 23359 6374 23379
rect 6396 23359 6398 23379
rect 6492 23359 6494 23379
rect 6516 23359 6518 23379
rect 6588 23359 6590 23379
rect 6612 23359 6614 23379
rect 6636 23359 6638 23379
rect 6708 23359 6710 23379
rect 6804 23359 6806 23379
rect 6900 23359 6902 23379
rect 7164 23359 7166 23379
rect 7404 23359 7406 23379
rect 7500 23359 7502 23379
rect 7596 23359 7598 23379
rect 7692 23359 7694 23379
rect 7908 23359 7910 23379
rect 8124 23359 8126 23379
rect 8220 23359 8222 23379
rect 8316 23359 8318 23379
rect 8412 23359 8414 23379
rect 8700 23359 8702 23379
rect 8748 23359 8750 23379
rect 8796 23359 8798 23379
rect 8844 23359 8846 23379
rect 8868 23359 8870 23379
rect 9516 23360 9518 23379
rect 9684 23360 9686 23379
rect 9721 23374 9724 23379
rect 9732 23374 9734 23379
rect 9769 23374 9772 23379
rect 9780 23374 9782 23379
rect 9913 23376 9917 23379
rect 9924 23376 9927 23379
rect 9731 23360 9734 23374
rect 9779 23360 9782 23374
rect 9793 23366 9797 23374
rect 9783 23360 9793 23366
rect 9409 23359 9443 23360
rect 3073 23355 9443 23359
rect 9505 23359 9539 23360
rect 9577 23359 9611 23360
rect 9505 23355 9611 23359
rect 9625 23359 9659 23360
rect 9673 23359 9707 23360
rect 9625 23355 9707 23359
rect 10033 23359 10067 23360
rect 10140 23359 10142 23379
rect 10236 23359 10238 23379
rect 10332 23359 10334 23379
rect 10428 23360 10430 23379
rect 10452 23360 10454 23379
rect 10524 23360 10526 23379
rect 10548 23360 10550 23379
rect 10620 23360 10622 23379
rect 10644 23360 10646 23379
rect 10716 23360 10718 23379
rect 10860 23360 10862 23379
rect 10956 23360 10958 23379
rect 11052 23360 11054 23379
rect 12553 23376 12557 23379
rect 12564 23376 12567 23379
rect 12780 23360 12782 23379
rect 12876 23360 12878 23379
rect 13153 23374 13156 23379
rect 13164 23374 13166 23379
rect 13163 23360 13166 23374
rect 13249 23374 13252 23379
rect 13260 23376 13262 23379
rect 13260 23374 13263 23376
rect 13321 23374 13324 23379
rect 13332 23376 13334 23379
rect 13332 23374 13335 23376
rect 13249 23366 13253 23374
rect 13239 23360 13249 23366
rect 13259 23360 13263 23374
rect 13331 23366 13335 23374
rect 13345 23366 13349 23374
rect 13331 23360 13345 23366
rect 10417 23359 10475 23360
rect 10513 23359 10571 23360
rect 10609 23359 10667 23360
rect 10705 23359 10739 23360
rect 10033 23355 10739 23359
rect 10753 23359 10787 23360
rect 10849 23359 10907 23360
rect 10945 23359 10979 23360
rect 10753 23355 10979 23359
rect 10993 23359 11027 23360
rect 11041 23359 11075 23360
rect 10993 23355 11075 23359
rect 12673 23359 12707 23360
rect 12745 23359 12803 23360
rect 12817 23359 12851 23360
rect 12673 23355 12851 23359
rect 12865 23359 12899 23360
rect 13057 23359 13091 23360
rect 12865 23355 13091 23359
rect 2617 23352 2621 23355
rect 2628 23352 2631 23355
rect 2724 23352 2726 23355
rect 2724 23336 2727 23352
rect 2713 23335 2747 23336
rect 2820 23335 2822 23355
rect 2905 23350 2908 23355
rect 2916 23350 2918 23355
rect 3073 23352 3077 23355
rect 3084 23352 3087 23355
rect 2915 23336 2918 23350
rect 2881 23335 2915 23336
rect 2713 23331 2915 23335
rect 3217 23335 3251 23336
rect 3324 23335 3326 23355
rect 3540 23335 3542 23355
rect 3780 23335 3782 23355
rect 4068 23335 4070 23355
rect 4164 23335 4166 23355
rect 4308 23335 4310 23355
rect 4932 23335 4934 23355
rect 5028 23335 5030 23355
rect 5124 23335 5126 23355
rect 5148 23335 5150 23355
rect 5196 23335 5198 23355
rect 5244 23335 5246 23355
rect 5292 23335 5294 23355
rect 5460 23335 5462 23355
rect 5508 23335 5510 23355
rect 5556 23335 5558 23355
rect 5652 23335 5654 23355
rect 5748 23335 5750 23355
rect 5772 23335 5774 23355
rect 5844 23335 5846 23355
rect 6108 23335 6110 23355
rect 6204 23335 6206 23355
rect 6276 23335 6278 23355
rect 6300 23335 6302 23355
rect 6372 23335 6374 23355
rect 6396 23335 6398 23355
rect 6492 23335 6494 23355
rect 6516 23335 6518 23355
rect 6588 23335 6590 23355
rect 6612 23335 6614 23355
rect 6636 23335 6638 23355
rect 6708 23335 6710 23355
rect 6804 23335 6806 23355
rect 6900 23335 6902 23355
rect 7164 23335 7166 23355
rect 7404 23335 7406 23355
rect 7500 23335 7502 23355
rect 7596 23335 7598 23355
rect 7692 23335 7694 23355
rect 7908 23335 7910 23355
rect 8124 23335 8126 23355
rect 8220 23335 8222 23355
rect 8316 23335 8318 23355
rect 8412 23335 8414 23355
rect 8700 23335 8702 23355
rect 8748 23335 8750 23355
rect 8796 23335 8798 23355
rect 8844 23335 8846 23355
rect 8868 23335 8870 23355
rect 9505 23350 9508 23355
rect 9516 23352 9518 23355
rect 9516 23350 9519 23352
rect 9673 23350 9676 23355
rect 9684 23352 9686 23355
rect 10140 23352 10142 23355
rect 9684 23350 9687 23352
rect 9515 23336 9519 23350
rect 9601 23342 9605 23350
rect 9591 23336 9601 23342
rect 9683 23336 9687 23350
rect 10140 23336 10143 23352
rect 9049 23335 9083 23336
rect 3217 23331 9083 23335
rect 10129 23335 10163 23336
rect 10236 23335 10238 23355
rect 10332 23336 10334 23355
rect 10417 23350 10420 23355
rect 10428 23350 10430 23355
rect 10441 23350 10444 23355
rect 10452 23350 10454 23355
rect 10513 23350 10516 23355
rect 10524 23352 10526 23355
rect 10524 23350 10527 23352
rect 10427 23336 10430 23350
rect 10451 23336 10454 23350
rect 10523 23342 10527 23350
rect 10537 23350 10540 23355
rect 10548 23352 10550 23355
rect 10548 23350 10551 23352
rect 10609 23350 10612 23355
rect 10620 23352 10622 23355
rect 10620 23350 10623 23352
rect 10537 23342 10541 23350
rect 10523 23336 10537 23342
rect 10547 23336 10551 23350
rect 10619 23342 10623 23350
rect 10633 23350 10636 23355
rect 10644 23352 10646 23355
rect 10644 23350 10647 23352
rect 10705 23350 10708 23355
rect 10716 23352 10718 23355
rect 10716 23350 10719 23352
rect 10849 23350 10852 23355
rect 10860 23352 10862 23355
rect 10860 23350 10863 23352
rect 10945 23350 10948 23355
rect 10956 23352 10958 23355
rect 10956 23350 10959 23352
rect 11041 23350 11044 23355
rect 11052 23352 11054 23355
rect 11052 23350 11055 23352
rect 10633 23342 10637 23350
rect 10619 23336 10633 23342
rect 10643 23336 10647 23350
rect 10715 23342 10719 23350
rect 10729 23342 10733 23350
rect 10715 23336 10729 23342
rect 10859 23336 10863 23350
rect 10955 23342 10959 23350
rect 10969 23342 10973 23350
rect 10955 23336 10969 23342
rect 11051 23336 11055 23350
rect 12769 23350 12772 23355
rect 12780 23352 12782 23355
rect 12780 23350 12783 23352
rect 12865 23350 12868 23355
rect 12876 23352 12878 23355
rect 12876 23350 12879 23352
rect 12769 23342 12773 23350
rect 12759 23336 12769 23342
rect 12779 23336 12783 23350
rect 12841 23342 12845 23350
rect 12831 23336 12841 23342
rect 12875 23336 12879 23350
rect 10321 23335 10379 23336
rect 10393 23335 10427 23336
rect 10129 23331 10427 23335
rect 12985 23335 13019 23336
rect 13033 23335 13067 23336
rect 12985 23331 13067 23335
rect 2713 23328 2717 23331
rect 2724 23328 2727 23331
rect 2820 23328 2822 23331
rect 3324 23328 3326 23331
rect 2820 23312 2823 23328
rect 3324 23312 3327 23328
rect 3540 23312 3542 23331
rect 2809 23311 2843 23312
rect 2857 23311 2891 23312
rect 2809 23307 2891 23311
rect 3313 23311 3347 23312
rect 3529 23311 3587 23312
rect 3780 23311 3782 23331
rect 4068 23311 4070 23331
rect 4164 23311 4166 23331
rect 4308 23311 4310 23331
rect 4932 23311 4934 23331
rect 5028 23311 5030 23331
rect 5124 23311 5126 23331
rect 5148 23311 5150 23331
rect 5196 23311 5198 23331
rect 5244 23311 5246 23331
rect 5292 23311 5294 23331
rect 5460 23311 5462 23331
rect 5508 23311 5510 23331
rect 5556 23311 5558 23331
rect 5652 23311 5654 23331
rect 5748 23311 5750 23331
rect 5772 23311 5774 23331
rect 5844 23311 5846 23331
rect 6108 23311 6110 23331
rect 6204 23311 6206 23331
rect 6276 23311 6278 23331
rect 6300 23311 6302 23331
rect 6372 23311 6374 23331
rect 6396 23311 6398 23331
rect 6492 23311 6494 23331
rect 6516 23311 6518 23331
rect 6588 23311 6590 23331
rect 6612 23311 6614 23331
rect 6636 23311 6638 23331
rect 6708 23311 6710 23331
rect 6804 23311 6806 23331
rect 6900 23312 6902 23331
rect 6889 23311 6923 23312
rect 3313 23307 6923 23311
rect 6937 23311 6971 23312
rect 7164 23311 7166 23331
rect 7404 23311 7406 23331
rect 7500 23311 7502 23331
rect 7596 23311 7598 23331
rect 7692 23311 7694 23331
rect 7908 23311 7910 23331
rect 8124 23311 8126 23331
rect 8220 23311 8222 23331
rect 8316 23311 8318 23331
rect 8412 23311 8414 23331
rect 8700 23311 8702 23331
rect 8748 23311 8750 23331
rect 8796 23311 8798 23331
rect 8844 23311 8846 23331
rect 8868 23312 8870 23331
rect 10129 23328 10133 23331
rect 10140 23328 10143 23331
rect 10236 23328 10238 23331
rect 10236 23312 10239 23328
rect 10321 23326 10324 23331
rect 10332 23326 10334 23331
rect 10331 23312 10334 23326
rect 10417 23318 10421 23326
rect 10407 23312 10417 23318
rect 8857 23311 8891 23312
rect 6937 23307 8891 23311
rect 10225 23311 10259 23312
rect 10273 23311 10307 23312
rect 10225 23307 10307 23311
rect 2809 23304 2813 23307
rect 2820 23304 2823 23307
rect 3313 23304 3317 23307
rect 3324 23304 3327 23307
rect 3529 23302 3532 23307
rect 3540 23302 3542 23307
rect 3539 23288 3542 23302
rect 3433 23287 3467 23288
rect 3505 23287 3539 23288
rect 3433 23283 3539 23287
rect 3673 23287 3707 23288
rect 3780 23287 3782 23307
rect 4068 23287 4070 23307
rect 4164 23287 4166 23307
rect 4308 23287 4310 23307
rect 4932 23287 4934 23307
rect 5028 23287 5030 23307
rect 5124 23288 5126 23307
rect 5148 23288 5150 23307
rect 5113 23287 5171 23288
rect 5196 23287 5198 23307
rect 5244 23287 5246 23307
rect 5292 23287 5294 23307
rect 5460 23287 5462 23307
rect 5508 23287 5510 23307
rect 5556 23287 5558 23307
rect 5652 23287 5654 23307
rect 5748 23287 5750 23307
rect 5772 23287 5774 23307
rect 5844 23287 5846 23307
rect 6108 23287 6110 23307
rect 6204 23287 6206 23307
rect 6276 23287 6278 23307
rect 6300 23287 6302 23307
rect 6372 23287 6374 23307
rect 6396 23287 6398 23307
rect 6492 23287 6494 23307
rect 6516 23287 6518 23307
rect 6588 23287 6590 23307
rect 6612 23287 6614 23307
rect 6636 23287 6638 23307
rect 6708 23287 6710 23307
rect 6804 23287 6806 23307
rect 6889 23302 6892 23307
rect 6900 23302 6902 23307
rect 6899 23288 6902 23302
rect 7164 23288 7166 23307
rect 6817 23287 6851 23288
rect 3673 23283 6851 23287
rect 7057 23287 7091 23288
rect 7153 23287 7211 23288
rect 7404 23287 7406 23307
rect 7500 23287 7502 23307
rect 7596 23287 7598 23307
rect 7692 23287 7694 23307
rect 7908 23287 7910 23307
rect 8124 23287 8126 23307
rect 8220 23287 8222 23307
rect 8316 23287 8318 23307
rect 8412 23287 8414 23307
rect 8700 23287 8702 23307
rect 8748 23287 8750 23307
rect 8796 23288 8798 23307
rect 8844 23288 8846 23307
rect 8857 23302 8860 23307
rect 8868 23302 8870 23307
rect 10225 23304 10229 23307
rect 10236 23304 10239 23307
rect 8867 23288 8870 23302
rect 8761 23287 8819 23288
rect 8833 23287 8867 23288
rect 7057 23283 8867 23287
rect 3780 23280 3782 23283
rect 3529 23270 3533 23278
rect 3519 23264 3529 23270
rect 3780 23264 3783 23280
rect 3769 23263 3803 23264
rect 4068 23263 4070 23283
rect 4164 23263 4166 23283
rect 4308 23263 4310 23283
rect 4932 23264 4934 23283
rect 5028 23264 5030 23283
rect 5113 23278 5116 23283
rect 5124 23278 5126 23283
rect 5137 23278 5140 23283
rect 5148 23278 5150 23283
rect 5123 23264 5126 23278
rect 5147 23264 5150 23278
rect 5196 23264 5198 23283
rect 5244 23280 5246 23283
rect 4489 23263 4523 23264
rect 4873 23263 4907 23264
rect 3769 23259 4907 23263
rect 4921 23263 4955 23264
rect 5017 23263 5075 23264
rect 5089 23263 5123 23264
rect 4921 23259 5123 23263
rect 5185 23259 5213 23264
rect 5244 23263 5247 23280
rect 5292 23263 5294 23283
rect 5460 23263 5462 23283
rect 5508 23263 5510 23283
rect 5556 23263 5558 23283
rect 5652 23263 5654 23283
rect 5748 23263 5750 23283
rect 5772 23263 5774 23283
rect 5844 23263 5846 23283
rect 6108 23263 6110 23283
rect 6204 23263 6206 23283
rect 6276 23263 6278 23283
rect 6300 23263 6302 23283
rect 6372 23263 6374 23283
rect 6396 23263 6398 23283
rect 6492 23263 6494 23283
rect 6516 23263 6518 23283
rect 6588 23263 6590 23283
rect 6612 23264 6614 23283
rect 6636 23264 6638 23283
rect 6708 23264 6710 23283
rect 6804 23264 6806 23283
rect 7153 23278 7156 23283
rect 7164 23280 7166 23283
rect 7164 23278 7167 23280
rect 7163 23264 7167 23278
rect 7404 23264 7406 23283
rect 7500 23264 7502 23283
rect 6601 23263 6659 23264
rect 6697 23263 6731 23264
rect 3769 23256 3773 23259
rect 3780 23256 3783 23259
rect 3961 23239 3995 23240
rect 4068 23239 4070 23259
rect 4164 23239 4166 23259
rect 4308 23239 4310 23259
rect 4921 23254 4924 23259
rect 4932 23254 4934 23259
rect 5017 23254 5020 23259
rect 5028 23256 5030 23259
rect 5028 23254 5031 23256
rect 5185 23254 5188 23259
rect 5196 23256 5198 23259
rect 5199 23256 5213 23259
rect 5223 23259 6731 23263
rect 6745 23263 6779 23264
rect 6793 23263 6827 23264
rect 6745 23259 6827 23263
rect 7297 23263 7331 23264
rect 7345 23263 7379 23264
rect 7297 23259 7379 23263
rect 7393 23263 7427 23264
rect 7465 23263 7523 23264
rect 7596 23263 7598 23283
rect 7692 23264 7694 23283
rect 7657 23263 7715 23264
rect 7908 23263 7910 23283
rect 8124 23263 8126 23283
rect 8220 23263 8222 23283
rect 8316 23263 8318 23283
rect 8412 23263 8414 23283
rect 8700 23263 8702 23283
rect 8748 23264 8750 23283
rect 8785 23278 8788 23283
rect 8796 23278 8798 23283
rect 8833 23278 8836 23283
rect 8844 23278 8846 23283
rect 8795 23264 8798 23278
rect 8843 23264 8846 23278
rect 8857 23270 8861 23278
rect 8847 23264 8857 23270
rect 8737 23263 8771 23264
rect 7393 23259 8771 23263
rect 5223 23256 5237 23259
rect 5244 23256 5247 23259
rect 5292 23256 5294 23259
rect 5196 23254 5199 23256
rect 4931 23240 4934 23254
rect 5027 23240 5031 23254
rect 5113 23246 5117 23254
rect 5103 23240 5113 23246
rect 5195 23240 5199 23254
rect 5292 23240 5295 23256
rect 5460 23240 5462 23259
rect 5508 23240 5510 23259
rect 5556 23240 5558 23259
rect 5652 23240 5654 23259
rect 5748 23240 5750 23259
rect 5772 23240 5774 23259
rect 5844 23240 5846 23259
rect 4513 23239 4547 23240
rect 3961 23235 4547 23239
rect 4561 23239 4595 23240
rect 4849 23239 4883 23240
rect 5281 23239 5315 23240
rect 4561 23235 4883 23239
rect 5271 23235 5315 23239
rect 5353 23239 5387 23240
rect 5401 23239 5435 23240
rect 5353 23235 5435 23239
rect 5449 23239 5483 23240
rect 5497 23239 5531 23240
rect 5449 23235 5531 23239
rect 5545 23239 5579 23240
rect 5641 23239 5699 23240
rect 5737 23239 5795 23240
rect 5833 23239 5867 23240
rect 5545 23235 5867 23239
rect 5881 23239 5915 23240
rect 6108 23239 6110 23259
rect 6204 23239 6206 23259
rect 6276 23239 6278 23259
rect 6300 23239 6302 23259
rect 6372 23239 6374 23259
rect 6396 23239 6398 23259
rect 6492 23239 6494 23259
rect 6516 23240 6518 23259
rect 6588 23240 6590 23259
rect 6601 23254 6604 23259
rect 6612 23254 6614 23259
rect 6625 23254 6628 23259
rect 6636 23254 6638 23259
rect 6697 23254 6700 23259
rect 6708 23256 6710 23259
rect 6708 23254 6711 23256
rect 6793 23254 6796 23259
rect 6804 23256 6806 23259
rect 6804 23254 6807 23256
rect 7393 23254 7396 23259
rect 7404 23256 7406 23259
rect 7404 23254 7407 23256
rect 6611 23240 6614 23254
rect 6635 23240 6638 23254
rect 6707 23246 6711 23254
rect 6721 23246 6725 23254
rect 6707 23240 6721 23246
rect 6803 23240 6807 23254
rect 7403 23240 7407 23254
rect 7489 23254 7492 23259
rect 7500 23256 7502 23259
rect 7596 23256 7598 23259
rect 7500 23254 7503 23256
rect 7489 23246 7493 23254
rect 7479 23240 7489 23246
rect 7499 23240 7503 23254
rect 7596 23240 7599 23256
rect 7681 23254 7684 23259
rect 7692 23254 7694 23259
rect 7691 23240 7694 23254
rect 7908 23240 7910 23259
rect 6505 23239 6563 23240
rect 6577 23239 6611 23240
rect 5881 23235 6611 23239
rect 7585 23239 7619 23240
rect 7633 23239 7667 23240
rect 7585 23235 7667 23239
rect 7801 23239 7835 23240
rect 7873 23239 7931 23240
rect 8124 23239 8126 23259
rect 8220 23239 8222 23259
rect 8316 23239 8318 23259
rect 8412 23239 8414 23259
rect 8700 23239 8702 23259
rect 8737 23254 8740 23259
rect 8748 23254 8750 23259
rect 8747 23240 8750 23254
rect 8713 23239 8747 23240
rect 7801 23235 8747 23239
rect 4068 23232 4070 23235
rect 4068 23216 4071 23232
rect 4057 23215 4091 23216
rect 4164 23215 4166 23235
rect 4308 23216 4310 23235
rect 4575 23232 4589 23235
rect 5271 23232 5285 23235
rect 5292 23232 5295 23235
rect 5449 23230 5452 23235
rect 5460 23232 5462 23235
rect 5460 23230 5463 23232
rect 5497 23230 5500 23235
rect 5508 23232 5510 23235
rect 5508 23230 5511 23232
rect 5545 23230 5548 23235
rect 5556 23232 5558 23235
rect 5556 23230 5559 23232
rect 5641 23230 5644 23235
rect 5652 23232 5654 23235
rect 5652 23230 5655 23232
rect 5737 23230 5740 23235
rect 5748 23232 5750 23235
rect 5748 23230 5751 23232
rect 5377 23222 5381 23230
rect 5367 23216 5377 23222
rect 5459 23216 5463 23230
rect 5507 23216 5511 23230
rect 5555 23216 5559 23230
rect 5651 23216 5655 23230
rect 5747 23222 5751 23230
rect 5761 23230 5764 23235
rect 5772 23232 5774 23235
rect 5772 23230 5775 23232
rect 5833 23230 5836 23235
rect 5844 23232 5846 23235
rect 5844 23230 5847 23232
rect 5761 23222 5765 23230
rect 5747 23216 5761 23222
rect 5771 23216 5775 23230
rect 5843 23222 5847 23230
rect 5857 23222 5861 23230
rect 5843 23216 5857 23222
rect 4297 23215 4331 23216
rect 4057 23211 4331 23215
rect 4681 23215 4715 23216
rect 4825 23215 4859 23216
rect 4681 23211 4859 23215
rect 6001 23215 6035 23216
rect 6108 23215 6110 23235
rect 6204 23215 6206 23235
rect 6276 23215 6278 23235
rect 6300 23215 6302 23235
rect 6372 23215 6374 23235
rect 6396 23216 6398 23235
rect 6492 23216 6494 23235
rect 6505 23230 6508 23235
rect 6516 23230 6518 23235
rect 6577 23230 6580 23235
rect 6588 23230 6590 23235
rect 7585 23232 7589 23235
rect 7596 23232 7599 23235
rect 7897 23230 7900 23235
rect 7908 23232 7910 23235
rect 7908 23230 7911 23232
rect 6515 23216 6518 23230
rect 6587 23216 6590 23230
rect 6601 23222 6605 23230
rect 7897 23222 7901 23230
rect 6591 23216 6601 23222
rect 7887 23216 7897 23222
rect 7907 23216 7911 23230
rect 8124 23216 8126 23235
rect 8220 23216 8222 23235
rect 6385 23215 6443 23216
rect 6481 23215 6515 23216
rect 6001 23211 6515 23215
rect 8017 23215 8051 23216
rect 8089 23215 8147 23216
rect 8161 23215 8195 23216
rect 8017 23211 8195 23215
rect 8209 23215 8243 23216
rect 8316 23215 8318 23235
rect 8412 23216 8414 23235
rect 8700 23216 8702 23235
rect 8377 23215 8435 23216
rect 8593 23215 8627 23216
rect 8209 23211 8627 23215
rect 8641 23215 8675 23216
rect 8689 23215 8723 23216
rect 8641 23211 8723 23215
rect 4057 23208 4061 23211
rect 4068 23208 4071 23211
rect 4164 23208 4166 23211
rect 4164 23192 4167 23208
rect 4297 23206 4300 23211
rect 4308 23206 4310 23211
rect 4307 23192 4310 23206
rect 6108 23208 6110 23211
rect 6108 23192 6111 23208
rect 6204 23192 6206 23211
rect 6276 23192 6278 23211
rect 6300 23192 6302 23211
rect 6372 23192 6374 23211
rect 6385 23206 6388 23211
rect 6396 23206 6398 23211
rect 6481 23206 6484 23211
rect 6492 23208 6494 23211
rect 6492 23206 6495 23208
rect 8113 23206 8116 23211
rect 8124 23208 8126 23211
rect 8124 23206 8127 23208
rect 8209 23206 8212 23211
rect 8220 23208 8222 23211
rect 8316 23208 8318 23211
rect 8220 23206 8223 23208
rect 6395 23192 6398 23206
rect 6491 23198 6495 23206
rect 6505 23198 6509 23206
rect 8113 23198 8117 23206
rect 6491 23192 6505 23198
rect 8103 23192 8113 23198
rect 8123 23192 8127 23206
rect 8185 23198 8189 23206
rect 8175 23192 8185 23198
rect 8219 23192 8223 23206
rect 8316 23192 8319 23208
rect 8401 23206 8404 23211
rect 8412 23206 8414 23211
rect 8689 23206 8692 23211
rect 8700 23208 8702 23211
rect 8700 23206 8703 23208
rect 8411 23192 8414 23206
rect 8699 23192 8703 23206
rect 4153 23191 4187 23192
rect 4201 23191 4235 23192
rect 4153 23187 4235 23191
rect 6097 23191 6131 23192
rect 6169 23191 6227 23192
rect 6265 23191 6323 23192
rect 6361 23191 6395 23192
rect 6097 23187 6395 23191
rect 8305 23191 8339 23192
rect 8353 23191 8387 23192
rect 8305 23187 8387 23191
rect 8521 23191 8555 23192
rect 8569 23191 8603 23192
rect 8521 23187 8603 23191
rect 4153 23184 4157 23187
rect 4164 23184 4167 23187
rect 6097 23184 6101 23187
rect 6108 23184 6111 23187
rect 6193 23182 6196 23187
rect 6204 23184 6206 23187
rect 6204 23182 6207 23184
rect 6265 23182 6268 23187
rect 6276 23184 6278 23187
rect 6276 23182 6279 23184
rect 6193 23174 6197 23182
rect 6183 23168 6193 23174
rect 6203 23168 6207 23182
rect 6275 23174 6279 23182
rect 6289 23182 6292 23187
rect 6300 23184 6302 23187
rect 6300 23182 6303 23184
rect 6361 23182 6364 23187
rect 6372 23184 6374 23187
rect 8305 23184 8309 23187
rect 8316 23184 8319 23187
rect 6372 23182 6375 23184
rect 6289 23174 6293 23182
rect 6275 23168 6289 23174
rect 6299 23168 6303 23182
rect 6371 23174 6375 23182
rect 6385 23174 6389 23182
rect 6371 23168 6385 23174
use Control/control_ROUTED control_ROUTED_0
timestamp 1394713725
transform -1 0 32208 0 -1 26565
box 23 -3488 51336 3397
use Control/control_ROUTED control_ROUTED_1
timestamp 1394713725
transform -1 0 32284 0 -1 26557
box 23 -3488 51336 3397
use Datapath/datapath datapath_0
timestamp 1394713977
transform 1 0 7142 0 1 0
box 0 0 25013 22218
<< end >>
