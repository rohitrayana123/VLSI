magic
tech c035u
timestamp 1395747878
<< metal1 >>
rect 12520 8180 12538 8194
rect 9784 8156 9802 8170
rect 11488 8156 11506 8170
rect 12040 8158 17102 8168
rect 8056 8134 16250 8144
rect 20224 8132 20242 8146
rect 5584 8108 5602 8122
rect 5728 8110 18806 8120
rect 18820 8110 22490 8120
rect 84 8086 1730 8096
rect 2440 8086 9818 8096
rect 10720 8084 10738 8098
rect 11056 8086 15398 8096
rect 18796 8086 24122 8096
rect 84 8062 1778 8072
rect 2608 8062 22214 8072
rect 23908 8062 24722 8072
rect 3304 8038 13706 8048
rect 14416 8036 14434 8050
rect 15388 8038 15410 8048
rect 16192 8038 21362 8048
rect 23800 8038 27314 8048
rect 4168 8014 4778 8024
rect 5008 8012 5026 8026
rect 5128 8014 12830 8024
rect 13072 8014 23918 8024
rect 24280 8014 25622 8024
rect 27208 8012 27226 8026
rect 27256 8014 27266 8024
rect 5392 7990 13010 8000
rect 13024 7990 18218 8000
rect 18232 7990 27651 8000
rect 5608 7966 6782 7976
rect 7672 7966 20510 7976
rect 27280 7966 27651 7976
rect 6760 7942 17018 7952
rect 19432 7942 27290 7952
rect 27328 7942 27651 7952
rect 8488 7918 8666 7928
rect 9352 7918 12962 7928
rect 19864 7918 24770 7928
rect 27280 7918 27651 7928
rect 8584 7894 27266 7904
rect 27304 7894 27651 7904
rect 13480 7061 14090 7071
rect 13336 7037 16970 7047
rect 26560 7037 26930 7047
rect 11800 7013 11810 7023
rect 11992 7013 26546 7023
rect 11680 6989 11714 6999
rect 11776 6989 25946 6999
rect 11584 6965 17066 6975
rect 11512 6941 22778 6951
rect 11488 6917 17906 6927
rect 20440 6917 20474 6927
rect 11008 6893 11030 6903
rect 11128 6893 11162 6903
rect 11368 6893 12818 6903
rect 13312 6893 13802 6903
rect 14752 6893 20426 6903
rect 10552 6869 21770 6879
rect 9664 6845 9914 6855
rect 9976 6845 23810 6855
rect 9592 6821 21698 6831
rect 21712 6821 21794 6831
rect 9352 6797 23522 6807
rect 23536 6797 23954 6807
rect 9328 6773 9794 6783
rect 9952 6773 19874 6783
rect 9256 6749 9698 6759
rect 9880 6749 16442 6759
rect 16456 6749 26090 6759
rect 8920 6725 9290 6735
rect 9304 6725 10778 6735
rect 10792 6725 11090 6735
rect 11104 6725 12314 6735
rect 12328 6725 14738 6735
rect 14752 6725 17594 6735
rect 17608 6725 21074 6735
rect 21088 6725 24194 6735
rect 8728 6701 13970 6711
rect 13984 6701 25706 6711
rect 8416 6677 15626 6687
rect 18712 6677 18722 6687
rect 8392 6653 18698 6663
rect 8368 6629 21002 6639
rect 8344 6605 17762 6615
rect 17776 6605 20330 6615
rect 21544 6605 21566 6615
rect 8320 6581 8402 6591
rect 8560 6581 11210 6591
rect 11224 6581 14210 6591
rect 14224 6581 14282 6591
rect 14296 6581 18962 6591
rect 18976 6581 23762 6591
rect 8272 6557 17210 6567
rect 20536 6557 22178 6567
rect 22192 6557 24314 6567
rect 25096 6557 25346 6567
rect 8032 6533 21530 6543
rect 21544 6533 25850 6543
rect 7792 6509 7898 6519
rect 8008 6509 26906 6519
rect 7744 6485 25082 6495
rect 7720 6461 16538 6471
rect 17632 6461 22130 6471
rect 7720 6437 16850 6447
rect 17536 6437 19730 6447
rect 19744 6437 23114 6447
rect 7672 6413 12866 6423
rect 13144 6413 13634 6423
rect 13648 6413 14162 6423
rect 14176 6413 20522 6423
rect 20536 6413 23618 6423
rect 7624 6389 14366 6399
rect 14488 6389 19346 6399
rect 7600 6365 9506 6375
rect 9520 6365 12722 6375
rect 12928 6365 20090 6375
rect 20104 6365 25202 6375
rect 7240 6341 8618 6351
rect 8632 6341 19106 6351
rect 19120 6341 22442 6351
rect 22456 6341 22826 6351
rect 7240 6317 10658 6327
rect 10864 6317 11570 6327
rect 11584 6317 17522 6327
rect 17536 6317 17618 6327
rect 17632 6317 18722 6327
rect 7192 6293 20498 6303
rect 20512 6293 22202 6303
rect 7168 6269 15218 6279
rect 7072 6245 7250 6255
rect 7264 6245 13370 6255
rect 13384 6245 19082 6255
rect 19096 6245 22850 6255
rect 6952 6221 16946 6231
rect 6928 6197 22682 6207
rect 6880 6173 12674 6183
rect 12904 6173 18818 6183
rect 18832 6173 19010 6183
rect 19024 6173 20882 6183
rect 20896 6173 24338 6183
rect 24352 6173 27074 6183
rect 6856 6149 9842 6159
rect 9856 6149 10346 6159
rect 10360 6149 14834 6159
rect 14848 6149 18506 6159
rect 18520 6149 23930 6159
rect 23944 6149 26066 6159
rect 26080 6149 26666 6159
rect 6472 6125 22250 6135
rect 6328 6101 21242 6111
rect 23056 6101 23138 6111
rect 23224 6101 23282 6111
rect 6232 6077 9266 6087
rect 9280 6077 10946 6087
rect 10960 6077 16862 6087
rect 21352 6077 22418 6087
rect 22432 6077 25754 6087
rect 6184 6053 25298 6063
rect 6136 6029 6362 6039
rect 6376 6029 6794 6039
rect 6808 6029 7442 6039
rect 7456 6029 10298 6039
rect 10312 6029 14714 6039
rect 14728 6029 19178 6039
rect 19192 6029 21266 6039
rect 21280 6029 23042 6039
rect 23056 6029 23066 6039
rect 23080 6029 23210 6039
rect 23224 6029 25778 6039
rect 25792 6029 26330 6039
rect 6040 6005 11762 6015
rect 11776 6005 21602 6015
rect 22984 6005 24410 6015
rect 5992 5981 7370 5991
rect 7504 5981 8474 5991
rect 8488 5981 10034 5991
rect 10048 5981 11330 5991
rect 11344 5981 13346 5991
rect 13360 5981 14258 5991
rect 14272 5981 20402 5991
rect 20416 5981 22970 5991
rect 22984 5981 23450 5991
rect 5944 5957 7922 5967
rect 7936 5957 10394 5967
rect 10408 5957 10922 5967
rect 10936 5957 12770 5967
rect 12784 5957 13586 5967
rect 13600 5957 21338 5967
rect 21352 5957 24842 5967
rect 24856 5957 25994 5967
rect 5728 5933 10010 5943
rect 10336 5933 23186 5943
rect 5656 5909 20786 5919
rect 20800 5909 22658 5919
rect 5368 5885 5378 5895
rect 5392 5885 9962 5895
rect 9976 5885 19826 5895
rect 19840 5885 25130 5895
rect 5320 5861 16994 5871
rect 5272 5837 7010 5847
rect 7024 5837 24890 5847
rect 5224 5813 14474 5823
rect 14536 5813 21566 5823
rect 25192 5813 25442 5823
rect 5200 5789 10874 5799
rect 10888 5789 13874 5799
rect 13936 5789 14306 5799
rect 14464 5789 25178 5799
rect 5104 5765 17474 5775
rect 5056 5741 23162 5751
rect 5032 5717 6602 5727
rect 6760 5717 8906 5727
rect 9016 5717 20186 5727
rect 23584 5717 23594 5727
rect 5008 5693 13850 5703
rect 13864 5693 13922 5703
rect 13936 5693 16682 5703
rect 16696 5693 20234 5703
rect 20248 5693 20690 5703
rect 20704 5693 20882 5703
rect 20896 5693 21674 5703
rect 21688 5693 23570 5703
rect 4936 5669 15746 5679
rect 15760 5669 16346 5679
rect 16360 5669 18830 5679
rect 18844 5669 19898 5679
rect 19912 5669 20762 5679
rect 20776 5669 23858 5679
rect 4864 5645 8186 5655
rect 8200 5645 8930 5655
rect 8944 5645 11258 5655
rect 11272 5645 15530 5655
rect 15544 5645 18578 5655
rect 18592 5645 18794 5655
rect 18808 5645 24842 5655
rect 4816 5621 6482 5631
rect 6544 5621 13778 5631
rect 13960 5621 17306 5631
rect 4768 5597 24794 5607
rect 4720 5573 9050 5583
rect 9232 5573 9626 5583
rect 9784 5573 22490 5583
rect 4672 5549 10370 5559
rect 10384 5549 16298 5559
rect 4672 5525 7802 5535
rect 7888 5525 12098 5535
rect 12112 5525 14450 5535
rect 14464 5525 16922 5535
rect 16936 5525 25562 5535
rect 4624 5501 26210 5511
rect 4504 5477 11786 5487
rect 11800 5477 21578 5487
rect 4504 5453 16370 5463
rect 16768 5453 26738 5463
rect 4456 5429 8030 5439
rect 8044 5429 10538 5439
rect 10552 5429 13682 5439
rect 13696 5429 17402 5439
rect 17416 5429 23426 5439
rect 4384 5405 18242 5415
rect 18256 5405 19274 5415
rect 19288 5405 25226 5415
rect 4384 5381 8450 5391
rect 8512 5381 23282 5391
rect 4360 5357 9650 5367
rect 9664 5357 16490 5367
rect 16504 5357 17186 5367
rect 4312 5333 14570 5343
rect 14872 5333 16130 5343
rect 16528 5333 16766 5343
rect 4288 5309 17570 5319
rect 4264 5285 7298 5295
rect 7360 5285 12602 5295
rect 12664 5285 13946 5295
rect 14248 5285 14426 5295
rect 14512 5285 14546 5295
rect 14632 5285 24074 5295
rect 4240 5261 8978 5271
rect 9040 5261 22802 5271
rect 4216 5237 9050 5247
rect 9112 5237 17282 5247
rect 17464 5237 17714 5247
rect 19048 5237 19922 5247
rect 19936 5237 22058 5247
rect 4168 5213 17642 5223
rect 18952 5213 20498 5223
rect 20512 5213 21650 5223
rect 4144 5189 5090 5199
rect 5104 5189 11450 5199
rect 11464 5189 14234 5199
rect 14416 5189 20642 5199
rect 4048 5165 5354 5175
rect 5368 5165 10226 5175
rect 10240 5165 11666 5175
rect 11680 5165 17738 5175
rect 18544 5165 20282 5175
rect 21160 5165 21494 5175
rect 4024 5141 6650 5151
rect 6712 5141 9098 5151
rect 9112 5141 12698 5151
rect 12784 5141 26690 5151
rect 3952 5117 10490 5127
rect 10624 5117 10670 5127
rect 10720 5117 21818 5127
rect 3928 5093 5522 5103
rect 5584 5093 8006 5103
rect 8020 5093 11474 5103
rect 11488 5093 14498 5103
rect 14512 5093 18002 5103
rect 18016 5093 18146 5103
rect 18160 5093 19922 5103
rect 19936 5093 24122 5103
rect 24136 5093 24194 5103
rect 3880 5069 13466 5079
rect 13744 5069 21938 5079
rect 21952 5069 24722 5079
rect 24736 5069 25394 5079
rect 3856 5045 15242 5055
rect 16288 5045 25274 5055
rect 25840 5045 25862 5055
rect 3712 5021 5426 5031
rect 5440 5021 15962 5031
rect 15976 5021 26234 5031
rect 3664 4997 4586 5007
rect 4600 4997 9026 5007
rect 9040 4997 10082 5007
rect 10096 4997 10898 5007
rect 10912 4997 11138 5007
rect 11152 4997 16322 5007
rect 16336 4997 16514 5007
rect 16528 4997 24938 5007
rect 24952 4997 25238 5007
rect 25252 4997 25826 5007
rect 25840 4997 26594 5007
rect 3592 4973 17450 4983
rect 17464 4973 23714 4983
rect 3568 4949 21146 4959
rect 3496 4925 13106 4935
rect 13120 4925 14282 4935
rect 14344 4925 24050 4935
rect 3472 4901 6458 4911
rect 6472 4901 7850 4911
rect 7864 4901 8786 4911
rect 8800 4901 9218 4911
rect 9232 4901 9866 4911
rect 9880 4901 11522 4911
rect 11536 4901 23642 4911
rect 23656 4901 23978 4911
rect 23992 4901 24626 4911
rect 24640 4901 24890 4911
rect 3424 4877 17498 4887
rect 17512 4877 21050 4887
rect 3400 4853 9338 4863
rect 9352 4853 13994 4863
rect 14008 4853 21122 4863
rect 21136 4853 23690 4863
rect 3304 4829 3770 4839
rect 3784 4829 7634 4839
rect 7648 4829 8954 4839
rect 8968 4829 9386 4839
rect 9400 4829 11378 4839
rect 11392 4829 20330 4839
rect 20968 4829 21098 4839
rect 3280 4805 19658 4815
rect 20824 4805 21626 4815
rect 3256 4781 13370 4791
rect 13384 4781 13514 4791
rect 13672 4781 13994 4791
rect 14128 4781 19706 4791
rect 20272 4781 20450 4791
rect 20632 4781 21410 4791
rect 3232 4757 7970 4767
rect 7984 4757 16274 4767
rect 16288 4757 18410 4767
rect 18424 4757 20354 4767
rect 20560 4757 21494 4767
rect 3184 4733 9986 4743
rect 10288 4733 15098 4743
rect 15112 4733 19514 4743
rect 19624 4733 22706 4743
rect 22720 4733 25346 4743
rect 3136 4709 8162 4719
rect 8176 4709 11930 4719
rect 11944 4709 12194 4719
rect 12208 4709 22946 4719
rect 3040 4685 24434 4695
rect 3016 4661 17042 4671
rect 17104 4661 26786 4671
rect 2992 4637 6074 4647
rect 6136 4637 7130 4647
rect 7144 4637 19850 4647
rect 20176 4637 24314 4647
rect 2920 4613 6146 4623
rect 6160 4613 9146 4623
rect 9160 4613 13610 4623
rect 13624 4613 15482 4623
rect 15496 4613 18890 4623
rect 18904 4613 24506 4623
rect 2896 4589 5282 4599
rect 5344 4589 17330 4599
rect 18496 4589 18626 4599
rect 18880 4589 19154 4599
rect 19216 4589 22262 4599
rect 2872 4565 12914 4575
rect 12928 4565 21554 4575
rect 2824 4541 6506 4551
rect 6712 4541 19778 4551
rect 19984 4541 23450 4551
rect 2752 4517 21194 4527
rect 22096 4517 22142 4527
rect 2680 4493 4586 4503
rect 4600 4493 4682 4503
rect 4696 4493 6626 4503
rect 6640 4493 13226 4503
rect 13240 4493 16250 4503
rect 16264 4493 21002 4503
rect 21016 4493 21314 4503
rect 21328 4493 22874 4503
rect 22888 4493 23786 4503
rect 2656 4469 6578 4479
rect 6592 4469 7778 4479
rect 7792 4469 9578 4479
rect 9592 4469 23306 4479
rect 2608 4445 11690 4455
rect 11752 4445 17138 4455
rect 17824 4445 26570 4455
rect 2584 4421 4514 4431
rect 4528 4421 23186 4431
rect 24376 4421 24578 4431
rect 26152 4421 26378 4431
rect 2560 4397 5762 4407
rect 5848 4397 16766 4407
rect 16780 4397 21194 4407
rect 21208 4397 22226 4407
rect 22240 4397 22298 4407
rect 23344 4397 23498 4407
rect 24232 4397 25610 4407
rect 26056 4397 26162 4407
rect 26320 4397 26474 4407
rect 26536 4397 26882 4407
rect 2536 4373 15338 4383
rect 15352 4373 21746 4383
rect 21760 4373 24026 4383
rect 24112 4373 24446 4383
rect 24688 4373 26762 4383
rect 2512 4349 9554 4359
rect 9568 4349 11426 4359
rect 11440 4349 15314 4359
rect 15328 4349 25058 4359
rect 25120 4349 27266 4359
rect 2440 4325 14642 4335
rect 14656 4325 22082 4335
rect 22096 4325 22418 4335
rect 22576 4325 22610 4335
rect 22768 4325 22922 4335
rect 23128 4325 26930 4335
rect 2344 4301 8666 4311
rect 8680 4301 8786 4311
rect 8800 4301 19826 4311
rect 19840 4301 23810 4311
rect 23824 4301 24866 4311
rect 25072 4301 25238 4311
rect 26008 4301 26066 4311
rect 2248 4277 9530 4287
rect 9616 4277 27314 4287
rect 2248 4253 20378 4263
rect 21496 4253 25634 4263
rect 2200 4229 7418 4239
rect 7504 4229 26186 4239
rect 26200 4229 26330 4239
rect 2128 4205 20714 4215
rect 20728 4205 22634 4215
rect 23320 4205 23426 4215
rect 23488 4205 26354 4215
rect 2080 4181 8210 4191
rect 8224 4181 20258 4191
rect 20320 4181 22898 4191
rect 23872 4181 23930 4191
rect 2008 4157 11858 4167
rect 11872 4157 12794 4167
rect 12808 4157 13394 4167
rect 13576 4157 17690 4167
rect 17992 4157 19130 4167
rect 19864 4157 20186 4167
rect 21880 4157 23354 4167
rect 1960 4133 2690 4143
rect 2704 4133 3986 4143
rect 4048 4133 4058 4143
rect 4120 4133 8642 4143
rect 8656 4133 12146 4143
rect 12232 4133 12602 4143
rect 12664 4133 14090 4143
rect 14104 4133 26042 4143
rect 1912 4109 3746 4119
rect 3760 4109 9410 4119
rect 9472 4109 26714 4119
rect 1864 4085 7394 4095
rect 7408 4085 26234 4095
rect 1840 4061 13418 4071
rect 13624 4061 14210 4071
rect 14992 4061 27026 4071
rect 1672 4037 2498 4047
rect 2512 4037 7274 4047
rect 7288 4037 10202 4047
rect 10312 4037 10346 4047
rect 10432 4037 10466 4047
rect 10648 4037 12290 4047
rect 12304 4037 22442 4047
rect 22456 4037 22538 4047
rect 22552 4037 23138 4047
rect 23152 4037 27122 4047
rect 1624 4013 6482 4023
rect 6496 4013 8234 4023
rect 8248 4013 11354 4023
rect 11368 4013 22106 4023
rect 22120 4013 26426 4023
rect 84 3989 10610 3999
rect 10624 3989 24554 3999
rect 26440 3989 27194 3999
rect 84 3965 6746 3975
rect 6832 3965 9194 3975
rect 9208 3965 10058 3975
rect 10072 3965 12578 3975
rect 12592 3965 13202 3975
rect 13216 3965 23354 3975
rect 1744 3941 2786 3951
rect 2848 3941 4274 3951
rect 4288 3941 20594 3951
rect 20608 3941 22142 3951
rect 22240 3941 22262 3951
rect 22312 3941 23258 3951
rect 1792 3917 9482 3927
rect 9544 3917 9842 3927
rect 10000 3917 15266 3927
rect 15280 3917 24266 3927
rect 2056 3893 4802 3903
rect 4816 3893 6338 3903
rect 6352 3893 24962 3903
rect 2104 3869 2306 3879
rect 2320 3869 3674 3879
rect 3688 3869 7058 3879
rect 7072 3869 7370 3879
rect 7384 3869 15434 3879
rect 15448 3869 16610 3879
rect 16624 3869 16706 3879
rect 16720 3869 18434 3879
rect 18448 3869 23066 3879
rect 23080 3869 23330 3879
rect 23344 3869 26306 3879
rect 2296 3845 8210 3855
rect 8224 3845 10754 3855
rect 10768 3845 11618 3855
rect 11632 3845 13154 3855
rect 13168 3845 26618 3855
rect 2320 3821 8690 3831
rect 8704 3821 9314 3831
rect 9328 3821 11234 3831
rect 11248 3821 13274 3831
rect 13288 3821 14330 3831
rect 14344 3821 15458 3831
rect 15472 3821 15986 3831
rect 16000 3821 16562 3831
rect 16576 3821 18770 3831
rect 18784 3821 20018 3831
rect 20032 3821 22754 3831
rect 22768 3821 23546 3831
rect 23560 3821 23666 3831
rect 23680 3821 26402 3831
rect 2368 3797 15986 3807
rect 16120 3797 22994 3807
rect 2368 3773 4466 3783
rect 4480 3773 5474 3783
rect 5488 3773 7394 3783
rect 7408 3773 13658 3783
rect 13672 3773 23090 3783
rect 23104 3773 25802 3783
rect 2416 3749 8066 3759
rect 8128 3749 8258 3759
rect 8272 3749 13898 3759
rect 13912 3749 14882 3759
rect 15208 3749 20666 3759
rect 20680 3749 22946 3759
rect 2416 3725 5498 3735
rect 5512 3725 5954 3735
rect 5968 3725 12866 3735
rect 12880 3725 17786 3735
rect 17800 3725 20042 3735
rect 20056 3725 22562 3735
rect 2440 3701 2858 3711
rect 2872 3701 6050 3711
rect 6064 3701 9242 3711
rect 9256 3701 10994 3711
rect 11008 3701 11402 3711
rect 11416 3701 15770 3711
rect 15784 3701 19226 3711
rect 19240 3701 20930 3711
rect 20944 3701 25922 3711
rect 2464 3677 12746 3687
rect 12832 3677 12962 3687
rect 13168 3677 26858 3687
rect 2464 3653 26498 3663
rect 2536 3629 5594 3639
rect 5608 3629 6818 3639
rect 6832 3629 10418 3639
rect 10432 3629 16586 3639
rect 16600 3629 16730 3639
rect 16744 3629 18314 3639
rect 18328 3629 25490 3639
rect 2632 3605 5066 3615
rect 5080 3605 26138 3615
rect 2656 3581 7946 3591
rect 7960 3581 11030 3591
rect 11044 3581 11114 3591
rect 11128 3581 20618 3591
rect 22000 3581 26450 3591
rect 2680 3557 15410 3567
rect 15472 3557 15530 3567
rect 15640 3557 16394 3567
rect 16600 3557 16970 3567
rect 17488 3557 17762 3567
rect 18064 3557 26834 3567
rect 2728 3533 24362 3543
rect 24376 3533 26474 3543
rect 2752 3509 5450 3519
rect 5464 3509 6386 3519
rect 6400 3509 6410 3519
rect 6424 3509 16226 3519
rect 16240 3509 26210 3519
rect 2776 3485 16442 3495
rect 16672 3485 26978 3495
rect 3016 3461 25658 3471
rect 3064 3437 18914 3447
rect 19024 3437 19346 3447
rect 20008 3437 26162 3447
rect 3088 3413 9746 3423
rect 10072 3413 21290 3423
rect 3160 3389 3554 3399
rect 3616 3389 24170 3399
rect 3328 3365 26762 3375
rect 3376 3341 20834 3351
rect 3376 3317 8450 3327
rect 8464 3317 9794 3327
rect 9808 3317 14066 3327
rect 14080 3317 14594 3327
rect 14608 3317 17546 3327
rect 17560 3317 18482 3327
rect 18496 3317 18602 3327
rect 18616 3317 19946 3327
rect 19960 3317 20138 3327
rect 3424 3293 8138 3303
rect 8152 3293 8858 3303
rect 8872 3293 9890 3303
rect 9904 3293 18674 3303
rect 18688 3293 21458 3303
rect 21472 3293 22610 3303
rect 3520 3269 22874 3279
rect 3616 3245 7610 3255
rect 7624 3245 15866 3255
rect 15880 3245 16634 3255
rect 16720 3245 16862 3255
rect 18760 3245 25418 3255
rect 3640 3221 6914 3231
rect 6928 3221 13706 3231
rect 13720 3221 16466 3231
rect 16480 3221 16802 3231
rect 16816 3221 26114 3231
rect 3760 3197 17234 3207
rect 18784 3197 18830 3207
rect 18904 3197 19274 3207
rect 20032 3197 20354 3207
rect 25432 3197 26258 3207
rect 3784 3173 20210 3183
rect 3808 3149 26810 3159
rect 3856 3125 6938 3135
rect 6952 3125 9818 3135
rect 9832 3125 13754 3135
rect 13768 3125 15890 3135
rect 15904 3125 16826 3135
rect 16840 3125 18554 3135
rect 18832 3125 26954 3135
rect 3880 3101 8882 3111
rect 8896 3101 9674 3111
rect 9688 3101 16034 3111
rect 16048 3101 17666 3111
rect 17680 3101 18458 3111
rect 18472 3101 20738 3111
rect 20752 3101 20978 3111
rect 20992 3101 22922 3111
rect 3904 3077 14522 3087
rect 15232 3077 17018 3087
rect 17032 3077 18098 3087
rect 18112 3077 19322 3087
rect 19336 3077 23402 3087
rect 23416 3077 24650 3087
rect 24664 3077 25442 3087
rect 25456 3077 25514 3087
rect 3928 3053 4778 3063
rect 4792 3053 7730 3063
rect 7744 3053 9626 3063
rect 9640 3053 12962 3063
rect 12976 3053 16202 3063
rect 16216 3053 17714 3063
rect 17728 3053 18578 3063
rect 18592 3053 19082 3063
rect 19096 3053 20714 3063
rect 3952 3029 5810 3039
rect 5896 3029 25370 3039
rect 4024 3005 11306 3015
rect 11320 3005 12386 3015
rect 12400 3005 18650 3015
rect 20224 3005 20402 3015
rect 20752 3005 21578 3015
rect 4120 2981 6554 2991
rect 6688 2981 11882 2991
rect 12256 2981 14546 2991
rect 15400 2981 16178 2991
rect 16240 2981 16298 2991
rect 16744 2981 17066 2991
rect 18472 2981 20906 2991
rect 4144 2957 6554 2967
rect 6568 2957 21386 2967
rect 21400 2957 26090 2967
rect 4216 2933 9722 2943
rect 9736 2933 12074 2943
rect 12088 2933 13082 2943
rect 13096 2933 13322 2943
rect 13336 2933 13826 2943
rect 13840 2933 18362 2943
rect 18376 2933 18866 2943
rect 18880 2933 21218 2943
rect 21232 2933 22538 2943
rect 22552 2933 24098 2943
rect 4240 2909 4874 2919
rect 4888 2909 6794 2919
rect 6808 2909 7466 2919
rect 7480 2909 7634 2919
rect 7648 2909 7826 2919
rect 7840 2909 8834 2919
rect 8848 2909 10178 2919
rect 10192 2909 17114 2919
rect 17128 2909 21026 2919
rect 4408 2885 10082 2895
rect 10336 2885 11546 2895
rect 11608 2885 27651 2895
rect 4432 2861 14138 2871
rect 14152 2861 22346 2871
rect 4456 2837 14114 2847
rect 14128 2837 16394 2847
rect 16408 2837 19058 2847
rect 19072 2837 24746 2847
rect 24760 2837 26378 2847
rect 4576 2813 17546 2823
rect 4696 2789 11810 2799
rect 12352 2789 21434 2799
rect 21448 2789 24446 2799
rect 4792 2765 6266 2775
rect 6280 2765 18626 2775
rect 4888 2741 6722 2751
rect 6736 2741 15506 2751
rect 15568 2741 20066 2751
rect 20080 2741 22178 2751
rect 4936 2717 10970 2727
rect 10984 2717 13490 2727
rect 14080 2717 14366 2727
rect 15496 2717 23234 2727
rect 4984 2693 25274 2703
rect 5008 2669 5474 2679
rect 5488 2669 9170 2679
rect 9184 2669 11714 2679
rect 11728 2669 14570 2679
rect 14584 2669 25862 2679
rect 5152 2645 13298 2655
rect 13312 2645 16898 2655
rect 16912 2645 21410 2655
rect 21424 2645 25730 2655
rect 5176 2621 21266 2631
rect 5224 2597 8738 2607
rect 8752 2597 14690 2607
rect 14704 2597 26282 2607
rect 5320 2573 9914 2583
rect 9928 2573 10826 2583
rect 10840 2573 14810 2583
rect 14824 2573 19154 2583
rect 5416 2549 26498 2559
rect 5584 2525 9698 2535
rect 9784 2525 19370 2535
rect 5608 2501 12506 2511
rect 12568 2501 25322 2511
rect 5704 2477 10106 2487
rect 10456 2477 24386 2487
rect 6088 2453 24290 2463
rect 6304 2429 6722 2439
rect 6736 2429 10154 2439
rect 10168 2429 11162 2439
rect 11176 2429 22586 2439
rect 6376 2405 10730 2415
rect 10744 2405 15578 2415
rect 15592 2405 20114 2415
rect 6520 2381 9458 2391
rect 9472 2381 19466 2391
rect 19480 2381 20810 2391
rect 6880 2357 14354 2367
rect 14368 2357 18218 2367
rect 18232 2357 18386 2367
rect 6976 2333 19802 2343
rect 7000 2309 13874 2319
rect 13888 2309 14186 2319
rect 14200 2309 21170 2319
rect 21184 2309 21362 2319
rect 21376 2309 25226 2319
rect 7168 2285 19250 2295
rect 7192 2261 14042 2271
rect 14704 2261 22730 2271
rect 22744 2261 24986 2271
rect 7264 2237 24002 2247
rect 7288 2213 20450 2223
rect 20464 2213 21626 2223
rect 7432 2189 7442 2199
rect 7528 2189 21890 2199
rect 7576 2165 23738 2175
rect 7768 2141 22346 2151
rect 7864 2117 8006 2127
rect 8104 2117 10466 2127
rect 10480 2117 26642 2127
rect 7960 2093 8030 2103
rect 8176 2093 8186 2103
rect 8296 2093 14426 2103
rect 14440 2093 16178 2103
rect 16192 2093 25970 2103
rect 7984 2069 25034 2079
rect 8032 2045 13538 2055
rect 13552 2045 18986 2055
rect 19264 2045 20474 2055
rect 25048 2045 25202 2055
rect 8320 2021 9434 2031
rect 9448 2021 22634 2031
rect 8368 1997 8810 2007
rect 8968 1997 8978 2007
rect 9088 1997 18266 2007
rect 19000 1997 19418 2007
rect 8392 1973 8930 1983
rect 8944 1973 10670 1983
rect 10684 1973 23594 1983
rect 8584 1949 12674 1959
rect 12688 1949 13010 1959
rect 13024 1949 13802 1959
rect 13816 1949 16418 1959
rect 16432 1949 21242 1959
rect 21256 1949 23378 1959
rect 23392 1949 24482 1959
rect 24496 1949 26642 1959
rect 8608 1925 26522 1935
rect 8776 1901 9362 1911
rect 9568 1901 10130 1911
rect 10144 1901 11834 1911
rect 11848 1901 17426 1911
rect 17440 1901 24530 1911
rect 9160 1877 11642 1887
rect 11848 1877 12026 1887
rect 12424 1877 12890 1887
rect 12904 1877 13250 1887
rect 13264 1877 18362 1887
rect 18376 1877 23882 1887
rect 23896 1877 24074 1887
rect 24088 1877 26018 1887
rect 26032 1877 26618 1887
rect 9688 1853 10034 1863
rect 10504 1853 21050 1863
rect 21064 1853 26882 1863
rect 9832 1829 19586 1839
rect 10840 1805 10946 1815
rect 11032 1805 20858 1815
rect 10936 1781 27290 1791
rect 11176 1757 11954 1767
rect 12472 1757 13754 1767
rect 15664 1757 20786 1767
rect 20800 1757 22850 1767
rect 22864 1757 23906 1767
rect 11200 1733 14018 1743
rect 16024 1733 25898 1743
rect 11248 1709 27242 1719
rect 11320 1685 13442 1695
rect 13456 1685 23498 1695
rect 23512 1685 24242 1695
rect 24256 1685 25154 1695
rect 11440 1661 11474 1671
rect 12472 1661 14306 1671
rect 16336 1661 16490 1671
rect 23920 1661 24410 1671
rect 25168 1661 25394 1671
rect 13216 1637 13634 1647
rect 27328 1637 27651 1647
rect 13432 1613 13970 1623
rect 27304 1613 27651 1623
rect 13552 1589 19298 1599
rect 19312 1589 24146 1599
rect 27280 1589 27651 1599
rect 26835 1560 27267 1570
rect 26835 1537 27267 1547
rect 26835 1499 27267 1524
rect 26835 854 27267 879
rect 13264 756 15530 766
rect 11944 732 20354 742
rect 11536 708 19946 718
rect 10384 684 21914 694
rect 10288 660 19130 670
rect 19144 660 26114 670
rect 9712 636 13586 646
rect 13840 636 14930 646
rect 16912 636 19658 646
rect 9016 612 10202 622
rect 10216 612 11066 622
rect 11080 612 26186 622
rect 8680 588 9914 598
rect 10024 588 16058 598
rect 16792 588 17642 598
rect 18136 588 20042 598
rect 21400 588 23954 598
rect 8488 564 10658 574
rect 11176 562 11194 576
rect 11272 564 16082 574
rect 16504 564 22010 574
rect 22600 564 23978 574
rect 7996 540 12602 550
rect 12808 540 18506 550
rect 21112 540 22898 550
rect 7888 516 14210 526
rect 15040 516 15074 526
rect 15376 516 23138 526
rect 7576 492 9434 502
rect 9616 492 26378 502
rect 7528 468 15818 478
rect 15928 468 21962 478
rect 22144 468 26834 478
rect 6664 444 13706 454
rect 13792 444 14402 454
rect 14968 444 20138 454
rect 20560 444 22658 454
rect 23272 444 23666 454
rect 26824 444 26858 454
rect 6424 420 7130 430
rect 7336 420 24482 430
rect 26776 420 27651 430
rect 6280 396 10778 406
rect 10888 396 15146 406
rect 15304 396 23402 406
rect 23920 394 23938 408
rect 26728 396 26810 406
rect 5560 372 6602 382
rect 6616 372 17858 382
rect 5272 348 7034 358
rect 7096 348 20402 358
rect 5248 324 8498 334
rect 8560 324 14162 334
rect 4744 300 11546 310
rect 11728 300 23690 310
rect 4480 276 18602 286
rect 4360 252 4826 262
rect 5032 252 26666 262
rect 4336 228 9410 238
rect 9424 228 15698 238
rect 4168 204 20594 214
rect 4072 180 7298 190
rect 7456 180 11642 190
rect 11896 180 17690 190
rect 3736 156 18170 166
rect 3712 132 22994 142
rect 3664 108 15002 118
rect 1696 84 20450 94
rect 84 60 23498 70
rect 26872 60 27651 70
rect 84 36 2234 46
rect 2560 36 4538 46
rect 4552 36 22778 46
rect 26824 36 27651 46
rect 3568 12 14426 22
rect 26848 12 27651 22
<< m2contact >>
rect 12506 8180 12520 8194
rect 9770 8156 9784 8170
rect 11474 8156 11488 8170
rect 12026 8156 12040 8170
rect 17102 8156 17116 8170
rect 8042 8132 8056 8146
rect 16250 8132 16264 8146
rect 20210 8132 20224 8146
rect 5570 8108 5584 8122
rect 5714 8108 5728 8122
rect 18806 8108 18820 8122
rect 22490 8108 22504 8122
rect 70 8084 84 8098
rect 1730 8084 1744 8098
rect 2426 8084 2440 8098
rect 9818 8084 9832 8098
rect 10706 8084 10720 8098
rect 11042 8084 11056 8098
rect 15398 8084 15412 8098
rect 18782 8084 18796 8098
rect 24122 8084 24136 8098
rect 70 8060 84 8074
rect 1778 8060 1792 8074
rect 2594 8060 2608 8074
rect 22214 8060 22228 8074
rect 23894 8060 23908 8074
rect 24722 8060 24736 8074
rect 3290 8036 3304 8050
rect 13706 8036 13720 8050
rect 14402 8036 14416 8050
rect 15374 8036 15388 8050
rect 15410 8036 15424 8050
rect 16178 8036 16192 8050
rect 21362 8036 21376 8050
rect 23786 8036 23800 8050
rect 27314 8036 27328 8050
rect 4154 8012 4168 8026
rect 4778 8012 4792 8026
rect 4994 8012 5008 8026
rect 5114 8012 5128 8026
rect 12830 8012 12844 8026
rect 13058 8012 13072 8026
rect 23918 8012 23932 8026
rect 24266 8012 24280 8026
rect 25622 8012 25636 8026
rect 27194 8012 27208 8026
rect 27242 8012 27256 8026
rect 27266 8012 27280 8026
rect 5378 7988 5392 8002
rect 13010 7988 13024 8002
rect 18218 7988 18232 8002
rect 27651 7988 27665 8002
rect 5594 7964 5608 7978
rect 6782 7964 6796 7978
rect 7658 7964 7672 7978
rect 20510 7964 20524 7978
rect 27266 7964 27280 7978
rect 27651 7964 27665 7978
rect 6746 7940 6760 7954
rect 17018 7940 17032 7954
rect 19418 7940 19432 7954
rect 27290 7940 27304 7954
rect 27314 7940 27328 7954
rect 27651 7940 27665 7954
rect 8474 7916 8488 7930
rect 8666 7916 8680 7930
rect 9338 7916 9352 7930
rect 12962 7916 12976 7930
rect 19850 7916 19864 7930
rect 24770 7916 24784 7930
rect 27266 7916 27280 7930
rect 27651 7916 27665 7930
rect 8570 7892 8584 7906
rect 27266 7892 27280 7906
rect 27290 7892 27304 7906
rect 27651 7892 27665 7906
rect 13466 7059 13480 7073
rect 14090 7059 14104 7073
rect 13322 7035 13336 7049
rect 16970 7035 16984 7049
rect 26546 7035 26560 7049
rect 26930 7035 26944 7049
rect 11786 7011 11800 7025
rect 11810 7011 11824 7025
rect 11978 7011 11992 7025
rect 26546 7011 26560 7025
rect 11666 6987 11680 7001
rect 11714 6987 11728 7001
rect 11762 6987 11776 7001
rect 25946 6987 25960 7001
rect 11570 6963 11584 6977
rect 17066 6963 17080 6977
rect 11498 6939 11512 6953
rect 22778 6939 22792 6953
rect 11474 6915 11488 6929
rect 17906 6915 17920 6929
rect 20426 6915 20440 6929
rect 20474 6915 20488 6929
rect 10994 6891 11008 6905
rect 11030 6891 11044 6905
rect 11114 6891 11128 6905
rect 11162 6891 11176 6905
rect 11354 6891 11368 6905
rect 12818 6891 12832 6905
rect 13298 6891 13312 6905
rect 13802 6891 13816 6905
rect 14738 6891 14752 6905
rect 20426 6891 20440 6905
rect 10538 6867 10552 6881
rect 21770 6867 21784 6881
rect 9650 6843 9664 6857
rect 9914 6843 9928 6857
rect 9962 6843 9976 6857
rect 23810 6843 23824 6857
rect 9578 6819 9592 6833
rect 21698 6819 21712 6833
rect 21794 6819 21808 6833
rect 9338 6795 9352 6809
rect 23522 6795 23536 6809
rect 23954 6795 23968 6809
rect 9314 6771 9328 6785
rect 9794 6771 9808 6785
rect 9938 6771 9952 6785
rect 19874 6771 19888 6785
rect 9242 6747 9256 6761
rect 9698 6747 9712 6761
rect 9866 6747 9880 6761
rect 16442 6747 16456 6761
rect 26090 6747 26104 6761
rect 8906 6723 8920 6737
rect 9290 6723 9304 6737
rect 10778 6723 10792 6737
rect 11090 6723 11104 6737
rect 12314 6723 12328 6737
rect 14738 6723 14752 6737
rect 17594 6723 17608 6737
rect 21074 6723 21088 6737
rect 24194 6723 24208 6737
rect 8714 6699 8728 6713
rect 13970 6699 13984 6713
rect 25706 6699 25720 6713
rect 8402 6675 8416 6689
rect 15626 6675 15640 6689
rect 18698 6675 18712 6689
rect 18722 6675 18736 6689
rect 8378 6651 8392 6665
rect 18698 6651 18712 6665
rect 8354 6627 8368 6641
rect 21002 6627 21016 6641
rect 8330 6603 8344 6617
rect 17762 6603 17776 6617
rect 20330 6603 20344 6617
rect 21530 6603 21544 6617
rect 21566 6603 21580 6617
rect 8306 6579 8320 6593
rect 8402 6579 8416 6593
rect 8546 6579 8560 6593
rect 11210 6579 11224 6593
rect 14210 6579 14224 6593
rect 14282 6579 14296 6593
rect 18962 6579 18976 6593
rect 23762 6579 23776 6593
rect 8258 6555 8272 6569
rect 17210 6555 17224 6569
rect 20522 6555 20536 6569
rect 22178 6555 22192 6569
rect 24314 6555 24328 6569
rect 25082 6555 25096 6569
rect 25346 6555 25360 6569
rect 8018 6531 8032 6545
rect 21530 6531 21544 6545
rect 25850 6531 25864 6545
rect 7778 6507 7792 6521
rect 7898 6507 7912 6521
rect 7994 6507 8008 6521
rect 26906 6507 26920 6521
rect 7730 6483 7744 6497
rect 25082 6483 25096 6497
rect 7706 6459 7720 6473
rect 16538 6459 16552 6473
rect 17618 6459 17632 6473
rect 22130 6459 22144 6473
rect 7706 6435 7720 6449
rect 16850 6435 16864 6449
rect 17522 6435 17536 6449
rect 19730 6435 19744 6449
rect 23114 6435 23128 6449
rect 7658 6411 7672 6425
rect 12866 6411 12880 6425
rect 13130 6411 13144 6425
rect 13634 6411 13648 6425
rect 14162 6411 14176 6425
rect 20522 6411 20536 6425
rect 23618 6411 23632 6425
rect 7610 6387 7624 6401
rect 14366 6387 14380 6401
rect 14474 6387 14488 6401
rect 19346 6387 19360 6401
rect 7586 6363 7600 6377
rect 9506 6363 9520 6377
rect 12722 6363 12736 6377
rect 12914 6363 12928 6377
rect 20090 6363 20104 6377
rect 25202 6363 25216 6377
rect 7226 6339 7240 6353
rect 8618 6339 8632 6353
rect 19106 6339 19120 6353
rect 22442 6339 22456 6353
rect 22826 6339 22840 6353
rect 7226 6315 7240 6329
rect 10658 6315 10672 6329
rect 10850 6315 10864 6329
rect 11570 6315 11584 6329
rect 17522 6315 17536 6329
rect 17618 6315 17632 6329
rect 18722 6315 18736 6329
rect 7178 6291 7192 6305
rect 20498 6291 20512 6305
rect 22202 6291 22216 6305
rect 7154 6267 7168 6281
rect 15218 6267 15232 6281
rect 7058 6243 7072 6257
rect 7250 6243 7264 6257
rect 13370 6243 13384 6257
rect 19082 6243 19096 6257
rect 22850 6243 22864 6257
rect 6938 6219 6952 6233
rect 16946 6219 16960 6233
rect 6914 6195 6928 6209
rect 22682 6195 22696 6209
rect 6866 6171 6880 6185
rect 12674 6171 12688 6185
rect 12890 6171 12904 6185
rect 18818 6171 18832 6185
rect 19010 6171 19024 6185
rect 20882 6171 20896 6185
rect 24338 6171 24352 6185
rect 27074 6171 27088 6185
rect 6842 6147 6856 6161
rect 9842 6147 9856 6161
rect 10346 6147 10360 6161
rect 14834 6147 14848 6161
rect 18506 6147 18520 6161
rect 23930 6147 23944 6161
rect 26066 6147 26080 6161
rect 26666 6147 26680 6161
rect 6458 6123 6472 6137
rect 22250 6123 22264 6137
rect 6314 6099 6328 6113
rect 21242 6099 21256 6113
rect 23042 6099 23056 6113
rect 23138 6099 23152 6113
rect 23210 6099 23224 6113
rect 23282 6099 23296 6113
rect 6218 6075 6232 6089
rect 9266 6075 9280 6089
rect 10946 6075 10960 6089
rect 16862 6075 16876 6089
rect 21338 6075 21352 6089
rect 22418 6075 22432 6089
rect 25754 6075 25768 6089
rect 6170 6051 6184 6065
rect 25298 6051 25312 6065
rect 6122 6027 6136 6041
rect 6362 6027 6376 6041
rect 6794 6027 6808 6041
rect 7442 6027 7456 6041
rect 10298 6027 10312 6041
rect 14714 6027 14728 6041
rect 19178 6027 19192 6041
rect 21266 6027 21280 6041
rect 23042 6027 23056 6041
rect 23066 6027 23080 6041
rect 23210 6027 23224 6041
rect 25778 6027 25792 6041
rect 26330 6027 26344 6041
rect 6026 6003 6040 6017
rect 11762 6003 11776 6017
rect 21602 6003 21616 6017
rect 22970 6003 22984 6017
rect 24410 6003 24424 6017
rect 5978 5979 5992 5993
rect 7370 5979 7384 5993
rect 7490 5979 7504 5993
rect 8474 5979 8488 5993
rect 10034 5979 10048 5993
rect 11330 5979 11344 5993
rect 13346 5979 13360 5993
rect 14258 5979 14272 5993
rect 20402 5979 20416 5993
rect 22970 5979 22984 5993
rect 23450 5979 23464 5993
rect 5930 5955 5944 5969
rect 7922 5955 7936 5969
rect 10394 5955 10408 5969
rect 10922 5955 10936 5969
rect 12770 5955 12784 5969
rect 13586 5955 13600 5969
rect 21338 5955 21352 5969
rect 24842 5955 24856 5969
rect 25994 5955 26008 5969
rect 5714 5931 5728 5945
rect 10010 5931 10024 5945
rect 10322 5931 10336 5945
rect 23186 5931 23200 5945
rect 5642 5907 5656 5921
rect 20786 5907 20800 5921
rect 22658 5907 22672 5921
rect 5354 5883 5368 5897
rect 5378 5883 5392 5897
rect 9962 5883 9976 5897
rect 19826 5883 19840 5897
rect 25130 5883 25144 5897
rect 5306 5859 5320 5873
rect 16994 5859 17008 5873
rect 5258 5835 5272 5849
rect 7010 5835 7024 5849
rect 24890 5835 24904 5849
rect 5210 5811 5224 5825
rect 14474 5811 14488 5825
rect 14522 5811 14536 5825
rect 21566 5811 21580 5825
rect 25178 5811 25192 5825
rect 25442 5811 25456 5825
rect 5186 5787 5200 5801
rect 10874 5787 10888 5801
rect 13874 5787 13888 5801
rect 13922 5787 13936 5801
rect 14306 5787 14320 5801
rect 14450 5787 14464 5801
rect 25178 5787 25192 5801
rect 5090 5763 5104 5777
rect 17474 5763 17488 5777
rect 5042 5739 5056 5753
rect 23162 5739 23176 5753
rect 5018 5715 5032 5729
rect 6602 5715 6616 5729
rect 6746 5715 6760 5729
rect 8906 5715 8920 5729
rect 9002 5715 9016 5729
rect 20186 5715 20200 5729
rect 23570 5715 23584 5729
rect 23594 5715 23608 5729
rect 4994 5691 5008 5705
rect 13850 5691 13864 5705
rect 13922 5691 13936 5705
rect 16682 5691 16696 5705
rect 20234 5691 20248 5705
rect 20690 5691 20704 5705
rect 20882 5691 20896 5705
rect 21674 5691 21688 5705
rect 23570 5691 23584 5705
rect 4922 5667 4936 5681
rect 15746 5667 15760 5681
rect 16346 5667 16360 5681
rect 18830 5667 18844 5681
rect 19898 5667 19912 5681
rect 20762 5667 20776 5681
rect 23858 5667 23872 5681
rect 4850 5643 4864 5657
rect 8186 5643 8200 5657
rect 8930 5643 8944 5657
rect 11258 5643 11272 5657
rect 15530 5643 15544 5657
rect 18578 5643 18592 5657
rect 18794 5643 18808 5657
rect 24842 5643 24856 5657
rect 4802 5619 4816 5633
rect 6482 5619 6496 5633
rect 6530 5619 6544 5633
rect 13778 5619 13792 5633
rect 13946 5619 13960 5633
rect 17306 5619 17320 5633
rect 4754 5595 4768 5609
rect 24794 5595 24808 5609
rect 4706 5571 4720 5585
rect 9050 5571 9064 5585
rect 9218 5571 9232 5585
rect 9626 5571 9640 5585
rect 9770 5571 9784 5585
rect 22490 5571 22504 5585
rect 4658 5547 4672 5561
rect 10370 5547 10384 5561
rect 16298 5547 16312 5561
rect 4658 5523 4672 5537
rect 7802 5523 7816 5537
rect 7874 5523 7888 5537
rect 12098 5523 12112 5537
rect 14450 5523 14464 5537
rect 16922 5523 16936 5537
rect 25562 5523 25576 5537
rect 4610 5499 4624 5513
rect 26210 5499 26224 5513
rect 4490 5475 4504 5489
rect 11786 5475 11800 5489
rect 21578 5475 21592 5489
rect 4490 5451 4504 5465
rect 16370 5451 16384 5465
rect 16754 5451 16768 5465
rect 26738 5451 26752 5465
rect 4442 5427 4456 5441
rect 8030 5427 8044 5441
rect 10538 5427 10552 5441
rect 13682 5427 13696 5441
rect 17402 5427 17416 5441
rect 23426 5427 23440 5441
rect 4370 5403 4384 5417
rect 18242 5403 18256 5417
rect 19274 5403 19288 5417
rect 25226 5403 25240 5417
rect 4370 5379 4384 5393
rect 8450 5379 8464 5393
rect 8498 5379 8512 5393
rect 23282 5379 23296 5393
rect 4346 5355 4360 5369
rect 9650 5355 9664 5369
rect 16490 5355 16504 5369
rect 17186 5355 17200 5369
rect 4298 5331 4312 5345
rect 14570 5331 14584 5345
rect 14858 5331 14872 5345
rect 16130 5331 16144 5345
rect 16514 5331 16528 5345
rect 16766 5331 16780 5345
rect 4274 5307 4288 5321
rect 17570 5307 17584 5321
rect 4250 5283 4264 5297
rect 7298 5283 7312 5297
rect 7346 5283 7360 5297
rect 12602 5283 12616 5297
rect 12650 5283 12664 5297
rect 13946 5283 13960 5297
rect 14234 5283 14248 5297
rect 14426 5283 14440 5297
rect 14498 5283 14512 5297
rect 14546 5283 14560 5297
rect 14618 5283 14632 5297
rect 24074 5283 24088 5297
rect 4226 5259 4240 5273
rect 8978 5259 8992 5273
rect 9026 5259 9040 5273
rect 22802 5259 22816 5273
rect 4202 5235 4216 5249
rect 9050 5235 9064 5249
rect 9098 5235 9112 5249
rect 17282 5235 17296 5249
rect 17450 5235 17464 5249
rect 17714 5235 17728 5249
rect 19034 5235 19048 5249
rect 19922 5235 19936 5249
rect 22058 5235 22072 5249
rect 4154 5211 4168 5225
rect 17642 5211 17656 5225
rect 18938 5211 18952 5225
rect 20498 5211 20512 5225
rect 21650 5211 21664 5225
rect 4130 5187 4144 5201
rect 5090 5187 5104 5201
rect 11450 5187 11464 5201
rect 14234 5187 14248 5201
rect 14402 5187 14416 5201
rect 20642 5187 20656 5201
rect 4034 5163 4048 5177
rect 5354 5163 5368 5177
rect 10226 5163 10240 5177
rect 11666 5163 11680 5177
rect 17738 5163 17752 5177
rect 18530 5163 18544 5177
rect 20282 5163 20296 5177
rect 21146 5163 21160 5177
rect 21494 5163 21508 5177
rect 4010 5139 4024 5153
rect 6650 5139 6664 5153
rect 6698 5139 6712 5153
rect 9098 5139 9112 5153
rect 12698 5139 12712 5153
rect 12770 5139 12784 5153
rect 26690 5139 26704 5153
rect 3938 5115 3952 5129
rect 10490 5115 10504 5129
rect 10610 5115 10624 5129
rect 10670 5115 10684 5129
rect 10706 5115 10720 5129
rect 21818 5115 21832 5129
rect 3914 5091 3928 5105
rect 5522 5091 5536 5105
rect 5570 5091 5584 5105
rect 8006 5091 8020 5105
rect 11474 5091 11488 5105
rect 14498 5091 14512 5105
rect 18002 5091 18016 5105
rect 18146 5091 18160 5105
rect 19922 5091 19936 5105
rect 24122 5091 24136 5105
rect 24194 5091 24208 5105
rect 3866 5067 3880 5081
rect 13466 5067 13480 5081
rect 13730 5067 13744 5081
rect 21938 5067 21952 5081
rect 24722 5067 24736 5081
rect 25394 5067 25408 5081
rect 3842 5043 3856 5057
rect 15242 5043 15256 5057
rect 16274 5043 16288 5057
rect 25274 5043 25288 5057
rect 25826 5043 25840 5057
rect 25862 5043 25876 5057
rect 3698 5019 3712 5033
rect 5426 5019 5440 5033
rect 15962 5019 15976 5033
rect 26234 5019 26248 5033
rect 3650 4995 3664 5009
rect 4586 4995 4600 5009
rect 9026 4995 9040 5009
rect 10082 4995 10096 5009
rect 10898 4995 10912 5009
rect 11138 4995 11152 5009
rect 16322 4995 16336 5009
rect 16514 4995 16528 5009
rect 24938 4995 24952 5009
rect 25238 4995 25252 5009
rect 25826 4995 25840 5009
rect 26594 4995 26608 5009
rect 3578 4971 3592 4985
rect 17450 4971 17464 4985
rect 23714 4971 23728 4985
rect 3554 4947 3568 4961
rect 21146 4947 21160 4961
rect 3482 4923 3496 4937
rect 13106 4923 13120 4937
rect 14282 4923 14296 4937
rect 14330 4923 14344 4937
rect 24050 4923 24064 4937
rect 3458 4899 3472 4913
rect 6458 4899 6472 4913
rect 7850 4899 7864 4913
rect 8786 4899 8800 4913
rect 9218 4899 9232 4913
rect 9866 4899 9880 4913
rect 11522 4899 11536 4913
rect 23642 4899 23656 4913
rect 23978 4899 23992 4913
rect 24626 4899 24640 4913
rect 24890 4899 24904 4913
rect 3410 4875 3424 4889
rect 17498 4875 17512 4889
rect 21050 4875 21064 4889
rect 3386 4851 3400 4865
rect 9338 4851 9352 4865
rect 13994 4851 14008 4865
rect 21122 4851 21136 4865
rect 23690 4851 23704 4865
rect 3290 4827 3304 4841
rect 3770 4827 3784 4841
rect 7634 4827 7648 4841
rect 8954 4827 8968 4841
rect 9386 4827 9400 4841
rect 11378 4827 11392 4841
rect 20330 4827 20344 4841
rect 20954 4827 20968 4841
rect 21098 4827 21112 4841
rect 3266 4803 3280 4817
rect 19658 4803 19672 4817
rect 20810 4803 20824 4817
rect 21626 4803 21640 4817
rect 3242 4779 3256 4793
rect 13370 4779 13384 4793
rect 13514 4779 13528 4793
rect 13658 4779 13672 4793
rect 13994 4779 14008 4793
rect 14114 4779 14128 4793
rect 19706 4779 19720 4793
rect 20258 4779 20272 4793
rect 20450 4779 20464 4793
rect 20618 4779 20632 4793
rect 21410 4779 21424 4793
rect 3218 4755 3232 4769
rect 7970 4755 7984 4769
rect 16274 4755 16288 4769
rect 18410 4755 18424 4769
rect 20354 4755 20368 4769
rect 20546 4755 20560 4769
rect 21494 4755 21508 4769
rect 3170 4731 3184 4745
rect 9986 4731 10000 4745
rect 10274 4731 10288 4745
rect 15098 4731 15112 4745
rect 19514 4731 19528 4745
rect 19610 4731 19624 4745
rect 22706 4731 22720 4745
rect 25346 4731 25360 4745
rect 3122 4707 3136 4721
rect 8162 4707 8176 4721
rect 11930 4707 11944 4721
rect 12194 4707 12208 4721
rect 22946 4707 22960 4721
rect 3026 4683 3040 4697
rect 24434 4683 24448 4697
rect 3002 4659 3016 4673
rect 17042 4659 17056 4673
rect 17090 4659 17104 4673
rect 26786 4659 26800 4673
rect 2978 4635 2992 4649
rect 6074 4635 6088 4649
rect 6122 4635 6136 4649
rect 7130 4635 7144 4649
rect 19850 4635 19864 4649
rect 20162 4635 20176 4649
rect 24314 4635 24328 4649
rect 2906 4611 2920 4625
rect 6146 4611 6160 4625
rect 9146 4611 9160 4625
rect 13610 4611 13624 4625
rect 15482 4611 15496 4625
rect 18890 4611 18904 4625
rect 24506 4611 24520 4625
rect 2882 4587 2896 4601
rect 5282 4587 5296 4601
rect 5330 4587 5344 4601
rect 17330 4587 17344 4601
rect 18482 4587 18496 4601
rect 18626 4587 18640 4601
rect 18866 4587 18880 4601
rect 19154 4587 19168 4601
rect 19202 4587 19216 4601
rect 22262 4587 22276 4601
rect 2858 4563 2872 4577
rect 12914 4563 12928 4577
rect 21554 4563 21568 4577
rect 2810 4539 2824 4553
rect 6506 4539 6520 4553
rect 6698 4539 6712 4553
rect 19778 4539 19792 4553
rect 19970 4539 19984 4553
rect 23450 4539 23464 4553
rect 2738 4515 2752 4529
rect 21194 4515 21208 4529
rect 22082 4515 22096 4529
rect 22142 4515 22156 4529
rect 2666 4491 2680 4505
rect 4586 4491 4600 4505
rect 4682 4491 4696 4505
rect 6626 4491 6640 4505
rect 13226 4491 13240 4505
rect 16250 4491 16264 4505
rect 21002 4491 21016 4505
rect 21314 4491 21328 4505
rect 22874 4491 22888 4505
rect 23786 4491 23800 4505
rect 2642 4467 2656 4481
rect 6578 4467 6592 4481
rect 7778 4467 7792 4481
rect 9578 4467 9592 4481
rect 23306 4467 23320 4481
rect 2594 4443 2608 4457
rect 11690 4443 11704 4457
rect 11738 4443 11752 4457
rect 17138 4443 17152 4457
rect 17810 4443 17824 4457
rect 26570 4443 26584 4457
rect 2570 4419 2584 4433
rect 4514 4419 4528 4433
rect 23186 4419 23200 4433
rect 24362 4419 24376 4433
rect 24578 4419 24592 4433
rect 26138 4419 26152 4433
rect 26378 4419 26392 4433
rect 2546 4395 2560 4409
rect 5762 4395 5776 4409
rect 5834 4395 5848 4409
rect 16766 4395 16780 4409
rect 21194 4395 21208 4409
rect 22226 4395 22240 4409
rect 22298 4395 22312 4409
rect 23330 4395 23344 4409
rect 23498 4395 23512 4409
rect 24218 4395 24232 4409
rect 25610 4395 25624 4409
rect 26042 4395 26056 4409
rect 26162 4395 26176 4409
rect 26306 4395 26320 4409
rect 26474 4395 26488 4409
rect 26522 4395 26536 4409
rect 26882 4395 26896 4409
rect 2522 4371 2536 4385
rect 15338 4371 15352 4385
rect 21746 4371 21760 4385
rect 24026 4371 24040 4385
rect 24098 4371 24112 4385
rect 24446 4371 24460 4385
rect 24674 4371 24688 4385
rect 26762 4371 26776 4385
rect 2498 4347 2512 4361
rect 9554 4347 9568 4361
rect 11426 4347 11440 4361
rect 15314 4347 15328 4361
rect 25058 4347 25072 4361
rect 25106 4347 25120 4361
rect 27266 4347 27280 4361
rect 2426 4323 2440 4337
rect 14642 4323 14656 4337
rect 22082 4323 22096 4337
rect 22418 4323 22432 4337
rect 22562 4323 22576 4337
rect 22610 4323 22624 4337
rect 22754 4323 22768 4337
rect 22922 4323 22936 4337
rect 23114 4323 23128 4337
rect 26930 4323 26944 4337
rect 2330 4299 2344 4313
rect 8666 4299 8680 4313
rect 8786 4299 8800 4313
rect 19826 4299 19840 4313
rect 23810 4299 23824 4313
rect 24866 4299 24880 4313
rect 25058 4299 25072 4313
rect 25238 4299 25252 4313
rect 25994 4299 26008 4313
rect 26066 4299 26080 4313
rect 2234 4275 2248 4289
rect 9530 4275 9544 4289
rect 9602 4275 9616 4289
rect 27314 4275 27328 4289
rect 2234 4251 2248 4265
rect 20378 4251 20392 4265
rect 21482 4251 21496 4265
rect 25634 4251 25648 4265
rect 2186 4227 2200 4241
rect 7418 4227 7432 4241
rect 7490 4227 7504 4241
rect 26186 4227 26200 4241
rect 26330 4227 26344 4241
rect 2114 4203 2128 4217
rect 20714 4203 20728 4217
rect 22634 4203 22648 4217
rect 23306 4203 23320 4217
rect 23426 4203 23440 4217
rect 23474 4203 23488 4217
rect 26354 4203 26368 4217
rect 2066 4179 2080 4193
rect 8210 4179 8224 4193
rect 20258 4179 20272 4193
rect 20306 4179 20320 4193
rect 22898 4179 22912 4193
rect 23858 4179 23872 4193
rect 23930 4179 23944 4193
rect 1994 4155 2008 4169
rect 11858 4155 11872 4169
rect 12794 4155 12808 4169
rect 13394 4155 13408 4169
rect 13562 4155 13576 4169
rect 17690 4155 17704 4169
rect 17978 4155 17992 4169
rect 19130 4155 19144 4169
rect 19850 4155 19864 4169
rect 20186 4155 20200 4169
rect 21866 4155 21880 4169
rect 23354 4155 23368 4169
rect 1946 4131 1960 4145
rect 2690 4131 2704 4145
rect 3986 4131 4000 4145
rect 4034 4131 4048 4145
rect 4058 4131 4072 4145
rect 4106 4131 4120 4145
rect 8642 4131 8656 4145
rect 12146 4131 12160 4145
rect 12218 4131 12232 4145
rect 12602 4131 12616 4145
rect 12650 4131 12664 4145
rect 14090 4131 14104 4145
rect 26042 4131 26056 4145
rect 1898 4107 1912 4121
rect 3746 4107 3760 4121
rect 9410 4107 9424 4121
rect 9458 4107 9472 4121
rect 26714 4107 26728 4121
rect 1850 4083 1864 4097
rect 7394 4083 7408 4097
rect 26234 4083 26248 4097
rect 1826 4059 1840 4073
rect 13418 4059 13432 4073
rect 13610 4059 13624 4073
rect 14210 4059 14224 4073
rect 14978 4059 14992 4073
rect 27026 4059 27040 4073
rect 1658 4035 1672 4049
rect 2498 4035 2512 4049
rect 7274 4035 7288 4049
rect 10202 4035 10216 4049
rect 10298 4035 10312 4049
rect 10346 4035 10360 4049
rect 10418 4035 10432 4049
rect 10466 4035 10480 4049
rect 10634 4035 10648 4049
rect 12290 4035 12304 4049
rect 22442 4035 22456 4049
rect 22538 4035 22552 4049
rect 23138 4035 23152 4049
rect 27122 4035 27136 4049
rect 1610 4011 1624 4025
rect 6482 4011 6496 4025
rect 8234 4011 8248 4025
rect 11354 4011 11368 4025
rect 22106 4011 22120 4025
rect 26426 4011 26440 4025
rect 70 3987 84 4001
rect 10610 3987 10624 4001
rect 24554 3987 24568 4001
rect 26426 3987 26440 4001
rect 27194 3987 27208 4001
rect 70 3963 84 3977
rect 6746 3963 6760 3977
rect 6818 3963 6832 3977
rect 9194 3963 9208 3977
rect 10058 3963 10072 3977
rect 12578 3963 12592 3977
rect 13202 3963 13216 3977
rect 23354 3963 23368 3977
rect 1730 3939 1744 3953
rect 2786 3939 2800 3953
rect 2834 3939 2848 3953
rect 4274 3939 4288 3953
rect 20594 3939 20608 3953
rect 22142 3939 22156 3953
rect 22226 3939 22240 3953
rect 22262 3939 22276 3953
rect 22298 3939 22312 3953
rect 23258 3939 23272 3953
rect 1778 3915 1792 3929
rect 9482 3915 9496 3929
rect 9530 3915 9544 3929
rect 9842 3915 9856 3929
rect 9986 3915 10000 3929
rect 15266 3915 15280 3929
rect 24266 3915 24280 3929
rect 2042 3891 2056 3905
rect 4802 3891 4816 3905
rect 6338 3891 6352 3905
rect 24962 3891 24976 3905
rect 2090 3867 2104 3881
rect 2306 3867 2320 3881
rect 3674 3867 3688 3881
rect 7058 3867 7072 3881
rect 7370 3867 7384 3881
rect 15434 3867 15448 3881
rect 16610 3867 16624 3881
rect 16706 3867 16720 3881
rect 18434 3867 18448 3881
rect 23066 3867 23080 3881
rect 23330 3867 23344 3881
rect 26306 3867 26320 3881
rect 2282 3843 2296 3857
rect 8210 3843 8224 3857
rect 10754 3843 10768 3857
rect 11618 3843 11632 3857
rect 13154 3843 13168 3857
rect 26618 3843 26632 3857
rect 2306 3819 2320 3833
rect 8690 3819 8704 3833
rect 9314 3819 9328 3833
rect 11234 3819 11248 3833
rect 13274 3819 13288 3833
rect 14330 3819 14344 3833
rect 15458 3819 15472 3833
rect 15986 3819 16000 3833
rect 16562 3819 16576 3833
rect 18770 3819 18784 3833
rect 20018 3819 20032 3833
rect 22754 3819 22768 3833
rect 23546 3819 23560 3833
rect 23666 3819 23680 3833
rect 26402 3819 26416 3833
rect 2354 3795 2368 3809
rect 15986 3795 16000 3809
rect 16106 3795 16120 3809
rect 22994 3795 23008 3809
rect 2354 3771 2368 3785
rect 4466 3771 4480 3785
rect 5474 3771 5488 3785
rect 7394 3771 7408 3785
rect 13658 3771 13672 3785
rect 23090 3771 23104 3785
rect 25802 3771 25816 3785
rect 2402 3747 2416 3761
rect 8066 3747 8080 3761
rect 8114 3747 8128 3761
rect 8258 3747 8272 3761
rect 13898 3747 13912 3761
rect 14882 3747 14896 3761
rect 15194 3747 15208 3761
rect 20666 3747 20680 3761
rect 22946 3747 22960 3761
rect 2402 3723 2416 3737
rect 5498 3723 5512 3737
rect 5954 3723 5968 3737
rect 12866 3723 12880 3737
rect 17786 3723 17800 3737
rect 20042 3723 20056 3737
rect 22562 3723 22576 3737
rect 2426 3699 2440 3713
rect 2858 3699 2872 3713
rect 6050 3699 6064 3713
rect 9242 3699 9256 3713
rect 10994 3699 11008 3713
rect 11402 3699 11416 3713
rect 15770 3699 15784 3713
rect 19226 3699 19240 3713
rect 20930 3699 20944 3713
rect 25922 3699 25936 3713
rect 2450 3675 2464 3689
rect 12746 3675 12760 3689
rect 12818 3675 12832 3689
rect 12962 3675 12976 3689
rect 13154 3675 13168 3689
rect 26858 3675 26872 3689
rect 2450 3651 2464 3665
rect 26498 3651 26512 3665
rect 2522 3627 2536 3641
rect 5594 3627 5608 3641
rect 6818 3627 6832 3641
rect 10418 3627 10432 3641
rect 16586 3627 16600 3641
rect 16730 3627 16744 3641
rect 18314 3627 18328 3641
rect 25490 3627 25504 3641
rect 2618 3603 2632 3617
rect 5066 3603 5080 3617
rect 26138 3603 26152 3617
rect 2642 3579 2656 3593
rect 7946 3579 7960 3593
rect 11030 3579 11044 3593
rect 11114 3579 11128 3593
rect 20618 3579 20632 3593
rect 21986 3579 22000 3593
rect 26450 3579 26464 3593
rect 2666 3555 2680 3569
rect 15410 3555 15424 3569
rect 15458 3555 15472 3569
rect 15530 3555 15544 3569
rect 15626 3555 15640 3569
rect 16394 3555 16408 3569
rect 16586 3555 16600 3569
rect 16970 3555 16984 3569
rect 17474 3555 17488 3569
rect 17762 3555 17776 3569
rect 18050 3555 18064 3569
rect 26834 3555 26848 3569
rect 2714 3531 2728 3545
rect 24362 3531 24376 3545
rect 26474 3531 26488 3545
rect 2738 3507 2752 3521
rect 5450 3507 5464 3521
rect 6386 3507 6400 3521
rect 6410 3507 6424 3521
rect 16226 3507 16240 3521
rect 26210 3507 26224 3521
rect 2762 3483 2776 3497
rect 16442 3483 16456 3497
rect 16658 3483 16672 3497
rect 26978 3483 26992 3497
rect 3002 3459 3016 3473
rect 25658 3459 25672 3473
rect 3050 3435 3064 3449
rect 18914 3435 18928 3449
rect 19010 3435 19024 3449
rect 19346 3435 19360 3449
rect 19994 3435 20008 3449
rect 26162 3435 26176 3449
rect 3074 3411 3088 3425
rect 9746 3411 9760 3425
rect 10058 3411 10072 3425
rect 21290 3411 21304 3425
rect 3146 3387 3160 3401
rect 3554 3387 3568 3401
rect 3602 3387 3616 3401
rect 24170 3387 24184 3401
rect 3314 3363 3328 3377
rect 26762 3363 26776 3377
rect 3362 3339 3376 3353
rect 20834 3339 20848 3353
rect 3362 3315 3376 3329
rect 8450 3315 8464 3329
rect 9794 3315 9808 3329
rect 14066 3315 14080 3329
rect 14594 3315 14608 3329
rect 17546 3315 17560 3329
rect 18482 3315 18496 3329
rect 18602 3315 18616 3329
rect 19946 3315 19960 3329
rect 20138 3315 20152 3329
rect 3410 3291 3424 3305
rect 8138 3291 8152 3305
rect 8858 3291 8872 3305
rect 9890 3291 9904 3305
rect 18674 3291 18688 3305
rect 21458 3291 21472 3305
rect 22610 3291 22624 3305
rect 3506 3267 3520 3281
rect 22874 3267 22888 3281
rect 3602 3243 3616 3257
rect 7610 3243 7624 3257
rect 15866 3243 15880 3257
rect 16634 3243 16648 3257
rect 16706 3243 16720 3257
rect 16862 3243 16876 3257
rect 18746 3243 18760 3257
rect 25418 3243 25432 3257
rect 3626 3219 3640 3233
rect 6914 3219 6928 3233
rect 13706 3219 13720 3233
rect 16466 3219 16480 3233
rect 16802 3219 16816 3233
rect 26114 3219 26128 3233
rect 3746 3195 3760 3209
rect 17234 3195 17248 3209
rect 18770 3195 18784 3209
rect 18830 3195 18844 3209
rect 18890 3195 18904 3209
rect 19274 3195 19288 3209
rect 20018 3195 20032 3209
rect 20354 3195 20368 3209
rect 25418 3195 25432 3209
rect 26258 3195 26272 3209
rect 3770 3171 3784 3185
rect 20210 3171 20224 3185
rect 3794 3147 3808 3161
rect 26810 3147 26824 3161
rect 3842 3123 3856 3137
rect 6938 3123 6952 3137
rect 9818 3123 9832 3137
rect 13754 3123 13768 3137
rect 15890 3123 15904 3137
rect 16826 3123 16840 3137
rect 18554 3123 18568 3137
rect 18818 3123 18832 3137
rect 26954 3123 26968 3137
rect 3866 3099 3880 3113
rect 8882 3099 8896 3113
rect 9674 3099 9688 3113
rect 16034 3099 16048 3113
rect 17666 3099 17680 3113
rect 18458 3099 18472 3113
rect 20738 3099 20752 3113
rect 20978 3099 20992 3113
rect 22922 3099 22936 3113
rect 3890 3075 3904 3089
rect 14522 3075 14536 3089
rect 15218 3075 15232 3089
rect 17018 3075 17032 3089
rect 18098 3075 18112 3089
rect 19322 3075 19336 3089
rect 23402 3075 23416 3089
rect 24650 3075 24664 3089
rect 25442 3075 25456 3089
rect 25514 3075 25528 3089
rect 3914 3051 3928 3065
rect 4778 3051 4792 3065
rect 7730 3051 7744 3065
rect 9626 3051 9640 3065
rect 12962 3051 12976 3065
rect 16202 3051 16216 3065
rect 17714 3051 17728 3065
rect 18578 3051 18592 3065
rect 19082 3051 19096 3065
rect 20714 3051 20728 3065
rect 3938 3027 3952 3041
rect 5810 3027 5824 3041
rect 5882 3027 5896 3041
rect 25370 3027 25384 3041
rect 4010 3003 4024 3017
rect 11306 3003 11320 3017
rect 12386 3003 12400 3017
rect 18650 3003 18664 3017
rect 20210 3003 20224 3017
rect 20402 3003 20416 3017
rect 20738 3003 20752 3017
rect 21578 3003 21592 3017
rect 4106 2979 4120 2993
rect 6554 2979 6568 2993
rect 6674 2979 6688 2993
rect 11882 2979 11896 2993
rect 12242 2979 12256 2993
rect 14546 2979 14560 2993
rect 15386 2979 15400 2993
rect 16178 2979 16192 2993
rect 16226 2979 16240 2993
rect 16298 2979 16312 2993
rect 16730 2979 16744 2993
rect 17066 2979 17080 2993
rect 18458 2979 18472 2993
rect 20906 2979 20920 2993
rect 4130 2955 4144 2969
rect 6554 2955 6568 2969
rect 21386 2955 21400 2969
rect 26090 2955 26104 2969
rect 4202 2931 4216 2945
rect 9722 2931 9736 2945
rect 12074 2931 12088 2945
rect 13082 2931 13096 2945
rect 13322 2931 13336 2945
rect 13826 2931 13840 2945
rect 18362 2931 18376 2945
rect 18866 2931 18880 2945
rect 21218 2931 21232 2945
rect 22538 2931 22552 2945
rect 24098 2931 24112 2945
rect 4226 2907 4240 2921
rect 4874 2907 4888 2921
rect 6794 2907 6808 2921
rect 7466 2907 7480 2921
rect 7634 2907 7648 2921
rect 7826 2907 7840 2921
rect 8834 2907 8848 2921
rect 10178 2907 10192 2921
rect 17114 2907 17128 2921
rect 21026 2907 21040 2921
rect 4394 2883 4408 2897
rect 10082 2883 10096 2897
rect 10322 2883 10336 2897
rect 11546 2883 11560 2897
rect 11594 2883 11608 2897
rect 27651 2883 27665 2897
rect 4418 2859 4432 2873
rect 14138 2859 14152 2873
rect 22346 2859 22360 2873
rect 4442 2835 4456 2849
rect 14114 2835 14128 2849
rect 16394 2835 16408 2849
rect 19058 2835 19072 2849
rect 24746 2835 24760 2849
rect 26378 2835 26392 2849
rect 4562 2811 4576 2825
rect 17546 2811 17560 2825
rect 4682 2787 4696 2801
rect 11810 2787 11824 2801
rect 12338 2787 12352 2801
rect 21434 2787 21448 2801
rect 24446 2787 24460 2801
rect 4778 2763 4792 2777
rect 6266 2763 6280 2777
rect 18626 2763 18640 2777
rect 4874 2739 4888 2753
rect 6722 2739 6736 2753
rect 15506 2739 15520 2753
rect 15554 2739 15568 2753
rect 20066 2739 20080 2753
rect 22178 2739 22192 2753
rect 4922 2715 4936 2729
rect 10970 2715 10984 2729
rect 13490 2715 13504 2729
rect 14066 2715 14080 2729
rect 14366 2715 14380 2729
rect 15482 2715 15496 2729
rect 23234 2715 23248 2729
rect 4970 2691 4984 2705
rect 25274 2691 25288 2705
rect 4994 2667 5008 2681
rect 5474 2667 5488 2681
rect 9170 2667 9184 2681
rect 11714 2667 11728 2681
rect 14570 2667 14584 2681
rect 25862 2667 25876 2681
rect 5138 2643 5152 2657
rect 13298 2643 13312 2657
rect 16898 2643 16912 2657
rect 21410 2643 21424 2657
rect 25730 2643 25744 2657
rect 5162 2619 5176 2633
rect 21266 2619 21280 2633
rect 5210 2595 5224 2609
rect 8738 2595 8752 2609
rect 14690 2595 14704 2609
rect 26282 2595 26296 2609
rect 5306 2571 5320 2585
rect 9914 2571 9928 2585
rect 10826 2571 10840 2585
rect 14810 2571 14824 2585
rect 19154 2571 19168 2585
rect 5402 2547 5416 2561
rect 26498 2547 26512 2561
rect 5570 2523 5584 2537
rect 9698 2523 9712 2537
rect 9770 2523 9784 2537
rect 19370 2523 19384 2537
rect 5594 2499 5608 2513
rect 12506 2499 12520 2513
rect 12554 2499 12568 2513
rect 25322 2499 25336 2513
rect 5690 2475 5704 2489
rect 10106 2475 10120 2489
rect 10442 2475 10456 2489
rect 24386 2475 24400 2489
rect 6074 2451 6088 2465
rect 24290 2451 24304 2465
rect 6290 2427 6304 2441
rect 6722 2427 6736 2441
rect 10154 2427 10168 2441
rect 11162 2427 11176 2441
rect 22586 2427 22600 2441
rect 6362 2403 6376 2417
rect 10730 2403 10744 2417
rect 15578 2403 15592 2417
rect 20114 2403 20128 2417
rect 6506 2379 6520 2393
rect 9458 2379 9472 2393
rect 19466 2379 19480 2393
rect 20810 2379 20824 2393
rect 6866 2355 6880 2369
rect 14354 2355 14368 2369
rect 18218 2355 18232 2369
rect 18386 2355 18400 2369
rect 6962 2331 6976 2345
rect 19802 2331 19816 2345
rect 6986 2307 7000 2321
rect 13874 2307 13888 2321
rect 14186 2307 14200 2321
rect 21170 2307 21184 2321
rect 21362 2307 21376 2321
rect 25226 2307 25240 2321
rect 7154 2283 7168 2297
rect 19250 2283 19264 2297
rect 7178 2259 7192 2273
rect 14042 2259 14056 2273
rect 14690 2259 14704 2273
rect 22730 2259 22744 2273
rect 24986 2259 25000 2273
rect 7250 2235 7264 2249
rect 24002 2235 24016 2249
rect 7274 2211 7288 2225
rect 20450 2211 20464 2225
rect 21626 2211 21640 2225
rect 7418 2187 7432 2201
rect 7442 2187 7456 2201
rect 7514 2187 7528 2201
rect 21890 2187 21904 2201
rect 7562 2163 7576 2177
rect 23738 2163 23752 2177
rect 7754 2139 7768 2153
rect 22346 2139 22360 2153
rect 7850 2115 7864 2129
rect 8006 2115 8020 2129
rect 8090 2115 8104 2129
rect 10466 2115 10480 2129
rect 26642 2115 26656 2129
rect 7946 2091 7960 2105
rect 8030 2091 8044 2105
rect 8162 2091 8176 2105
rect 8186 2091 8200 2105
rect 8282 2091 8296 2105
rect 14426 2091 14440 2105
rect 16178 2091 16192 2105
rect 25970 2091 25984 2105
rect 7970 2067 7984 2081
rect 25034 2067 25048 2081
rect 8018 2043 8032 2057
rect 13538 2043 13552 2057
rect 18986 2043 19000 2057
rect 19250 2043 19264 2057
rect 20474 2043 20488 2057
rect 25034 2043 25048 2057
rect 25202 2043 25216 2057
rect 8306 2019 8320 2033
rect 9434 2019 9448 2033
rect 22634 2019 22648 2033
rect 8354 1995 8368 2009
rect 8810 1995 8824 2009
rect 8954 1995 8968 2009
rect 8978 1995 8992 2009
rect 9074 1995 9088 2009
rect 18266 1995 18280 2009
rect 18986 1995 19000 2009
rect 19418 1995 19432 2009
rect 8378 1971 8392 1985
rect 8930 1971 8944 1985
rect 10670 1971 10684 1985
rect 23594 1971 23608 1985
rect 8570 1947 8584 1961
rect 12674 1947 12688 1961
rect 13010 1947 13024 1961
rect 13802 1947 13816 1961
rect 16418 1947 16432 1961
rect 21242 1947 21256 1961
rect 23378 1947 23392 1961
rect 24482 1947 24496 1961
rect 26642 1947 26656 1961
rect 8594 1923 8608 1937
rect 26522 1923 26536 1937
rect 8762 1899 8776 1913
rect 9362 1899 9376 1913
rect 9554 1899 9568 1913
rect 10130 1899 10144 1913
rect 11834 1899 11848 1913
rect 17426 1899 17440 1913
rect 24530 1899 24544 1913
rect 9146 1875 9160 1889
rect 11642 1875 11656 1889
rect 11834 1875 11848 1889
rect 12026 1875 12040 1889
rect 12410 1875 12424 1889
rect 12890 1875 12904 1889
rect 13250 1875 13264 1889
rect 18362 1875 18376 1889
rect 23882 1875 23896 1889
rect 24074 1875 24088 1889
rect 26018 1875 26032 1889
rect 26618 1875 26632 1889
rect 9674 1851 9688 1865
rect 10034 1851 10048 1865
rect 10490 1851 10504 1865
rect 21050 1851 21064 1865
rect 26882 1851 26896 1865
rect 9818 1827 9832 1841
rect 19586 1827 19600 1841
rect 10826 1803 10840 1817
rect 10946 1803 10960 1817
rect 11018 1803 11032 1817
rect 20858 1803 20872 1817
rect 10922 1779 10936 1793
rect 27290 1779 27304 1793
rect 11162 1755 11176 1769
rect 11954 1755 11968 1769
rect 12458 1755 12472 1769
rect 13754 1755 13768 1769
rect 15650 1755 15664 1769
rect 20786 1755 20800 1769
rect 22850 1755 22864 1769
rect 23906 1755 23920 1769
rect 11186 1731 11200 1745
rect 14018 1731 14032 1745
rect 16010 1731 16024 1745
rect 25898 1731 25912 1745
rect 11234 1707 11248 1721
rect 27242 1707 27256 1721
rect 11306 1683 11320 1697
rect 13442 1683 13456 1697
rect 23498 1683 23512 1697
rect 24242 1683 24256 1697
rect 25154 1683 25168 1697
rect 11426 1659 11440 1673
rect 11474 1659 11488 1673
rect 12458 1659 12472 1673
rect 14306 1659 14320 1673
rect 16322 1659 16336 1673
rect 16490 1659 16504 1673
rect 23906 1659 23920 1673
rect 24410 1659 24424 1673
rect 25154 1659 25168 1673
rect 25394 1659 25408 1673
rect 13202 1635 13216 1649
rect 13634 1635 13648 1649
rect 27314 1635 27328 1649
rect 27651 1635 27665 1649
rect 13418 1611 13432 1625
rect 13970 1611 13984 1625
rect 27290 1611 27304 1625
rect 27651 1611 27665 1625
rect 13538 1587 13552 1601
rect 19298 1587 19312 1601
rect 24146 1587 24160 1601
rect 27266 1587 27280 1601
rect 27651 1587 27665 1601
rect 13250 754 13264 768
rect 15530 754 15544 768
rect 11930 730 11944 744
rect 20354 730 20368 744
rect 11522 706 11536 720
rect 19946 706 19960 720
rect 10370 682 10384 696
rect 21914 682 21928 696
rect 10274 658 10288 672
rect 19130 658 19144 672
rect 26114 658 26128 672
rect 9698 634 9712 648
rect 13586 634 13600 648
rect 13826 634 13840 648
rect 14930 634 14944 648
rect 16898 634 16912 648
rect 19658 634 19672 648
rect 9002 610 9016 624
rect 10202 610 10216 624
rect 11066 610 11080 624
rect 26186 610 26200 624
rect 8666 586 8680 600
rect 9914 586 9928 600
rect 10010 586 10024 600
rect 16058 586 16072 600
rect 16778 586 16792 600
rect 17642 586 17656 600
rect 18122 586 18136 600
rect 20042 586 20056 600
rect 21386 586 21400 600
rect 23954 586 23968 600
rect 8474 562 8488 576
rect 10658 562 10672 576
rect 11162 562 11176 576
rect 11258 562 11272 576
rect 16082 562 16096 576
rect 16490 562 16504 576
rect 22010 562 22024 576
rect 22586 562 22600 576
rect 23978 562 23992 576
rect 7982 538 7996 552
rect 12602 538 12616 552
rect 12794 538 12808 552
rect 18506 538 18520 552
rect 21098 538 21112 552
rect 22898 538 22912 552
rect 7874 514 7888 528
rect 14210 514 14224 528
rect 15026 514 15040 528
rect 15074 514 15088 528
rect 15362 514 15376 528
rect 23138 514 23152 528
rect 7562 490 7576 504
rect 9434 490 9448 504
rect 9602 490 9616 504
rect 26378 490 26392 504
rect 7514 466 7528 480
rect 15818 466 15832 480
rect 15914 466 15928 480
rect 21962 466 21976 480
rect 22130 466 22144 480
rect 26834 466 26848 480
rect 6650 442 6664 456
rect 13706 442 13720 456
rect 13778 442 13792 456
rect 14402 442 14416 456
rect 14954 442 14968 456
rect 20138 442 20152 456
rect 20546 442 20560 456
rect 22658 442 22672 456
rect 23258 442 23272 456
rect 23666 442 23680 456
rect 26810 442 26824 456
rect 26858 442 26872 456
rect 6410 418 6424 432
rect 7130 418 7144 432
rect 7322 418 7336 432
rect 24482 418 24496 432
rect 26762 418 26776 432
rect 27651 418 27665 432
rect 6266 394 6280 408
rect 10778 394 10792 408
rect 10874 394 10888 408
rect 15146 394 15160 408
rect 15290 394 15304 408
rect 23402 394 23416 408
rect 23906 394 23920 408
rect 26714 394 26728 408
rect 26810 394 26824 408
rect 5546 370 5560 384
rect 6602 370 6616 384
rect 17858 370 17872 384
rect 5258 346 5272 360
rect 7034 346 7048 360
rect 7082 346 7096 360
rect 20402 346 20416 360
rect 5234 322 5248 336
rect 8498 322 8512 336
rect 8546 322 8560 336
rect 14162 322 14176 336
rect 4730 298 4744 312
rect 11546 298 11560 312
rect 11714 298 11728 312
rect 23690 298 23704 312
rect 4466 274 4480 288
rect 18602 274 18616 288
rect 4346 250 4360 264
rect 4826 250 4840 264
rect 5018 250 5032 264
rect 26666 250 26680 264
rect 4322 226 4336 240
rect 9410 226 9424 240
rect 15698 226 15712 240
rect 4154 202 4168 216
rect 20594 202 20608 216
rect 4058 178 4072 192
rect 7298 178 7312 192
rect 7442 178 7456 192
rect 11642 178 11656 192
rect 11882 178 11896 192
rect 17690 178 17704 192
rect 3722 154 3736 168
rect 18170 154 18184 168
rect 3698 130 3712 144
rect 22994 130 23008 144
rect 3650 106 3664 120
rect 15002 106 15016 120
rect 1682 82 1696 96
rect 20450 82 20464 96
rect 70 58 84 72
rect 23498 58 23512 72
rect 26858 58 26872 72
rect 27651 58 27665 72
rect 70 34 84 48
rect 2234 34 2248 48
rect 2546 34 2560 48
rect 4538 34 4552 48
rect 22778 34 22792 48
rect 26810 34 26824 48
rect 27651 34 27665 48
rect 3554 10 3568 24
rect 14426 10 14440 24
rect 26834 10 26848 24
rect 27651 10 27665 24
<< metal2 >>
rect 0 8085 70 8097
rect 0 8061 70 8073
rect 123 7882 323 8204
rect 339 7882 351 8204
rect 363 7882 375 8204
rect 387 7882 399 8204
rect 411 7882 423 8204
rect 2427 8098 2439 8204
rect 1731 7882 1743 8084
rect 1779 7882 1791 8060
rect 2595 7882 2607 8060
rect 3291 8050 3303 8204
rect 4155 8026 4167 8204
rect 5007 8026 5019 8204
rect 5583 8122 5595 8204
rect 5584 8108 5602 8122
rect 5008 8012 5026 8026
rect 4779 7882 4791 8012
rect 4995 7882 5007 8012
rect 5115 7882 5127 8012
rect 5379 7882 5391 7988
rect 5571 7882 5583 8108
rect 5595 7882 5607 7964
rect 5715 7882 5727 8108
rect 6747 7954 6759 8204
rect 6783 7978 6795 8204
rect 7659 7882 7671 7964
rect 8043 7882 8055 8132
rect 8475 7930 8487 8204
rect 9339 7930 9351 8204
rect 9783 8170 9795 8204
rect 9784 8156 9802 8170
rect 8571 7882 8583 7892
rect 8667 7882 8679 7916
rect 9771 7882 9783 8156
rect 10719 8098 10731 8204
rect 11487 8170 11499 8204
rect 12519 8194 12531 8204
rect 12520 8180 12538 8194
rect 11488 8156 11506 8170
rect 10720 8084 10738 8098
rect 9819 7882 9831 8084
rect 10707 7882 10719 8084
rect 11043 7882 11055 8084
rect 11475 7882 11487 8156
rect 12027 7882 12039 8156
rect 12507 7882 12519 8180
rect 12831 8026 12843 8204
rect 14415 8050 14427 8204
rect 15375 8050 15387 8204
rect 15399 8098 15411 8204
rect 16251 8146 16263 8204
rect 17103 8170 17115 8204
rect 18783 8098 18795 8204
rect 18807 8122 18819 8204
rect 20223 8146 20235 8204
rect 20224 8132 20242 8146
rect 14416 8036 14434 8050
rect 12963 7882 12975 7916
rect 13011 7882 13023 7988
rect 13059 7882 13071 8012
rect 13707 7882 13719 8036
rect 14403 7882 14415 8036
rect 15411 7882 15423 8036
rect 16179 7882 16191 8036
rect 17019 7882 17031 7940
rect 18219 7882 18231 7988
rect 19419 7882 19431 7940
rect 19851 7882 19863 7916
rect 20211 7882 20223 8132
rect 20511 7978 20523 8204
rect 21363 8050 21375 8204
rect 22215 8074 22227 8204
rect 22491 7882 22503 8108
rect 23895 8074 23907 8204
rect 23787 7882 23799 8036
rect 23919 8026 23931 8204
rect 24123 7882 24135 8084
rect 24267 7882 24279 8012
rect 24723 7882 24735 8060
rect 24771 7930 24783 8204
rect 25623 8026 25635 8204
rect 27207 8026 27219 8204
rect 27208 8012 27226 8026
rect 27195 7882 27207 8012
rect 27243 7882 27255 8012
rect 27267 7978 27279 8012
rect 27315 7954 27327 8036
rect 27267 7906 27279 7916
rect 27291 7906 27303 7940
rect 27387 7882 27587 8204
rect 27665 7989 27735 8001
rect 27665 7965 27735 7977
rect 27665 7941 27735 7953
rect 27665 7917 27735 7929
rect 27665 7893 27735 7905
rect 0 3988 70 4000
rect 0 3964 70 3976
rect 123 1577 323 7083
rect 339 1577 351 7083
rect 363 1577 375 7083
rect 387 1577 399 7083
rect 411 1577 423 7083
rect 1611 4025 1623 7083
rect 1659 4049 1671 7083
rect 1731 3953 1743 7083
rect 1779 3929 1791 7083
rect 1827 4073 1839 7083
rect 1851 4097 1863 7083
rect 1899 4121 1911 7083
rect 1947 4145 1959 7083
rect 1995 4169 2007 7083
rect 2067 4193 2079 7083
rect 2115 4217 2127 7083
rect 2187 4241 2199 7083
rect 2235 4289 2247 7083
rect 2043 1577 2055 3891
rect 2091 1577 2103 3867
rect 2235 1577 2247 4251
rect 2307 3881 2319 7083
rect 2331 4313 2343 7083
rect 2283 1577 2295 3843
rect 2307 1577 2319 3819
rect 2355 3809 2367 7083
rect 2355 1577 2367 3771
rect 2403 3761 2415 7083
rect 2427 4337 2439 7083
rect 2403 1577 2415 3723
rect 2427 1577 2439 3699
rect 2451 3689 2463 7083
rect 2499 4361 2511 7083
rect 2523 4385 2535 7083
rect 2547 4409 2559 7083
rect 2571 4433 2583 7083
rect 2643 4481 2655 7083
rect 2667 4505 2679 7083
rect 2451 1577 2463 3651
rect 2499 1577 2511 4035
rect 2523 1577 2535 3627
rect 2595 1577 2607 4443
rect 2691 4145 2703 7083
rect 2739 4529 2751 7083
rect 2619 1577 2631 3603
rect 2643 1577 2655 3579
rect 2667 1577 2679 3555
rect 2715 1577 2727 3531
rect 2739 1577 2751 3507
rect 2763 3497 2775 7083
rect 2811 4553 2823 7083
rect 2859 4577 2871 7083
rect 2907 4625 2919 7083
rect 2979 4649 2991 7083
rect 3003 4673 3015 7083
rect 3027 4697 3039 7083
rect 2787 1577 2799 3939
rect 2835 1577 2847 3939
rect 2859 1577 2871 3699
rect 2883 1577 2895 4587
rect 3003 1577 3015 3459
rect 3051 3449 3063 7083
rect 3075 3425 3087 7083
rect 3123 4721 3135 7083
rect 3147 3401 3159 7083
rect 3171 4745 3183 7083
rect 3219 4769 3231 7083
rect 3243 4793 3255 7083
rect 3267 4817 3279 7083
rect 3291 4841 3303 7083
rect 3315 3377 3327 7083
rect 3363 3353 3375 7083
rect 3387 4865 3399 7083
rect 3411 4889 3423 7083
rect 3459 4913 3471 7083
rect 3483 4937 3495 7083
rect 3363 1577 3375 3315
rect 3411 1577 3423 3291
rect 3507 3281 3519 7083
rect 3555 4961 3567 7083
rect 3579 4985 3591 7083
rect 3603 3401 3615 7083
rect 3651 5009 3663 7083
rect 3675 3881 3687 7083
rect 3699 5033 3711 7083
rect 3747 4121 3759 7083
rect 3771 4841 3783 7083
rect 3555 1577 3567 3387
rect 3603 1577 3615 3243
rect 3627 1577 3639 3219
rect 3747 1577 3759 3195
rect 3771 1577 3783 3171
rect 3795 3161 3807 7083
rect 3843 5057 3855 7083
rect 3867 5081 3879 7083
rect 3843 1577 3855 3123
rect 3867 1577 3879 3099
rect 3891 3089 3903 7083
rect 3915 5105 3927 7083
rect 3939 5129 3951 7083
rect 3987 4145 3999 7083
rect 4011 5153 4023 7083
rect 4035 5177 4047 7083
rect 4059 4145 4071 7083
rect 4107 4145 4119 7083
rect 4131 5201 4143 7083
rect 4155 5225 4167 7083
rect 4203 5249 4215 7083
rect 4227 5273 4239 7083
rect 4251 5297 4263 7083
rect 4275 5321 4287 7083
rect 4299 5345 4311 7083
rect 4347 5369 4359 7083
rect 4371 5417 4383 7083
rect 3915 1577 3927 3051
rect 3939 1577 3951 3027
rect 4011 1577 4023 3003
rect 4035 1577 4047 4131
rect 4107 1577 4119 2979
rect 4131 1577 4143 2955
rect 4203 1577 4215 2931
rect 4227 1577 4239 2907
rect 4275 1577 4287 3939
rect 4371 1577 4383 5379
rect 4395 2897 4407 7083
rect 4443 5441 4455 7083
rect 4467 3785 4479 7083
rect 4491 5489 4503 7083
rect 4419 1577 4431 2859
rect 4443 1577 4455 2835
rect 4491 1577 4503 5451
rect 4515 4433 4527 7083
rect 4563 2825 4575 7083
rect 4587 5009 4599 7083
rect 4611 5513 4623 7083
rect 4659 5561 4671 7083
rect 4587 1577 4599 4491
rect 4659 1577 4671 5523
rect 4683 4505 4695 7083
rect 4707 5585 4719 7083
rect 4755 5609 4767 7083
rect 4779 3065 4791 7083
rect 4803 5633 4815 7083
rect 4851 5657 4863 7083
rect 4683 1577 4695 2787
rect 4779 1577 4791 2763
rect 4803 1577 4815 3891
rect 4875 2921 4887 7083
rect 4923 5681 4935 7083
rect 4875 1577 4887 2739
rect 4923 1577 4935 2715
rect 4971 2705 4983 7083
rect 4995 5705 5007 7083
rect 5019 5729 5031 7083
rect 4995 1577 5007 2667
rect 5043 1577 5055 5739
rect 5067 3617 5079 7083
rect 5091 5777 5103 7083
rect 5091 1577 5103 5187
rect 5139 1577 5151 2643
rect 5163 2633 5175 7083
rect 5187 5801 5199 7083
rect 5211 5825 5223 7083
rect 5259 5849 5271 7083
rect 5283 4601 5295 7083
rect 5307 5873 5319 7083
rect 5355 5897 5367 7083
rect 5211 1577 5223 2595
rect 5307 1577 5319 2571
rect 5331 1577 5343 4587
rect 5355 1577 5367 5163
rect 5379 1577 5391 5883
rect 5403 2561 5415 7083
rect 5427 1577 5439 5019
rect 5451 3521 5463 7083
rect 5475 3785 5487 7083
rect 5499 3737 5511 7083
rect 5523 5105 5535 7083
rect 5571 5105 5583 7083
rect 5595 3641 5607 7083
rect 5643 5921 5655 7083
rect 5475 1577 5487 2667
rect 5571 1577 5583 2523
rect 5595 1577 5607 2499
rect 5691 2489 5703 7083
rect 5715 1577 5727 5931
rect 5763 4409 5775 7083
rect 5811 3041 5823 7083
rect 5835 4409 5847 7083
rect 5883 3041 5895 7083
rect 5931 5969 5943 7083
rect 5955 3737 5967 7083
rect 5979 5993 5991 7083
rect 6027 6017 6039 7083
rect 6051 3713 6063 7083
rect 6075 4649 6087 7083
rect 6123 6041 6135 7083
rect 6075 1577 6087 2451
rect 6123 1577 6135 4635
rect 6147 4625 6159 7083
rect 6171 6065 6183 7083
rect 6219 6089 6231 7083
rect 6267 2777 6279 7083
rect 6291 1577 6303 2427
rect 6315 1577 6327 6099
rect 6339 3905 6351 7083
rect 6363 6041 6375 7083
rect 6411 3521 6423 7083
rect 6459 6137 6471 7083
rect 6483 5633 6495 7083
rect 6363 1577 6375 2403
rect 6387 1577 6399 3507
rect 6459 1577 6471 4899
rect 6507 4553 6519 7083
rect 6531 5633 6543 7083
rect 6483 1577 6495 4011
rect 6555 2993 6567 7083
rect 6603 5729 6615 7083
rect 6627 4505 6639 7083
rect 6651 5153 6663 7083
rect 6699 5153 6711 7083
rect 6507 1577 6519 2379
rect 6555 1577 6567 2955
rect 6579 1577 6591 4467
rect 6675 1577 6687 2979
rect 6699 1577 6711 4539
rect 6723 2753 6735 7083
rect 6747 5729 6759 7083
rect 6795 6041 6807 7083
rect 6819 3977 6831 7083
rect 6843 6161 6855 7083
rect 6867 6185 6879 7083
rect 6915 6209 6927 7083
rect 6939 6233 6951 7083
rect 6723 1577 6735 2427
rect 6747 1577 6759 3963
rect 6795 1577 6807 2907
rect 6819 1577 6831 3627
rect 6867 1577 6879 2355
rect 6915 1577 6927 3219
rect 6939 1577 6951 3123
rect 6963 2345 6975 7083
rect 7011 5849 7023 7083
rect 7059 6257 7071 7083
rect 7131 4649 7143 7083
rect 7155 6281 7167 7083
rect 7179 6305 7191 7083
rect 7227 6353 7239 7083
rect 6987 1577 6999 2307
rect 7059 1577 7071 3867
rect 7155 1577 7167 2283
rect 7179 1577 7191 2259
rect 7227 1577 7239 6315
rect 7251 6257 7263 7083
rect 7275 4049 7287 7083
rect 7299 5297 7311 7083
rect 7347 5297 7359 7083
rect 7371 5993 7383 7083
rect 7395 4097 7407 7083
rect 7419 4241 7431 7083
rect 7251 1577 7263 2235
rect 7275 1577 7287 2211
rect 7371 1577 7383 3867
rect 7395 1577 7407 3771
rect 7443 2201 7455 6027
rect 7467 2921 7479 7083
rect 7491 5993 7503 7083
rect 7419 1577 7431 2187
rect 7491 1577 7503 4227
rect 7515 2201 7527 7083
rect 7563 2177 7575 7083
rect 7587 6377 7599 7083
rect 7611 6401 7623 7083
rect 7635 4841 7647 7083
rect 7707 6473 7719 7083
rect 7731 6497 7743 7083
rect 7611 1577 7623 3243
rect 7635 1577 7647 2907
rect 7659 1577 7671 6411
rect 7707 1577 7719 6435
rect 7731 1577 7743 3051
rect 7755 2153 7767 7083
rect 7779 6521 7791 7083
rect 7803 5537 7815 7083
rect 7851 4913 7863 7083
rect 7875 5537 7887 7083
rect 7899 6521 7911 7083
rect 7779 1577 7791 4467
rect 7827 1577 7839 2907
rect 7851 1577 7863 2115
rect 7923 1577 7935 5955
rect 7947 3593 7959 7083
rect 7971 4769 7983 7083
rect 7995 6521 8007 7083
rect 8019 6545 8031 7083
rect 8007 2129 8019 5091
rect 8031 2105 8043 5427
rect 7947 1577 7959 2091
rect 7971 1577 7983 2067
rect 8019 1577 8031 2043
rect 8067 1577 8079 3747
rect 8091 2129 8103 7083
rect 8115 3761 8127 7083
rect 8163 4721 8175 7083
rect 8139 1577 8151 3291
rect 8187 2105 8199 5643
rect 8211 4193 8223 7083
rect 8235 4025 8247 7083
rect 8259 6569 8271 7083
rect 8307 6593 8319 7083
rect 8331 6617 8343 7083
rect 8355 6641 8367 7083
rect 8379 6665 8391 7083
rect 8403 6689 8415 7083
rect 8163 1577 8175 2091
rect 8211 1577 8223 3843
rect 8259 1577 8271 3747
rect 8283 1577 8295 2091
rect 8307 1577 8319 2019
rect 8355 1577 8367 1995
rect 8379 1577 8391 1971
rect 8403 1577 8415 6579
rect 8451 5393 8463 7083
rect 8475 5993 8487 7083
rect 8499 5393 8511 7083
rect 8547 6593 8559 7083
rect 8451 1577 8463 3315
rect 8571 1577 8583 1947
rect 8595 1937 8607 7083
rect 8619 1577 8631 6339
rect 8643 4145 8655 7083
rect 8667 4313 8679 7083
rect 8715 6713 8727 7083
rect 8691 1577 8703 3819
rect 8739 1577 8751 2595
rect 8763 1913 8775 7083
rect 8787 4913 8799 7083
rect 8787 1577 8799 4299
rect 8811 2009 8823 7083
rect 8859 3305 8871 7083
rect 8883 3113 8895 7083
rect 8907 6737 8919 7083
rect 8835 1577 8847 2907
rect 8907 1577 8919 5715
rect 8931 5657 8943 7083
rect 8955 4841 8967 7083
rect 9003 5729 9015 7083
rect 9027 5273 9039 7083
rect 9051 5585 9063 7083
rect 8979 2009 8991 5259
rect 8931 1577 8943 1971
rect 8955 1577 8967 1995
rect 9027 1577 9039 4995
rect 9051 1577 9063 5235
rect 9075 2009 9087 7083
rect 9099 5249 9111 7083
rect 9099 1577 9111 5139
rect 9147 4625 9159 7083
rect 9171 2681 9183 7083
rect 9195 3977 9207 7083
rect 9219 5585 9231 7083
rect 9243 6761 9255 7083
rect 9291 6737 9303 7083
rect 9315 6785 9327 7083
rect 9339 6809 9351 7083
rect 9147 1577 9159 1875
rect 9219 1577 9231 4899
rect 9243 1577 9255 3699
rect 9267 1577 9279 6075
rect 9315 1577 9327 3819
rect 9339 1577 9351 4851
rect 9387 4841 9399 7083
rect 9411 4121 9423 7083
rect 9435 2033 9447 7083
rect 9459 4121 9471 7083
rect 9507 6377 9519 7083
rect 9531 4289 9543 7083
rect 9555 4361 9567 7083
rect 9579 6833 9591 7083
rect 9363 1577 9375 1899
rect 9459 1577 9471 2379
rect 9483 1577 9495 3915
rect 9531 1577 9543 3915
rect 9555 1577 9567 1899
rect 9579 1577 9591 4467
rect 9603 4289 9615 7083
rect 9651 6857 9663 7083
rect 9627 3065 9639 5571
rect 9651 1577 9663 5355
rect 9675 3113 9687 7083
rect 9699 2537 9711 6747
rect 9723 2945 9735 7083
rect 9771 5585 9783 7083
rect 9675 1577 9687 1851
rect 9747 1577 9759 3411
rect 9795 3329 9807 6771
rect 9819 3137 9831 7083
rect 9867 6761 9879 7083
rect 9843 3929 9855 6147
rect 9771 1577 9783 2523
rect 9819 1577 9831 1827
rect 9867 1577 9879 4899
rect 9891 1577 9903 3291
rect 9915 2585 9927 6843
rect 9939 6785 9951 7083
rect 9963 6857 9975 7083
rect 9963 1577 9975 5883
rect 9987 4745 9999 7083
rect 10011 5945 10023 7083
rect 9987 1577 9999 3915
rect 10035 1865 10047 5979
rect 10059 3977 10071 7083
rect 10083 5009 10095 7083
rect 10059 1577 10071 3411
rect 10083 1577 10095 2883
rect 10107 1577 10119 2475
rect 10131 1913 10143 7083
rect 10179 2921 10191 7083
rect 10203 4049 10215 7083
rect 10227 5177 10239 7083
rect 10275 4745 10287 7083
rect 10299 6041 10311 7083
rect 10323 5945 10335 7083
rect 10347 4049 10359 6147
rect 10371 5561 10383 7083
rect 10155 1577 10167 2427
rect 10299 1577 10311 4035
rect 10323 1577 10335 2883
rect 10395 1577 10407 5955
rect 10419 4049 10431 7083
rect 10491 5129 10503 7083
rect 10539 6881 10551 7083
rect 10419 1577 10431 3627
rect 10443 1577 10455 2475
rect 10467 2129 10479 4035
rect 10491 1577 10503 1851
rect 10539 1577 10551 5427
rect 10611 5129 10623 7083
rect 10635 4049 10647 7083
rect 10659 6329 10671 7083
rect 10707 5129 10719 7083
rect 10611 1577 10623 3987
rect 10671 1985 10683 5115
rect 10755 3857 10767 7083
rect 10779 6737 10791 7083
rect 10731 1577 10743 2403
rect 10755 1577 10767 3843
rect 10827 2585 10839 7083
rect 10827 1577 10839 1803
rect 10851 1577 10863 6315
rect 10875 5801 10887 7083
rect 10923 5969 10935 7083
rect 10995 6905 11007 7083
rect 11115 6905 11127 7083
rect 10899 1577 10911 4995
rect 10947 1817 10959 6075
rect 10923 1577 10935 1779
rect 10971 1577 10983 2715
rect 10995 1577 11007 3699
rect 11031 3593 11043 6891
rect 11019 1577 11031 1803
rect 11091 1577 11103 6723
rect 11139 5009 11151 7083
rect 11115 1577 11127 3579
rect 11163 2441 11175 6891
rect 11163 1577 11175 1755
rect 11187 1745 11199 7083
rect 11211 1577 11223 6579
rect 11235 3833 11247 7083
rect 11259 5657 11271 7083
rect 11307 3017 11319 7083
rect 11355 6905 11367 7083
rect 11235 1577 11247 1707
rect 11307 1577 11319 1683
rect 11331 1577 11343 5979
rect 11379 4841 11391 7083
rect 11427 4361 11439 7083
rect 11475 6929 11487 7083
rect 11355 1577 11367 4011
rect 11403 1577 11415 3699
rect 11427 1577 11439 1659
rect 11451 1577 11463 5187
rect 11475 1673 11487 5091
rect 11499 1577 11511 6939
rect 11523 4913 11535 7083
rect 11547 2897 11559 7083
rect 11571 6977 11583 7083
rect 11571 1577 11583 6315
rect 11619 3857 11631 7083
rect 11595 1577 11607 2883
rect 11643 1889 11655 7083
rect 11667 7001 11679 7083
rect 11667 1577 11679 5163
rect 11691 4457 11703 7083
rect 11715 2681 11727 6987
rect 11739 4457 11751 7083
rect 11763 7001 11775 7083
rect 11787 7025 11799 7083
rect 11763 1577 11775 6003
rect 11787 1577 11799 5475
rect 11811 2801 11823 7011
rect 11835 1913 11847 7083
rect 11859 4169 11871 7083
rect 11883 2993 11895 7083
rect 11931 4721 11943 7083
rect 11835 1577 11847 1875
rect 11955 1769 11967 7083
rect 11979 7025 11991 7083
rect 12027 1889 12039 7083
rect 12075 2945 12087 7083
rect 12099 5537 12111 7083
rect 12147 4145 12159 7083
rect 12195 4721 12207 7083
rect 12219 4145 12231 7083
rect 12243 2993 12255 7083
rect 12291 4049 12303 7083
rect 12315 6737 12327 7083
rect 12339 2801 12351 7083
rect 12387 3017 12399 7083
rect 12411 1889 12423 7083
rect 12459 1769 12471 7083
rect 12507 2513 12519 7083
rect 12555 2513 12567 7083
rect 12579 3977 12591 7083
rect 12603 5297 12615 7083
rect 12651 5297 12663 7083
rect 12675 6185 12687 7083
rect 12723 6377 12735 7083
rect 12771 5969 12783 7083
rect 12459 1577 12471 1659
rect 12603 1577 12615 4131
rect 12651 1577 12663 4131
rect 12675 1577 12687 1947
rect 12699 1577 12711 5139
rect 12747 1577 12759 3675
rect 12771 1577 12783 5139
rect 12795 4169 12807 7083
rect 12819 6905 12831 7083
rect 12867 6425 12879 7083
rect 12891 6185 12903 7083
rect 12915 6377 12927 7083
rect 12819 1577 12831 3675
rect 12867 1577 12879 3723
rect 12891 1577 12903 1875
rect 12915 1577 12927 4563
rect 12963 3689 12975 7083
rect 13131 6425 13143 7083
rect 12963 1577 12975 3051
rect 13011 1577 13023 1947
rect 13083 1577 13095 2931
rect 13107 1577 13119 4923
rect 13155 3857 13167 7083
rect 13203 3977 13215 7083
rect 13155 1577 13167 3675
rect 13203 1577 13215 1635
rect 13227 1577 13239 4491
rect 13251 1889 13263 7083
rect 13275 3833 13287 7083
rect 13299 6905 13311 7083
rect 13323 7049 13335 7083
rect 13371 6257 13383 7083
rect 13299 1577 13311 2643
rect 13323 1577 13335 2931
rect 13347 1577 13359 5979
rect 13371 1577 13383 4779
rect 13395 4169 13407 7083
rect 13419 4073 13431 7083
rect 13467 7073 13479 7083
rect 13419 1577 13431 1611
rect 13443 1577 13455 1683
rect 13467 1577 13479 5067
rect 13491 2729 13503 7083
rect 13515 1577 13527 4779
rect 13539 2057 13551 7083
rect 13587 5969 13599 7083
rect 13611 4625 13623 7083
rect 13539 1577 13551 1587
rect 13563 1577 13575 4155
rect 13611 1577 13623 4059
rect 13635 1649 13647 6411
rect 13659 4793 13671 7083
rect 13659 1577 13671 3771
rect 13683 1577 13695 5427
rect 13707 3233 13719 7083
rect 13731 5081 13743 7083
rect 13755 3137 13767 7083
rect 13779 5633 13791 7083
rect 13803 1961 13815 6891
rect 13827 2945 13839 7083
rect 13851 5705 13863 7083
rect 13875 5801 13887 7083
rect 13923 5801 13935 7083
rect 13755 1577 13767 1755
rect 13875 1577 13887 2307
rect 13899 1577 13911 3747
rect 13923 1577 13935 5691
rect 13947 5633 13959 7083
rect 13947 1577 13959 5283
rect 13971 1625 13983 6699
rect 13995 4865 14007 7083
rect 13995 1577 14007 4779
rect 14043 2273 14055 7083
rect 14067 3329 14079 7083
rect 14091 4145 14103 7059
rect 14115 4793 14127 7083
rect 14163 6425 14175 7083
rect 14019 1577 14031 1731
rect 14067 1577 14079 2715
rect 14115 1577 14127 2835
rect 14139 1577 14151 2859
rect 14187 2321 14199 7083
rect 14211 4073 14223 6579
rect 14235 5297 14247 7083
rect 14283 6593 14295 7083
rect 14235 1577 14247 5187
rect 14259 1577 14271 5979
rect 14283 1577 14295 4923
rect 14307 1673 14319 5787
rect 14331 4937 14343 7083
rect 14331 1577 14343 3819
rect 14367 2729 14379 6387
rect 14403 5201 14415 7083
rect 14451 5801 14463 7083
rect 14475 6401 14487 7083
rect 14355 1577 14367 2355
rect 14427 2105 14439 5283
rect 14451 1577 14463 5523
rect 14475 1577 14487 5811
rect 14499 5297 14511 7083
rect 14523 5825 14535 7083
rect 14571 5345 14583 7083
rect 14619 5297 14631 7083
rect 14499 1577 14511 5091
rect 14523 1577 14535 3075
rect 14547 2993 14559 5283
rect 14571 1577 14583 2667
rect 14595 1577 14607 3315
rect 14643 1577 14655 4323
rect 14691 2609 14703 7083
rect 14715 6041 14727 7083
rect 14739 6905 14751 7083
rect 14691 1577 14703 2259
rect 14739 1577 14751 6723
rect 14811 1577 14823 2571
rect 14835 1577 14847 6147
rect 14859 5345 14871 7083
rect 15219 6281 15231 7083
rect 14883 1577 14895 3747
rect 14979 1577 14991 4059
rect 15099 1577 15111 4731
rect 15195 1577 15207 3747
rect 15219 1577 15231 3075
rect 15243 1577 15255 5043
rect 15267 3929 15279 7083
rect 15315 1577 15327 4347
rect 15339 1577 15351 4371
rect 15411 3569 15423 7083
rect 15387 1577 15399 2979
rect 15435 1577 15447 3867
rect 15459 3833 15471 7083
rect 15483 4625 15495 7083
rect 15459 1577 15471 3555
rect 15507 2753 15519 7083
rect 15627 6689 15639 7083
rect 15531 3569 15543 5643
rect 15483 1577 15495 2715
rect 15555 1577 15567 2739
rect 15579 1577 15591 2403
rect 15627 1577 15639 3555
rect 15651 1577 15663 1755
rect 15747 1577 15759 5667
rect 15771 1577 15783 3699
rect 15867 1577 15879 3243
rect 15891 1577 15903 3123
rect 15963 1577 15975 5019
rect 15987 3833 15999 7083
rect 15987 1577 15999 3795
rect 16035 3113 16047 7083
rect 16011 1577 16023 1731
rect 16107 1577 16119 3795
rect 16131 1577 16143 5331
rect 16179 2993 16191 7083
rect 16227 3521 16239 7083
rect 16251 4505 16263 7083
rect 16275 5057 16287 7083
rect 16179 1577 16191 2091
rect 16203 1577 16215 3051
rect 16227 1577 16239 2979
rect 16275 1577 16287 4755
rect 16299 2993 16311 5547
rect 16323 5009 16335 7083
rect 16347 5681 16359 7083
rect 16371 5465 16383 7083
rect 16395 3569 16407 7083
rect 16443 6761 16455 7083
rect 16323 1577 16335 1659
rect 16395 1577 16407 2835
rect 16419 1577 16431 1947
rect 16443 1577 16455 3483
rect 16467 3233 16479 7083
rect 16491 1673 16503 5355
rect 16515 5345 16527 7083
rect 16515 1577 16527 4995
rect 16539 1577 16551 6459
rect 16563 3833 16575 7083
rect 16587 3641 16599 7083
rect 16587 1577 16599 3555
rect 16611 1577 16623 3867
rect 16635 3257 16647 7083
rect 16683 5705 16695 7083
rect 16707 3881 16719 7083
rect 16731 3641 16743 7083
rect 16755 5465 16767 7083
rect 16767 4409 16779 5331
rect 16659 1577 16671 3483
rect 16707 1577 16719 3243
rect 16803 3233 16815 7083
rect 16827 3137 16839 7083
rect 16851 6449 16863 7083
rect 16863 3257 16875 6075
rect 16731 1577 16743 2979
rect 16899 2657 16911 7083
rect 16923 5537 16935 7083
rect 16947 6233 16959 7083
rect 16971 3569 16983 7035
rect 16995 5873 17007 7083
rect 17019 3089 17031 7083
rect 17043 4673 17055 7083
rect 17067 2993 17079 6963
rect 17091 4673 17103 7083
rect 17115 2921 17127 7083
rect 17139 4457 17151 7083
rect 17187 5369 17199 7083
rect 17211 6569 17223 7083
rect 17235 3209 17247 7083
rect 17283 5249 17295 7083
rect 17307 1577 17319 5619
rect 17331 4601 17343 7083
rect 17403 5441 17415 7083
rect 17427 1913 17439 7083
rect 17451 5249 17463 7083
rect 17475 5777 17487 7083
rect 17523 6449 17535 7083
rect 17451 1577 17463 4971
rect 17475 1577 17487 3555
rect 17499 1577 17511 4875
rect 17523 1577 17535 6315
rect 17547 3329 17559 7083
rect 17571 5321 17583 7083
rect 17547 1577 17559 2811
rect 17595 1577 17607 6723
rect 17619 6473 17631 7083
rect 17619 1577 17631 6315
rect 17643 5225 17655 7083
rect 17691 4169 17703 7083
rect 17667 1577 17679 3099
rect 17715 3065 17727 5235
rect 17739 1577 17751 5163
rect 17763 3569 17775 6603
rect 17811 4457 17823 7083
rect 17787 1577 17799 3723
rect 17907 1577 17919 6915
rect 17979 1577 17991 4155
rect 18003 1577 18015 5091
rect 18051 1577 18063 3555
rect 18099 1577 18111 3075
rect 18147 1577 18159 5091
rect 18219 1577 18231 2355
rect 18243 1577 18255 5403
rect 18267 1577 18279 1995
rect 18315 1577 18327 3627
rect 18363 2945 18375 7083
rect 18387 2369 18399 7083
rect 18411 4769 18423 7083
rect 18363 1577 18375 1875
rect 18435 1577 18447 3867
rect 18459 3113 18471 7083
rect 18483 4601 18495 7083
rect 18507 6161 18519 7083
rect 18531 5177 18543 7083
rect 18579 5657 18591 7083
rect 18603 3329 18615 7083
rect 18699 6689 18711 7083
rect 18459 1577 18471 2979
rect 18483 1577 18495 3315
rect 18555 1577 18567 3123
rect 18579 1577 18591 3051
rect 18627 2777 18639 4587
rect 18651 1577 18663 3003
rect 18675 1577 18687 3291
rect 18699 1577 18711 6651
rect 18723 6329 18735 6675
rect 18771 3833 18783 7083
rect 18795 5657 18807 7083
rect 18819 6185 18831 7083
rect 18747 1577 18759 3243
rect 18831 3209 18843 5667
rect 18867 4601 18879 7083
rect 18891 4625 18903 7083
rect 18939 5225 18951 7083
rect 18771 1577 18783 3195
rect 18819 1577 18831 3123
rect 18867 1577 18879 2931
rect 18891 1577 18903 3195
rect 18915 1577 18927 3435
rect 18963 1577 18975 6579
rect 18987 2057 18999 7083
rect 19011 6185 19023 7083
rect 19035 5249 19047 7083
rect 19083 6257 19095 7083
rect 19107 6353 19119 7083
rect 19131 4169 19143 7083
rect 19179 6041 19191 7083
rect 19203 4601 19215 7083
rect 18987 1577 18999 1995
rect 19011 1577 19023 3435
rect 19059 1577 19071 2835
rect 19083 1577 19095 3051
rect 19155 2585 19167 4587
rect 19227 3713 19239 7083
rect 19251 2297 19263 7083
rect 19275 3209 19287 5403
rect 19251 1577 19263 2043
rect 19299 1601 19311 7083
rect 19323 3089 19335 7083
rect 19347 3449 19359 6387
rect 19371 2537 19383 7083
rect 19419 2009 19431 7083
rect 19467 2393 19479 7083
rect 19515 4745 19527 7083
rect 19587 1841 19599 7083
rect 19611 4745 19623 7083
rect 19659 4817 19671 7083
rect 19707 4793 19719 7083
rect 19731 6449 19743 7083
rect 19779 4553 19791 7083
rect 19827 5897 19839 7083
rect 19851 4649 19863 7083
rect 19875 6785 19887 7083
rect 19803 1577 19815 2331
rect 19827 1577 19839 4299
rect 19851 1577 19863 4155
rect 19899 1577 19911 5667
rect 19923 5249 19935 7083
rect 19923 1577 19935 5091
rect 19947 3329 19959 7083
rect 19971 4553 19983 7083
rect 20019 3833 20031 7083
rect 20043 3737 20055 7083
rect 19995 1577 20007 3435
rect 20019 1577 20031 3195
rect 20067 2753 20079 7083
rect 20091 1577 20103 6363
rect 20115 2417 20127 7083
rect 20139 3329 20151 7083
rect 20163 4649 20175 7083
rect 20187 4169 20199 5715
rect 20211 3185 20223 7083
rect 20211 1577 20223 3003
rect 20235 1577 20247 5691
rect 20259 4793 20271 7083
rect 20283 5177 20295 7083
rect 20331 6617 20343 7083
rect 20259 1577 20271 4179
rect 20307 1577 20319 4179
rect 20331 1577 20343 4827
rect 20355 3209 20367 4755
rect 20379 4265 20391 7083
rect 20427 6929 20439 7083
rect 20403 3017 20415 5979
rect 20427 1577 20439 6891
rect 20451 2225 20463 4779
rect 20475 2057 20487 6915
rect 20499 6305 20511 7083
rect 20523 6569 20535 7083
rect 20499 1577 20511 5211
rect 20523 1577 20535 6411
rect 20547 4769 20559 7083
rect 20595 3953 20607 7083
rect 20619 4793 20631 7083
rect 20619 1577 20631 3579
rect 20643 1577 20655 5187
rect 20667 3761 20679 7083
rect 20691 1577 20703 5691
rect 20715 4217 20727 7083
rect 20739 3113 20751 7083
rect 20763 5681 20775 7083
rect 20787 5921 20799 7083
rect 20811 4817 20823 7083
rect 20715 1577 20727 3051
rect 20739 1577 20751 3003
rect 20787 1577 20799 1755
rect 20811 1577 20823 2379
rect 20835 1577 20847 3339
rect 20859 1817 20871 7083
rect 20883 6185 20895 7083
rect 20883 1577 20895 5691
rect 20907 2993 20919 7083
rect 20955 4841 20967 7083
rect 20931 1577 20943 3699
rect 20979 3113 20991 7083
rect 21003 6641 21015 7083
rect 21051 4889 21063 7083
rect 21075 6737 21087 7083
rect 21099 4841 21111 7083
rect 21147 5177 21159 7083
rect 21003 1577 21015 4491
rect 21027 1577 21039 2907
rect 21051 1577 21063 1851
rect 21123 1577 21135 4851
rect 21147 1577 21159 4947
rect 21171 2321 21183 7083
rect 21195 4529 21207 7083
rect 21243 6113 21255 7083
rect 21267 6041 21279 7083
rect 21195 1577 21207 4395
rect 21291 3425 21303 7083
rect 21339 6089 21351 7083
rect 21219 1577 21231 2931
rect 21243 1577 21255 1947
rect 21267 1577 21279 2619
rect 21315 1577 21327 4491
rect 21339 1577 21351 5955
rect 21387 2969 21399 7083
rect 21531 6617 21543 7083
rect 21411 2657 21423 4779
rect 21495 4769 21507 5163
rect 21363 1577 21375 2307
rect 21435 1577 21447 2787
rect 21459 1577 21471 3291
rect 21483 1577 21495 4251
rect 21531 1577 21543 6531
rect 21567 5825 21579 6603
rect 21555 1577 21567 4563
rect 21579 3017 21591 5475
rect 21603 1577 21615 6003
rect 21627 2225 21639 4803
rect 21651 1577 21663 5211
rect 21675 1577 21687 5691
rect 21699 1577 21711 6819
rect 21747 1577 21759 4371
rect 21771 1577 21783 6867
rect 21795 1577 21807 6819
rect 21819 1577 21831 5115
rect 21939 5081 21951 7083
rect 21867 1577 21879 4155
rect 21891 1577 21903 2187
rect 21987 1577 21999 3579
rect 22059 1577 22071 5235
rect 22083 4529 22095 7083
rect 22083 1577 22095 4323
rect 22107 4025 22119 7083
rect 22131 6473 22143 7083
rect 22179 6569 22191 7083
rect 22203 6305 22215 7083
rect 22143 3953 22155 4515
rect 22227 4409 22239 7083
rect 22251 6137 22263 7083
rect 22263 3953 22275 4587
rect 22299 4409 22311 7083
rect 22179 1577 22191 2739
rect 22227 1577 22239 3939
rect 22299 1577 22311 3939
rect 22347 2873 22359 7083
rect 22419 6089 22431 7083
rect 22443 6353 22455 7083
rect 22347 1577 22359 2139
rect 22419 1577 22431 4323
rect 22443 1577 22455 4035
rect 22491 1577 22503 5571
rect 22539 4049 22551 7083
rect 22563 4337 22575 7083
rect 22539 1577 22551 2931
rect 22563 1577 22575 3723
rect 22587 2441 22599 7083
rect 22611 3305 22623 4323
rect 22635 4217 22647 7083
rect 22659 5921 22671 7083
rect 22683 6209 22695 7083
rect 22635 1577 22647 2019
rect 22707 1577 22719 4731
rect 22731 2273 22743 7083
rect 22755 4337 22767 7083
rect 22779 6953 22791 7083
rect 22827 6353 22839 7083
rect 22851 6257 22863 7083
rect 22755 1577 22767 3819
rect 22803 1577 22815 5259
rect 22875 4505 22887 7083
rect 22899 4193 22911 7083
rect 22947 4721 22959 7083
rect 22971 6017 22983 7083
rect 22851 1577 22863 1755
rect 22875 1577 22887 3267
rect 22923 3113 22935 4323
rect 22947 1577 22959 3747
rect 22971 1577 22983 5979
rect 22995 3809 23007 7083
rect 23043 6113 23055 7083
rect 23067 6041 23079 7083
rect 23115 6449 23127 7083
rect 23043 1577 23055 6027
rect 23067 1577 23079 3867
rect 23091 1577 23103 3771
rect 23115 1577 23127 4323
rect 23139 4049 23151 6099
rect 23163 5753 23175 7083
rect 23187 5945 23199 7083
rect 23211 6113 23223 7083
rect 23187 1577 23199 4419
rect 23211 1577 23223 6027
rect 23235 2729 23247 7083
rect 23259 3953 23271 7083
rect 23283 5393 23295 6099
rect 23307 4481 23319 7083
rect 23331 4409 23343 7083
rect 23307 1577 23319 4203
rect 23355 4169 23367 7083
rect 23331 1577 23343 3867
rect 23355 1577 23367 3963
rect 23403 3089 23415 7083
rect 23451 5993 23463 7083
rect 23523 6809 23535 7083
rect 23571 5729 23583 7083
rect 23427 4217 23439 5427
rect 23379 1577 23391 1947
rect 23451 1577 23463 4539
rect 23475 1577 23487 4203
rect 23499 1697 23511 4395
rect 23547 1577 23559 3819
rect 23571 1577 23583 5691
rect 23595 1985 23607 5715
rect 23619 1577 23631 6411
rect 23643 4913 23655 7083
rect 23667 3833 23679 7083
rect 23691 4865 23703 7083
rect 23715 4985 23727 7083
rect 23763 6593 23775 7083
rect 23811 6857 23823 7083
rect 23859 5681 23871 7083
rect 23739 1577 23751 2163
rect 23787 1577 23799 4491
rect 23811 1577 23823 4299
rect 23859 1577 23871 4179
rect 23883 1889 23895 7083
rect 23907 1769 23919 7083
rect 23955 6809 23967 7083
rect 23931 4193 23943 6147
rect 23979 4913 23991 7083
rect 24003 2249 24015 7083
rect 24051 4937 24063 7083
rect 24075 5297 24087 7083
rect 24099 4385 24111 7083
rect 23907 1577 23919 1659
rect 24027 1577 24039 4371
rect 24075 1577 24087 1875
rect 24099 1577 24111 2931
rect 24123 1577 24135 5091
rect 24171 3401 24183 7083
rect 24195 6737 24207 7083
rect 24147 1577 24159 1587
rect 24195 1577 24207 5091
rect 24219 4409 24231 7083
rect 24267 3929 24279 7083
rect 24291 2465 24303 7083
rect 24315 6569 24327 7083
rect 24243 1577 24255 1683
rect 24315 1577 24327 4635
rect 24339 1577 24351 6171
rect 24363 4433 24375 7083
rect 24363 1577 24375 3531
rect 24387 2489 24399 7083
rect 24411 1673 24423 6003
rect 24435 4697 24447 7083
rect 24447 2801 24459 4371
rect 24483 1961 24495 7083
rect 24507 4625 24519 7083
rect 24531 1913 24543 7083
rect 24555 4001 24567 7083
rect 24579 4433 24591 7083
rect 24627 4913 24639 7083
rect 24651 3089 24663 7083
rect 24675 4385 24687 7083
rect 24723 5081 24735 7083
rect 24747 2849 24759 7083
rect 24795 5609 24807 7083
rect 24843 5969 24855 7083
rect 24843 1577 24855 5643
rect 24867 4313 24879 7083
rect 24891 5849 24903 7083
rect 24939 5009 24951 7083
rect 24891 1577 24903 4899
rect 24963 3905 24975 7083
rect 24987 2273 24999 7083
rect 25035 2081 25047 7083
rect 25059 4361 25071 7083
rect 25083 6569 25095 7083
rect 25035 1577 25047 2043
rect 25059 1577 25071 4299
rect 25083 1577 25095 6483
rect 25107 4361 25119 7083
rect 25131 1577 25143 5883
rect 25155 1697 25167 7083
rect 25179 5825 25191 7083
rect 25155 1577 25167 1659
rect 25179 1577 25191 5787
rect 25203 2057 25215 6363
rect 25227 5417 25239 7083
rect 25275 5057 25287 7083
rect 25299 6065 25311 7083
rect 25239 4313 25251 4995
rect 25227 1577 25239 2307
rect 25275 1577 25287 2691
rect 25323 2513 25335 7083
rect 25347 4745 25359 6555
rect 25371 3041 25383 7083
rect 25395 1673 25407 5067
rect 25419 3257 25431 7083
rect 25419 1577 25431 3195
rect 25443 3089 25455 5811
rect 25491 3641 25503 7083
rect 25515 3089 25527 7083
rect 25563 5537 25575 7083
rect 25611 4409 25623 7083
rect 25635 4265 25647 7083
rect 25659 3473 25671 7083
rect 25707 6713 25719 7083
rect 25731 2657 25743 7083
rect 25755 6089 25767 7083
rect 25779 1577 25791 6027
rect 25803 3785 25815 7083
rect 25827 5057 25839 7083
rect 25851 6545 25863 7083
rect 25827 1577 25839 4995
rect 25863 2681 25875 5043
rect 25899 1745 25911 7083
rect 25923 3713 25935 7083
rect 25947 7001 25959 7083
rect 25995 5969 26007 7083
rect 25971 1577 25983 2091
rect 25995 1577 26007 4299
rect 26019 1889 26031 7083
rect 26043 4409 26055 7083
rect 26091 6761 26103 7083
rect 26067 4313 26079 6147
rect 26043 1577 26055 4131
rect 26115 3233 26127 7083
rect 26139 4433 26151 7083
rect 26091 1577 26103 2955
rect 26139 1577 26151 3603
rect 26163 3449 26175 4395
rect 26187 4241 26199 7083
rect 26211 5513 26223 7083
rect 26235 5033 26247 7083
rect 26211 1577 26223 3507
rect 26235 1577 26247 4083
rect 26259 3209 26271 7083
rect 26307 4409 26319 7083
rect 26331 6041 26343 7083
rect 26283 1577 26295 2595
rect 26307 1577 26319 3867
rect 26331 1577 26343 4227
rect 26355 4217 26367 7083
rect 26379 2849 26391 4419
rect 26403 3833 26415 7083
rect 26427 4025 26439 7083
rect 26427 1577 26439 3987
rect 26451 3593 26463 7083
rect 26475 3545 26487 4395
rect 26499 3665 26511 7083
rect 26523 4409 26535 7083
rect 26547 7049 26559 7083
rect 26499 1577 26511 2547
rect 26523 1577 26535 1923
rect 26547 1577 26559 7011
rect 26595 5009 26607 7083
rect 26571 1577 26583 4443
rect 26619 3857 26631 7083
rect 26643 2129 26655 7083
rect 26667 6161 26679 7083
rect 26691 5153 26703 7083
rect 26739 5465 26751 7083
rect 26763 4385 26775 7083
rect 26787 4673 26799 7083
rect 26619 1577 26631 1875
rect 26643 1577 26655 1947
rect 26715 1577 26727 4107
rect 26835 3569 26847 7083
rect 26859 3689 26871 7083
rect 26907 6521 26919 7083
rect 26763 1577 26775 3363
rect 26811 1577 26823 3147
rect 26883 1865 26895 4395
rect 26931 4337 26943 7035
rect 26955 3137 26967 7083
rect 26979 3497 26991 7083
rect 27027 4073 27039 7083
rect 27075 6185 27087 7083
rect 27123 4049 27135 7083
rect 27195 4001 27207 7083
rect 27243 1721 27255 7083
rect 27267 1601 27279 4347
rect 27291 1625 27303 1779
rect 27315 1649 27327 4275
rect 27387 1577 27587 7083
rect 27665 2884 27735 2896
rect 27665 1636 27735 1648
rect 27665 1612 27735 1624
rect 27665 1588 27735 1600
rect 0 59 70 71
rect 0 35 70 47
rect 123 0 323 778
rect 339 0 351 778
rect 363 0 375 778
rect 387 0 399 778
rect 411 0 423 778
rect 1683 96 1695 778
rect 2235 48 2247 778
rect 2547 48 2559 778
rect 3555 24 3567 778
rect 3651 120 3663 778
rect 3699 144 3711 778
rect 3723 168 3735 778
rect 4059 192 4071 778
rect 4155 216 4167 778
rect 4323 240 4335 778
rect 4347 264 4359 778
rect 4467 288 4479 778
rect 4539 48 4551 778
rect 4731 312 4743 778
rect 4827 264 4839 778
rect 5019 264 5031 778
rect 5235 336 5247 778
rect 5259 360 5271 778
rect 5547 384 5559 778
rect 6267 408 6279 778
rect 6411 432 6423 778
rect 6603 384 6615 778
rect 6651 456 6663 778
rect 7035 360 7047 778
rect 7083 360 7095 778
rect 7131 432 7143 778
rect 7299 192 7311 778
rect 7323 432 7335 778
rect 7443 192 7455 778
rect 7515 480 7527 778
rect 7563 504 7575 778
rect 7875 528 7887 778
rect 8475 576 8487 778
rect 7983 0 7995 538
rect 8499 336 8511 778
rect 8547 336 8559 778
rect 8667 600 8679 778
rect 9003 624 9015 778
rect 9411 240 9423 778
rect 9435 504 9447 778
rect 9603 504 9615 778
rect 9699 648 9711 778
rect 9915 600 9927 778
rect 10011 600 10023 778
rect 10203 624 10215 778
rect 10275 672 10287 778
rect 10371 696 10383 778
rect 10659 576 10671 778
rect 10779 408 10791 778
rect 10875 408 10887 778
rect 11067 624 11079 778
rect 11163 576 11175 778
rect 11259 576 11271 778
rect 11523 720 11535 778
rect 11176 562 11194 576
rect 11175 0 11187 562
rect 11547 312 11559 778
rect 11643 192 11655 778
rect 11715 312 11727 778
rect 11883 192 11895 778
rect 11931 744 11943 778
rect 12603 552 12615 778
rect 12795 552 12807 778
rect 13251 768 13263 778
rect 13587 648 13599 778
rect 13707 456 13719 778
rect 13779 456 13791 778
rect 13827 648 13839 778
rect 14163 336 14175 778
rect 14211 528 14223 778
rect 14403 456 14415 778
rect 14931 648 14943 778
rect 14955 456 14967 778
rect 15003 120 15015 778
rect 15027 528 15039 778
rect 15075 528 15087 778
rect 15147 408 15159 778
rect 15291 408 15303 778
rect 15363 528 15375 778
rect 15531 768 15543 778
rect 15699 240 15711 778
rect 15819 480 15831 778
rect 15915 480 15927 778
rect 16059 600 16071 778
rect 16083 576 16095 778
rect 16491 576 16503 778
rect 16779 600 16791 778
rect 16899 648 16911 778
rect 17643 600 17655 778
rect 17691 192 17703 778
rect 17859 384 17871 778
rect 18123 600 18135 778
rect 18171 168 18183 778
rect 18507 552 18519 778
rect 18603 288 18615 778
rect 19131 672 19143 778
rect 19659 648 19671 778
rect 19947 720 19959 778
rect 20043 600 20055 778
rect 20139 456 20151 778
rect 20355 744 20367 778
rect 20403 360 20415 778
rect 20451 96 20463 778
rect 20547 456 20559 778
rect 20595 216 20607 778
rect 21099 552 21111 778
rect 21387 600 21399 778
rect 21915 696 21927 778
rect 21963 480 21975 778
rect 22011 576 22023 778
rect 22131 480 22143 778
rect 22587 576 22599 778
rect 22659 456 22671 778
rect 22779 48 22791 778
rect 22899 552 22911 778
rect 22995 144 23007 778
rect 23139 528 23151 778
rect 23259 456 23271 778
rect 23403 408 23415 778
rect 23499 72 23511 778
rect 23667 456 23679 778
rect 23691 312 23703 778
rect 23907 408 23919 778
rect 23955 600 23967 778
rect 23979 576 23991 778
rect 24483 432 24495 778
rect 26115 672 26127 778
rect 26187 624 26199 778
rect 26379 504 26391 778
rect 23920 394 23938 408
rect 14427 0 14439 10
rect 23919 0 23931 394
rect 26667 264 26679 778
rect 26715 408 26727 778
rect 26763 432 26775 778
rect 26811 456 26823 778
rect 26811 48 26823 394
rect 26835 24 26847 466
rect 26859 72 26871 442
rect 27387 0 27587 778
rect 27665 419 27735 431
rect 27665 59 27735 71
rect 27665 35 27735 47
rect 27665 11 27735 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 7083
box 0 0 1464 799
use inv g8182
timestamp 1386238110
transform 1 0 1587 0 1 7083
box 0 0 120 799
use rowcrosser StatusRegEn
timestamp 1386086759
transform 1 0 1707 0 1 7083
box 0 0 48 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 1755 0 1 7083
box 0 0 48 799
use and2 g8369
timestamp 1386234845
transform 1 0 1803 0 1 7083
box 0 0 120 799
use inv g8462
timestamp 1386238110
transform 1 0 1923 0 1 7083
box 0 0 120 799
use inv g8169
timestamp 1386238110
transform 1 0 2043 0 1 7083
box 0 0 120 799
use inv g8469
timestamp 1386238110
transform 1 0 2163 0 1 7083
box 0 0 120 799
use nand2 g8229
timestamp 1386234792
transform 1 0 2283 0 1 7083
box 0 0 96 799
use nand2 g8107
timestamp 1386234792
transform 1 0 2379 0 1 7083
box 0 0 96 799
use nand4 g8370
timestamp 1386234936
transform 1 0 2475 0 1 7083
box 0 0 144 799
use nand2 g8313
timestamp 1386234792
transform 1 0 2619 0 1 7083
box 0 0 96 799
use and2 g8344
timestamp 1386234845
transform 1 0 2715 0 1 7083
box 0 0 120 799
use inv g8123
timestamp 1386238110
transform 1 0 2835 0 1 7083
box 0 0 120 799
use nand4 g8222
timestamp 1386234936
transform 1 0 2955 0 1 7083
box 0 0 144 799
use nand2 g8098
timestamp 1386234792
transform 1 0 3099 0 1 7083
box 0 0 96 799
use nand4 g8314
timestamp 1386234936
transform 1 0 3195 0 1 7083
box 0 0 144 799
use nand2 g8327
timestamp 1386234792
transform 1 0 3339 0 1 7083
box 0 0 96 799
use nand2 g8187
timestamp 1386234792
transform 1 0 3435 0 1 7083
box 0 0 96 799
use nand2 g8477
timestamp 1386234792
transform 1 0 3531 0 1 7083
box 0 0 96 799
use nand2 g8171
timestamp 1386234792
transform 1 0 3627 0 1 7083
box 0 0 96 799
use nand2 g8135
timestamp 1386234792
transform 1 0 3723 0 1 7083
box 0 0 96 799
use nand4 g8295
timestamp 1386234936
transform 1 0 3819 0 1 7083
box 0 0 144 799
use nand3 g8287
timestamp 1386234893
transform 1 0 3963 0 1 7083
box 0 0 120 799
use nand2 g8154
timestamp 1386234792
transform 1 0 4083 0 1 7083
box 0 0 96 799
use nand4 g8276
timestamp 1386234936
transform 1 0 4179 0 1 7083
box 0 0 144 799
use nand2 g8261
timestamp 1386234792
transform 1 0 4323 0 1 7083
box 0 0 96 799
use nand3 g8130
timestamp 1386234893
transform 1 0 4419 0 1 7083
box 0 0 120 799
use nand2 g8318
timestamp 1386234792
transform 1 0 4539 0 1 7083
box 0 0 96 799
use nand2 g8377
timestamp 1386234792
transform 1 0 4635 0 1 7083
box 0 0 96 799
use nand2 g8474
timestamp 1386234792
transform 1 0 4731 0 1 7083
box 0 0 96 799
use nor2 g8390
timestamp 1386235306
transform 1 0 4827 0 1 7083
box 0 0 120 799
use nand2 g8168
timestamp 1386234792
transform 1 0 4947 0 1 7083
box 0 0 96 799
use nand2 g8238
timestamp 1386234792
transform 1 0 5043 0 1 7083
box 0 0 96 799
use nand2 g8225
timestamp 1386234792
transform 1 0 5139 0 1 7083
box 0 0 96 799
use nand2 g8143
timestamp 1386234792
transform 1 0 5235 0 1 7083
box 0 0 96 799
use nand2 g8333
timestamp 1386234792
transform 1 0 5331 0 1 7083
box 0 0 96 799
use nand3 g8472
timestamp 1386234893
transform 1 0 5427 0 1 7083
box 0 0 120 799
use and2 g8149
timestamp 1386234845
transform 1 0 5547 0 1 7083
box 0 0 120 799
use nor2 g8338
timestamp 1386235306
transform 1 0 5667 0 1 7083
box 0 0 120 799
use nor2 g8280
timestamp 1386235306
transform 1 0 5787 0 1 7083
box 0 0 120 799
use nand2 g8249
timestamp 1386234792
transform 1 0 5907 0 1 7083
box 0 0 96 799
use nand2 g8310
timestamp 1386234792
transform 1 0 6003 0 1 7083
box 0 0 96 799
use nand2 g8456
timestamp 1386234792
transform 1 0 6099 0 1 7083
box 0 0 96 799
use inv g8450
timestamp 1386238110
transform 1 0 6195 0 1 7083
box 0 0 120 799
use and2 g8235
timestamp 1386234845
transform 1 0 6315 0 1 7083
box 0 0 120 799
use nand4 g8362
timestamp 1386234936
transform 1 0 6435 0 1 7083
box 0 0 144 799
use nand2 g8214
timestamp 1386234792
transform 1 0 6579 0 1 7083
box 0 0 96 799
use nand2 g8281
timestamp 1386234792
transform 1 0 6675 0 1 7083
box 0 0 96 799
use nand3 g8366
timestamp 1386234893
transform 1 0 6771 0 1 7083
box 0 0 120 799
use nand2 g8269
timestamp 1386234792
transform 1 0 6891 0 1 7083
box 0 0 96 799
use inv g8440
timestamp 1386238110
transform 1 0 6987 0 1 7083
box 0 0 120 799
use nand2 g8183
timestamp 1386234792
transform 1 0 7107 0 1 7083
box 0 0 96 799
use nand3 g8170
timestamp 1386234893
transform 1 0 7203 0 1 7083
box 0 0 120 799
use nand3 g8449
timestamp 1386234893
transform 1 0 7323 0 1 7083
box 0 0 120 799
use nand2 g8124
timestamp 1386234792
transform 1 0 7443 0 1 7083
box 0 0 96 799
use nand4 g8106
timestamp 1386234936
transform 1 0 7539 0 1 7083
box 0 0 144 799
use nand4 g8414
timestamp 1386234936
transform 1 0 7683 0 1 7083
box 0 0 144 799
use nand2 g8119
timestamp 1386234792
transform 1 0 7827 0 1 7083
box 0 0 96 799
use nand4 g8275
timestamp 1386234936
transform 1 0 7923 0 1 7083
box 0 0 144 799
use and2 g8418
timestamp 1386234845
transform 1 0 8067 0 1 7083
box 0 0 120 799
use nand2 g8146
timestamp 1386234792
transform 1 0 8187 0 1 7083
box 0 0 96 799
use nand4 g8155
timestamp 1386234936
transform 1 0 8283 0 1 7083
box 0 0 144 799
use nand2 g8127
timestamp 1386234792
transform 1 0 8427 0 1 7083
box 0 0 96 799
use nand2 g8290
timestamp 1386234792
transform 1 0 8523 0 1 7083
box 0 0 96 799
use and2 g8252
timestamp 1386234845
transform 1 0 8619 0 1 7083
box 0 0 120 799
use nand2 g8334
timestamp 1386234792
transform 1 0 8739 0 1 7083
box 0 0 96 799
use nand4 g8244
timestamp 1386234936
transform 1 0 8835 0 1 7083
box 0 0 144 799
use nand4 g8240
timestamp 1386234936
transform 1 0 8979 0 1 7083
box 0 0 144 799
use nand4 g8407
timestamp 1386234936
transform 1 0 9123 0 1 7083
box 0 0 144 799
use nand2 g8139
timestamp 1386234792
transform 1 0 9267 0 1 7083
box 0 0 96 799
use nand3 g8118
timestamp 1386234893
transform 1 0 9363 0 1 7083
box 0 0 120 799
use nand4 g8363
timestamp 1386234936
transform 1 0 9483 0 1 7083
box 0 0 144 799
use and2 g8489
timestamp 1386234845
transform 1 0 9627 0 1 7083
box 0 0 120 799
use rowcrosser nME
timestamp 1386086759
transform 1 0 9747 0 1 7083
box 0 0 48 799
use inv g8111
timestamp 1386238110
transform 1 0 9795 0 1 7083
box 0 0 120 799
use nand3 g8381
timestamp 1386234893
transform 1 0 9915 0 1 7083
box 0 0 120 799
use and2 g8403
timestamp 1386234845
transform 1 0 10035 0 1 7083
box 0 0 120 799
use nand2 g8347
timestamp 1386234792
transform 1 0 10155 0 1 7083
box 0 0 96 799
use nand2 g8357
timestamp 1386234792
transform 1 0 10251 0 1 7083
box 0 0 96 799
use inv g8134
timestamp 1386238110
transform 1 0 10347 0 1 7083
box 0 0 120 799
use inv g8386
timestamp 1386238110
transform 1 0 10467 0 1 7083
box 0 0 120 799
use nand2 g8425
timestamp 1386234792
transform 1 0 10587 0 1 7083
box 0 0 96 799
use rowcrosser Flags_91_3_93_
timestamp 1386086759
transform 1 0 10683 0 1 7083
box 0 0 48 799
use and2 g8320
timestamp 1386234845
transform 1 0 10731 0 1 7083
box 0 0 120 799
use inv g8374
timestamp 1386238110
transform 1 0 10851 0 1 7083
box 0 0 120 799
use inv g8354
timestamp 1386238110
transform 1 0 10971 0 1 7083
box 0 0 120 799
use nor2 g8479
timestamp 1386235306
transform 1 0 11091 0 1 7083
box 0 0 120 799
use nor2 g8218
timestamp 1386235306
transform 1 0 11211 0 1 7083
box 0 0 120 799
use and2 g8284
timestamp 1386234845
transform 1 0 11331 0 1 7083
box 0 0 120 799
use rowcrosser Flags_91_0_93_
timestamp 1386086759
transform 1 0 11451 0 1 7083
box 0 0 48 799
use nand2 g8198
timestamp 1386234792
transform 1 0 11499 0 1 7083
box 0 0 96 799
use nand3 g8272
timestamp 1386234893
transform 1 0 11595 0 1 7083
box 0 0 120 799
use nand2 g8306
timestamp 1386234792
transform 1 0 11715 0 1 7083
box 0 0 96 799
use nand2 g8221
timestamp 1386234792
transform 1 0 11811 0 1 7083
box 0 0 96 799
use nand2 g8319
timestamp 1386234792
transform 1 0 11907 0 1 7083
box 0 0 96 799
use rowcrosser LrWe
timestamp 1386086759
transform 1 0 12003 0 1 7083
box 0 0 48 799
use and2 g8220
timestamp 1386234845
transform 1 0 12051 0 1 7083
box 0 0 120 799
use nand2 g8431
timestamp 1386234792
transform 1 0 12171 0 1 7083
box 0 0 96 799
use nand2 g8392
timestamp 1386234792
transform 1 0 12267 0 1 7083
box 0 0 96 799
use and2 g8230
timestamp 1386234845
transform 1 0 12363 0 1 7083
box 0 0 120 799
use rowcrosser AluWe
timestamp 1386086759
transform 1 0 12483 0 1 7083
box 0 0 48 799
use nand2 g8194
timestamp 1386234792
transform 1 0 12531 0 1 7083
box 0 0 96 799
use and2 g8271
timestamp 1386234845
transform 1 0 12627 0 1 7083
box 0 0 120 799
use nand2 g8340
timestamp 1386234792
transform 1 0 12747 0 1 7083
box 0 0 96 799
use nand2 rm_assigns_buf_StatusReg_1
timestamp 1386234792
transform 1 0 12843 0 1 7083
box 0 0 96 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 12939 0 1 7083
box 0 0 48 799
use buffer g8421
timestamp 1386236986
transform 1 0 12987 0 1 7083
box 0 0 120 799
use and2 g8399
timestamp 1386234845
transform 1 0 13107 0 1 7083
box 0 0 120 799
use nand3 g8209
timestamp 1386234893
transform 1 0 13227 0 1 7083
box 0 0 120 799
use nand2 g8283
timestamp 1386234792
transform 1 0 13347 0 1 7083
box 0 0 96 799
use nor2 g8268
timestamp 1386235306
transform 1 0 13443 0 1 7083
box 0 0 120 799
use and2 g8411
timestamp 1386234845
transform 1 0 13563 0 1 7083
box 0 0 120 799
use nand3 g8321
timestamp 1386234893
transform 1 0 13683 0 1 7083
box 0 0 120 799
use nand2 g8379
timestamp 1386234792
transform 1 0 13803 0 1 7083
box 0 0 96 799
use and2 g8180
timestamp 1386234845
transform 1 0 13899 0 1 7083
box 0 0 120 799
use and2 g8417
timestamp 1386234845
transform 1 0 14019 0 1 7083
box 0 0 120 799
use and2 g8136
timestamp 1386234845
transform 1 0 14139 0 1 7083
box 0 0 120 799
use inv g8110
timestamp 1386238110
transform 1 0 14259 0 1 7083
box 0 0 120 799
use rowcrosser stateSub_reg_91_0_93_
timestamp 1386086759
transform 1 0 14379 0 1 7083
box 0 0 48 799
use nand3 g8153
timestamp 1386234893
transform 1 0 14427 0 1 7083
box 0 0 120 799
use inv g8361
timestamp 1386238110
transform 1 0 14547 0 1 7083
box 0 0 120 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 14667 0 1 7083
box 0 0 96 799
use scandtype g8308
timestamp 1386241841
transform 1 0 14763 0 1 7083
box 0 0 624 799
use rowcrosser Op2Sel_91_0_93_
timestamp 1386086759
transform 1 0 15387 0 1 7083
box 0 0 48 799
use nand2 stateSub_reg_91_2_93_
timestamp 1386234792
transform 1 0 15435 0 1 7083
box 0 0 96 799
use scandtype g8372
timestamp 1386241841
transform 1 0 15531 0 1 7083
box 0 0 624 799
use rowcrosser MemEn
timestamp 1386086759
transform 1 0 16155 0 1 7083
box 0 0 48 799
use nand2 g8294
timestamp 1386234792
transform 1 0 16203 0 1 7083
box 0 0 96 799
use nand3 g8444
timestamp 1386234893
transform 1 0 16299 0 1 7083
box 0 0 120 799
use nor2 g8466
timestamp 1386235306
transform 1 0 16419 0 1 7083
box 0 0 120 799
use and2 g8433
timestamp 1386234845
transform 1 0 16539 0 1 7083
box 0 0 120 799
use nand3 g8468
timestamp 1386234893
transform 1 0 16659 0 1 7083
box 0 0 120 799
use nand2 g8420
timestamp 1386234792
transform 1 0 16779 0 1 7083
box 0 0 96 799
use nand2 g8190
timestamp 1386234792
transform 1 0 16875 0 1 7083
box 0 0 96 799
use nand2 g8304
timestamp 1386234792
transform 1 0 16971 0 1 7083
box 0 0 96 799
use nand2 g8277
timestamp 1386234792
transform 1 0 17067 0 1 7083
box 0 0 96 799
use nand2 g8243
timestamp 1386234792
transform 1 0 17163 0 1 7083
box 0 0 96 799
use inv g8296
timestamp 1386238110
transform 1 0 17259 0 1 7083
box 0 0 120 799
use nand3 g8348
timestamp 1386234893
transform 1 0 17379 0 1 7083
box 0 0 120 799
use nand2 g8234
timestamp 1386234792
transform 1 0 17499 0 1 7083
box 0 0 96 799
use and2 StatusReg_reg_91_1_93_
timestamp 1386234845
transform 1 0 17595 0 1 7083
box 0 0 120 799
use scandtype g8324
timestamp 1386241841
transform 1 0 17715 0 1 7083
box 0 0 624 799
use nand2 g8293
timestamp 1386234792
transform 1 0 18339 0 1 7083
box 0 0 96 799
use nand3 g8435
timestamp 1386234893
transform 1 0 18435 0 1 7083
box 0 0 120 799
use xor2 g8452
timestamp 1386237344
transform 1 0 18555 0 1 7083
box 0 0 192 799
use nand2 g8312
timestamp 1386234792
transform 1 0 18747 0 1 7083
box 0 0 96 799
use and2 g8213
timestamp 1386234845
transform 1 0 18843 0 1 7083
box 0 0 120 799
use nand2 g8212
timestamp 1386234792
transform 1 0 18963 0 1 7083
box 0 0 96 799
use nand2 g8265
timestamp 1386234792
transform 1 0 19059 0 1 7083
box 0 0 96 799
use nand3 g8200
timestamp 1386234893
transform 1 0 19155 0 1 7083
box 0 0 120 799
use nor2 g8400
timestamp 1386235306
transform 1 0 19275 0 1 7083
box 0 0 120 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 19395 0 1 7083
box 0 0 48 799
use inv g8108
timestamp 1386238110
transform 1 0 19443 0 1 7083
box 0 0 120 799
use and2 g8159
timestamp 1386234845
transform 1 0 19563 0 1 7083
box 0 0 120 799
use nor2 g8144
timestamp 1386235306
transform 1 0 19683 0 1 7083
box 0 0 120 799
use nand2 g8177
timestamp 1386234792
transform 1 0 19803 0 1 7083
box 0 0 96 799
use nand2 g8356
timestamp 1386234792
transform 1 0 19899 0 1 7083
box 0 0 96 799
use nand2 g8251
timestamp 1386234792
transform 1 0 19995 0 1 7083
box 0 0 96 799
use nand2 g8226
timestamp 1386234792
transform 1 0 20091 0 1 7083
box 0 0 96 799
use rowcrosser LrSel
timestamp 1386086759
transform 1 0 20187 0 1 7083
box 0 0 48 799
use and2 g8480
timestamp 1386234845
transform 1 0 20235 0 1 7083
box 0 0 120 799
use inv g8436
timestamp 1386238110
transform 1 0 20355 0 1 7083
box 0 0 120 799
use nand2 g8264
timestamp 1386234792
transform 1 0 20475 0 1 7083
box 0 0 96 799
use and2 g8332
timestamp 1386234845
transform 1 0 20571 0 1 7083
box 0 0 120 799
use nand4 g8206
timestamp 1386234936
transform 1 0 20691 0 1 7083
box 0 0 144 799
use nand2 g8237
timestamp 1386234792
transform 1 0 20835 0 1 7083
box 0 0 96 799
use nand2 g8278
timestamp 1386234792
transform 1 0 20931 0 1 7083
box 0 0 96 799
use nand2 g8376
timestamp 1386234792
transform 1 0 21027 0 1 7083
box 0 0 96 799
use nand2 g8181
timestamp 1386234792
transform 1 0 21123 0 1 7083
box 0 0 96 799
use nand2 g8216
timestamp 1386234792
transform 1 0 21219 0 1 7083
box 0 0 96 799
use inv StatusReg_reg_91_0_93_
timestamp 1386238110
transform 1 0 21315 0 1 7083
box 0 0 120 799
use scandtype g8253
timestamp 1386241841
transform 1 0 21435 0 1 7083
box 0 0 624 799
use nand2 g8373
timestamp 1386234792
transform 1 0 22059 0 1 7083
box 0 0 96 799
use nand3 g8443
timestamp 1386234893
transform 1 0 22155 0 1 7083
box 0 0 120 799
use inv g8186
timestamp 1386238110
transform 1 0 22275 0 1 7083
box 0 0 120 799
use nor2 g8427
timestamp 1386235306
transform 1 0 22395 0 1 7083
box 0 0 120 799
use nand2 g8432
timestamp 1386234792
transform 1 0 22515 0 1 7083
box 0 0 96 799
use nand2 g8424
timestamp 1386234792
transform 1 0 22611 0 1 7083
box 0 0 96 799
use nand2 g8195
timestamp 1386234792
transform 1 0 22707 0 1 7083
box 0 0 96 799
use nand3 g8223
timestamp 1386234893
transform 1 0 22803 0 1 7083
box 0 0 120 799
use nand2 g8410
timestamp 1386234792
transform 1 0 22923 0 1 7083
box 0 0 96 799
use and2 g8133
timestamp 1386234845
transform 1 0 23019 0 1 7083
box 0 0 120 799
use nand4 g8341
timestamp 1386234936
transform 1 0 23139 0 1 7083
box 0 0 144 799
use nand2 g8495
timestamp 1386234792
transform 1 0 23283 0 1 7083
box 0 0 96 799
use inv g8406
timestamp 1386238110
transform 1 0 23379 0 1 7083
box 0 0 120 799
use inv g8289
timestamp 1386238110
transform 1 0 23499 0 1 7083
box 0 0 120 799
use nand3 g8128
timestamp 1386234893
transform 1 0 23619 0 1 7083
box 0 0 120 799
use nand2 g8397
timestamp 1386234792
transform 1 0 23739 0 1 7083
box 0 0 96 799
use nand2 g8350
timestamp 1386234792
transform 1 0 23835 0 1 7083
box 0 0 96 799
use nand2 g8117
timestamp 1386234792
transform 1 0 23931 0 1 7083
box 0 0 96 799
use nand3 g8167
timestamp 1386234893
transform 1 0 24027 0 1 7083
box 0 0 120 799
use nand2 g8439
timestamp 1386234792
transform 1 0 24147 0 1 7083
box 0 0 96 799
use nand2 g8191
timestamp 1386234792
transform 1 0 24243 0 1 7083
box 0 0 96 799
use and2 g8227
timestamp 1386234845
transform 1 0 24339 0 1 7083
box 0 0 120 799
use nand4 g8473
timestamp 1386234936
transform 1 0 24459 0 1 7083
box 0 0 144 799
use nand2 g8387
timestamp 1386234792
transform 1 0 24603 0 1 7083
box 0 0 96 799
use nor2 g8270
timestamp 1386235306
transform 1 0 24699 0 1 7083
box 0 0 120 799
use nand2 g8465
timestamp 1386234792
transform 1 0 24819 0 1 7083
box 0 0 96 799
use nand2 g8163
timestamp 1386234792
transform 1 0 24915 0 1 7083
box 0 0 96 799
use nand3 g8455
timestamp 1386234893
transform 1 0 25011 0 1 7083
box 0 0 120 799
use and2 g8273
timestamp 1386234845
transform 1 0 25131 0 1 7083
box 0 0 120 799
use nand2 g8337
timestamp 1386234792
transform 1 0 25251 0 1 7083
box 0 0 96 799
use inv g8478
timestamp 1386238110
transform 1 0 25347 0 1 7083
box 0 0 120 799
use and2 g8147
timestamp 1386234845
transform 1 0 25467 0 1 7083
box 0 0 120 799
use nand2 g8217
timestamp 1386234792
transform 1 0 25587 0 1 7083
box 0 0 96 799
use nand2 g8367
timestamp 1386234792
transform 1 0 25683 0 1 7083
box 0 0 96 799
use nand2 g8353
timestamp 1386234792
transform 1 0 25779 0 1 7083
box 0 0 96 799
use nand2 g8248
timestamp 1386234792
transform 1 0 25875 0 1 7083
box 0 0 96 799
use nand2 g8447
timestamp 1386234792
transform 1 0 25971 0 1 7083
box 0 0 96 799
use nand2 g8114
timestamp 1386234792
transform 1 0 26067 0 1 7083
box 0 0 96 799
use nand3 g8174
timestamp 1386234893
transform 1 0 26163 0 1 7083
box 0 0 120 799
use nand2 g8393
timestamp 1386234792
transform 1 0 26283 0 1 7083
box 0 0 96 799
use nand2 g8305
timestamp 1386234792
transform 1 0 26379 0 1 7083
box 0 0 96 799
use nand2 g8241
timestamp 1386234792
transform 1 0 26475 0 1 7083
box 0 0 96 799
use nand4 g8382
timestamp 1386234936
transform 1 0 26571 0 1 7083
box 0 0 144 799
use nand2 g8158
timestamp 1386234792
transform 1 0 26715 0 1 7083
box 0 0 96 799
use nor2 g8257
timestamp 1386235306
transform 1 0 26811 0 1 7083
box 0 0 120 799
use nor2 g8451
timestamp 1386235306
transform 1 0 26931 0 1 7083
box 0 0 120 799
use inv PcSel_91_1_93_
timestamp 1386238110
transform 1 0 27051 0 1 7083
box 0 0 120 799
use rowcrosser PcSel_91_0_93_
timestamp 1386086759
transform 1 0 27171 0 1 7083
box 0 0 48 799
use rowcrosser ALE
timestamp 1386086759
transform 1 0 27219 0 1 7083
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27267 0 1 7083
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 778
box 0 0 1464 799
use scandtype g8409
timestamp 1386241841
transform 1 0 1587 0 1 778
box 0 0 624 799
use rowcrosser SysBus_91_2_93_
timestamp 1386086759
transform 1 0 2211 0 1 778
box 0 0 48 799
use and2 g8352
timestamp 1386234845
transform 1 0 2259 0 1 778
box 0 0 120 799
use nand2 g8430
timestamp 1386234792
transform 1 0 2379 0 1 778
box 0 0 96 799
use nand2 g8150
timestamp 1386234792
transform 1 0 2475 0 1 778
box 0 0 96 799
use nand3 g8178
timestamp 1386234893
transform 1 0 2571 0 1 778
box 0 0 120 799
use and2 g8250
timestamp 1386234845
transform 1 0 2691 0 1 778
box 0 0 120 799
use nand2 state_reg_91_1_93_
timestamp 1386234792
transform 1 0 2811 0 1 778
box 0 0 96 799
use scandtype g8416
timestamp 1386241841
transform 1 0 2907 0 1 778
box 0 0 624 799
use rowcrosser SysBus_91_0_93_
timestamp 1386086759
transform 1 0 3531 0 1 778
box 0 0 48 799
use nand2 g8148
timestamp 1386234792
transform 1 0 3579 0 1 778
box 0 0 96 799
use nand3 g8434
timestamp 1386234893
transform 1 0 3675 0 1 778
box 0 0 120 799
use mux2 g8211
timestamp 1386235218
transform 1 0 3795 0 1 778
box 0 0 192 799
use nand2 g8196
timestamp 1386234792
transform 1 0 3987 0 1 778
box 0 0 96 799
use nand2 g8300
timestamp 1386234792
transform 1 0 4083 0 1 778
box 0 0 96 799
use and2 g8175
timestamp 1386234845
transform 1 0 4179 0 1 778
box 0 0 120 799
use nand2 g8359
timestamp 1386234792
transform 1 0 4299 0 1 778
box 0 0 96 799
use nand3 g8429
timestamp 1386234893
transform 1 0 4395 0 1 778
box 0 0 120 799
use inv g8104
timestamp 1386238110
transform 1 0 4515 0 1 778
box 0 0 120 799
use nor2 g8391
timestamp 1386235306
transform 1 0 4635 0 1 778
box 0 0 120 799
use nand2 g8307
timestamp 1386234792
transform 1 0 4755 0 1 778
box 0 0 96 799
use inv g8389
timestamp 1386238110
transform 1 0 4851 0 1 778
box 0 0 120 799
use nand2 g8458
timestamp 1386234792
transform 1 0 4971 0 1 778
box 0 0 96 799
use inv g8335
timestamp 1386238110
transform 1 0 5067 0 1 778
box 0 0 120 799
use nand2 g8160
timestamp 1386234792
transform 1 0 5187 0 1 778
box 0 0 96 799
use nand3 g8476
timestamp 1386234893
transform 1 0 5283 0 1 778
box 0 0 120 799
use inv g8161
timestamp 1386238110
transform 1 0 5403 0 1 778
box 0 0 120 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 5523 0 1 778
box 0 0 96 799
use scandtype g8224
timestamp 1386241841
transform 1 0 5619 0 1 778
box 0 0 624 799
use nand2 g8266
timestamp 1386234792
transform 1 0 6243 0 1 778
box 0 0 96 799
use nand2 g8401
timestamp 1386234792
transform 1 0 6339 0 1 778
box 0 0 96 799
use nand2 g8189
timestamp 1386234792
transform 1 0 6435 0 1 778
box 0 0 96 799
use nand2 g8125
timestamp 1386234792
transform 1 0 6531 0 1 778
box 0 0 96 799
use nand4 g8454
timestamp 1386234936
transform 1 0 6627 0 1 778
box 0 0 144 799
use nor2 g8442
timestamp 1386235306
transform 1 0 6771 0 1 778
box 0 0 120 799
use nor2 g8297
timestamp 1386235306
transform 1 0 6891 0 1 778
box 0 0 120 799
use nand2 g8232
timestamp 1386234792
transform 1 0 7011 0 1 778
box 0 0 96 799
use nand2 g8152
timestamp 1386234792
transform 1 0 7107 0 1 778
box 0 0 96 799
use nand4 g8328
timestamp 1386234936
transform 1 0 7203 0 1 778
box 0 0 144 799
use nand3 g8303
timestamp 1386234893
transform 1 0 7347 0 1 778
box 0 0 120 799
use nor2 g8394
timestamp 1386235306
transform 1 0 7467 0 1 778
box 0 0 120 799
use nand2 g8395
timestamp 1386234792
transform 1 0 7587 0 1 778
box 0 0 96 799
use nor2 g8453
timestamp 1386235306
transform 1 0 7683 0 1 778
box 0 0 120 799
use nand2 g8267
timestamp 1386234792
transform 1 0 7803 0 1 778
box 0 0 96 799
use nand2 g8282
timestamp 1386234792
transform 1 0 7899 0 1 778
box 0 0 96 799
use inv g8461
timestamp 1386238110
transform 1 0 7995 0 1 778
box 0 0 120 799
use nor2 g8274
timestamp 1386235306
transform 1 0 8115 0 1 778
box 0 0 120 799
use nand2 g8236
timestamp 1386234792
transform 1 0 8235 0 1 778
box 0 0 96 799
use nand2 g8438
timestamp 1386234792
transform 1 0 8331 0 1 778
box 0 0 96 799
use nand2 g8349
timestamp 1386234792
transform 1 0 8427 0 1 778
box 0 0 96 799
use and2 g8412
timestamp 1386234845
transform 1 0 8523 0 1 778
box 0 0 120 799
use and2 g8481
timestamp 1386234845
transform 1 0 8643 0 1 778
box 0 0 120 799
use inv g8185
timestamp 1386238110
transform 1 0 8763 0 1 778
box 0 0 120 799
use nand2 g8365
timestamp 1386234792
transform 1 0 8883 0 1 778
box 0 0 96 799
use nand2 g8255
timestamp 1386234792
transform 1 0 8979 0 1 778
box 0 0 96 799
use inv g8457
timestamp 1386238110
transform 1 0 9075 0 1 778
box 0 0 120 799
use nand2 g8301
timestamp 1386234792
transform 1 0 9195 0 1 778
box 0 0 96 799
use nand2 g8192
timestamp 1386234792
transform 1 0 9291 0 1 778
box 0 0 96 799
use nand3 g8292
timestamp 1386234893
transform 1 0 9387 0 1 778
box 0 0 120 799
use nand3 g8254
timestamp 1386234893
transform 1 0 9507 0 1 778
box 0 0 120 799
use nand2 g8116
timestamp 1386234792
transform 1 0 9627 0 1 778
box 0 0 96 799
use nor2 g8470
timestamp 1386235306
transform 1 0 9723 0 1 778
box 0 0 120 799
use nand2 g8145
timestamp 1386234792
transform 1 0 9843 0 1 778
box 0 0 96 799
use nand2 g8166
timestamp 1386234792
transform 1 0 9939 0 1 778
box 0 0 96 799
use nand2 g8426
timestamp 1386234792
transform 1 0 10035 0 1 778
box 0 0 96 799
use inv g8315
timestamp 1386238110
transform 1 0 10131 0 1 778
box 0 0 120 799
use nand2 g8228
timestamp 1386234792
transform 1 0 10251 0 1 778
box 0 0 96 799
use nand3 g8342
timestamp 1386234893
transform 1 0 10347 0 1 778
box 0 0 120 799
use inv g8490
timestamp 1386238110
transform 1 0 10467 0 1 778
box 0 0 120 799
use inv g8279
timestamp 1386238110
transform 1 0 10587 0 1 778
box 0 0 120 799
use nand2 g8105
timestamp 1386234792
transform 1 0 10707 0 1 778
box 0 0 96 799
use nand4 g8259
timestamp 1386234936
transform 1 0 10803 0 1 778
box 0 0 144 799
use nand2 g8375
timestamp 1386234792
transform 1 0 10947 0 1 778
box 0 0 96 799
use nand2 g8129
timestamp 1386234792
transform 1 0 11043 0 1 778
box 0 0 96 799
use rowcrosser AluOR_91_1_93_
timestamp 1386086759
transform 1 0 11139 0 1 778
box 0 0 48 799
use nand2 g8446
timestamp 1386234792
transform 1 0 11187 0 1 778
box 0 0 96 799
use nand2 g8459
timestamp 1386234792
transform 1 0 11283 0 1 778
box 0 0 96 799
use nand2 g8097
timestamp 1386234792
transform 1 0 11379 0 1 778
box 0 0 96 799
use nand4 g8247
timestamp 1386234936
transform 1 0 11475 0 1 778
box 0 0 144 799
use nor2 g8263
timestamp 1386235306
transform 1 0 11619 0 1 778
box 0 0 120 799
use and2 IntStatus_reg
timestamp 1386234845
transform 1 0 11739 0 1 778
box 0 0 120 799
use scanreg g8256
timestamp 1386241447
transform 1 0 11859 0 1 778
box 0 0 720 799
use rowcrosser SysBus_91_3_93_
timestamp 1386086759
transform 1 0 12579 0 1 778
box 0 0 48 799
use nand2 g8131
timestamp 1386234792
transform 1 0 12627 0 1 778
box 0 0 96 799
use nand3 g8345
timestamp 1386234893
transform 1 0 12723 0 1 778
box 0 0 120 799
use nand2 g8491
timestamp 1386234792
transform 1 0 12843 0 1 778
box 0 0 96 799
use inv g8322
timestamp 1386238110
transform 1 0 12939 0 1 778
box 0 0 120 799
use and2 g8368
timestamp 1386234845
transform 1 0 13059 0 1 778
box 0 0 120 799
use nand2 g8286
timestamp 1386234792
transform 1 0 13179 0 1 778
box 0 0 96 799
use nand3 g8201
timestamp 1386234893
transform 1 0 13275 0 1 778
box 0 0 120 799
use nand2 g8137
timestamp 1386234792
transform 1 0 13395 0 1 778
box 0 0 96 799
use nand4 g8331
timestamp 1386234936
transform 1 0 13491 0 1 778
box 0 0 144 799
use nand2 g8336
timestamp 1386234792
transform 1 0 13635 0 1 778
box 0 0 96 799
use nor2 g8242
timestamp 1386235306
transform 1 0 13731 0 1 778
box 0 0 120 799
use nand3 g8207
timestamp 1386234893
transform 1 0 13851 0 1 778
box 0 0 120 799
use nor2 g8423
timestamp 1386235306
transform 1 0 13971 0 1 778
box 0 0 120 799
use nand2 g8383
timestamp 1386234792
transform 1 0 14091 0 1 778
box 0 0 96 799
use nand3 g8405
timestamp 1386234893
transform 1 0 14187 0 1 778
box 0 0 120 799
use and2 g8173
timestamp 1386234845
transform 1 0 14307 0 1 778
box 0 0 120 799
use nand3 g8398
timestamp 1386234893
transform 1 0 14427 0 1 778
box 0 0 120 799
use and2 g8464
timestamp 1386234845
transform 1 0 14547 0 1 778
box 0 0 120 799
use inv g8325
timestamp 1386238110
transform 1 0 14667 0 1 778
box 0 0 120 799
use and2 g8157
timestamp 1386234845
transform 1 0 14787 0 1 778
box 0 0 120 799
use nand4 g8140
timestamp 1386234936
transform 1 0 14907 0 1 778
box 0 0 144 799
use nor2 g8210
timestamp 1386235306
transform 1 0 15051 0 1 778
box 0 0 120 799
use nand2 g8141
timestamp 1386234792
transform 1 0 15171 0 1 778
box 0 0 96 799
use nand4 g8460
timestamp 1386234936
transform 1 0 15267 0 1 778
box 0 0 144 799
use nand2 g8317
timestamp 1386234792
transform 1 0 15411 0 1 778
box 0 0 96 799
use nand2 g8203
timestamp 1386234792
transform 1 0 15507 0 1 778
box 0 0 96 799
use and2 g8404
timestamp 1386234845
transform 1 0 15603 0 1 778
box 0 0 120 799
use and2 g8413
timestamp 1386234845
transform 1 0 15723 0 1 778
box 0 0 120 799
use nand2 g8428
timestamp 1386234792
transform 1 0 15843 0 1 778
box 0 0 96 799
use nand2 g8113
timestamp 1386234792
transform 1 0 15939 0 1 778
box 0 0 96 799
use nand3 g8358
timestamp 1386234893
transform 1 0 16035 0 1 778
box 0 0 120 799
use nand2 g8323
timestamp 1386234792
transform 1 0 16155 0 1 778
box 0 0 96 799
use inv g8408
timestamp 1386238110
transform 1 0 16251 0 1 778
box 0 0 120 799
use nand2 g8309
timestamp 1386234792
transform 1 0 16371 0 1 778
box 0 0 96 799
use nand2 g8380
timestamp 1386234792
transform 1 0 16467 0 1 778
box 0 0 96 799
use and2 g8233
timestamp 1386234845
transform 1 0 16563 0 1 778
box 0 0 120 799
use and2 IRQ2_reg
timestamp 1386234845
transform 1 0 16683 0 1 778
box 0 0 120 799
use scandtype g8151
timestamp 1386241841
transform 1 0 16803 0 1 778
box 0 0 624 799
use nand4 g8138
timestamp 1386234936
transform 1 0 17427 0 1 778
box 0 0 144 799
use nand4 g8402
timestamp 1386234936
transform 1 0 17571 0 1 778
box 0 0 144 799
use inv g8188
timestamp 1386238110
transform 1 0 17715 0 1 778
box 0 0 120 799
use inv g8176
timestamp 1386238110
transform 1 0 17835 0 1 778
box 0 0 120 799
use nor2 g8172
timestamp 1386235306
transform 1 0 17955 0 1 778
box 0 0 120 799
use nand3 g8422
timestamp 1386234893
transform 1 0 18075 0 1 778
box 0 0 120 799
use nand2 g8488
timestamp 1386234792
transform 1 0 18195 0 1 778
box 0 0 96 799
use inv g8162
timestamp 1386238110
transform 1 0 18291 0 1 778
box 0 0 120 799
use nand3 g8475
timestamp 1386234893
transform 1 0 18411 0 1 778
box 0 0 120 799
use nand2 g8415
timestamp 1386234792
transform 1 0 18531 0 1 778
box 0 0 96 799
use nand2 g8299
timestamp 1386234792
transform 1 0 18627 0 1 778
box 0 0 96 799
use and2 g8326
timestamp 1386234845
transform 1 0 18723 0 1 778
box 0 0 120 799
use nand2 g8126
timestamp 1386234792
transform 1 0 18843 0 1 778
box 0 0 96 799
use nand2 g8396
timestamp 1386234792
transform 1 0 18939 0 1 778
box 0 0 96 799
use nor2 IRQ1_reg
timestamp 1386235306
transform 1 0 19035 0 1 778
box 0 0 120 799
use scandtype g8329
timestamp 1386241841
transform 1 0 19155 0 1 778
box 0 0 624 799
use nand2 g8419
timestamp 1386234792
transform 1 0 19779 0 1 778
box 0 0 96 799
use nand2 g8205
timestamp 1386234792
transform 1 0 19875 0 1 778
box 0 0 96 799
use nand2 g8339
timestamp 1386234792
transform 1 0 19971 0 1 778
box 0 0 96 799
use inv g8463
timestamp 1386238110
transform 1 0 20067 0 1 778
box 0 0 120 799
use nand2 g8164
timestamp 1386234792
transform 1 0 20187 0 1 778
box 0 0 96 799
use nand2 g8245
timestamp 1386234792
transform 1 0 20283 0 1 778
box 0 0 96 799
use nand2 g8260
timestamp 1386234792
transform 1 0 20379 0 1 778
box 0 0 96 799
use nand2 g8165
timestamp 1386234792
transform 1 0 20475 0 1 778
box 0 0 96 799
use nand2 g8471
timestamp 1386234792
transform 1 0 20571 0 1 778
box 0 0 96 799
use nand2 g8351
timestamp 1386234792
transform 1 0 20667 0 1 778
box 0 0 96 799
use nand2 g8492
timestamp 1386234792
transform 1 0 20763 0 1 778
box 0 0 96 799
use inv g8343
timestamp 1386238110
transform 1 0 20859 0 1 778
box 0 0 120 799
use nand2 g8215
timestamp 1386234792
transform 1 0 20979 0 1 778
box 0 0 96 799
use nand2 g8288
timestamp 1386234792
transform 1 0 21075 0 1 778
box 0 0 96 799
use nand3 g8239
timestamp 1386234893
transform 1 0 21171 0 1 778
box 0 0 120 799
use nand3 g8384
timestamp 1386234893
transform 1 0 21291 0 1 778
box 0 0 120 799
use nand2 g8311
timestamp 1386234792
transform 1 0 21411 0 1 778
box 0 0 96 799
use nor2 g8262
timestamp 1386235306
transform 1 0 21507 0 1 778
box 0 0 120 799
use nand2 g8109
timestamp 1386234792
transform 1 0 21627 0 1 778
box 0 0 96 799
use nand3 g8298
timestamp 1386234893
transform 1 0 21723 0 1 778
box 0 0 120 799
use nand2 g8346
timestamp 1386234792
transform 1 0 21843 0 1 778
box 0 0 96 799
use nand2 g8184
timestamp 1386234792
transform 1 0 21939 0 1 778
box 0 0 96 799
use and2 g8355
timestamp 1386234845
transform 1 0 22035 0 1 778
box 0 0 120 799
use inv g8132
timestamp 1386238110
transform 1 0 22155 0 1 778
box 0 0 120 799
use inv g8385
timestamp 1386238110
transform 1 0 22275 0 1 778
box 0 0 120 799
use and2 g8330
timestamp 1386234845
transform 1 0 22395 0 1 778
box 0 0 120 799
use nand2 g8219
timestamp 1386234792
transform 1 0 22515 0 1 778
box 0 0 96 799
use and2 g8360
timestamp 1386234845
transform 1 0 22611 0 1 778
box 0 0 120 799
use nand2 g8258
timestamp 1386234792
transform 1 0 22731 0 1 778
box 0 0 96 799
use nand2 g8202
timestamp 1386234792
transform 1 0 22827 0 1 778
box 0 0 96 799
use nand2 g8246
timestamp 1386234792
transform 1 0 22923 0 1 778
box 0 0 96 799
use nand4 g8208
timestamp 1386234936
transform 1 0 23019 0 1 778
box 0 0 144 799
use nor2 g8231
timestamp 1386235306
transform 1 0 23163 0 1 778
box 0 0 120 799
use nand4 g8156
timestamp 1386234936
transform 1 0 23283 0 1 778
box 0 0 144 799
use nand2 g8467
timestamp 1386234792
transform 1 0 23427 0 1 778
box 0 0 96 799
use and2 g8179
timestamp 1386234845
transform 1 0 23523 0 1 778
box 0 0 120 799
use nor2 g8371
timestamp 1386235306
transform 1 0 23643 0 1 778
box 0 0 120 799
use and2 g8193
timestamp 1386234845
transform 1 0 23763 0 1 778
box 0 0 120 799
use rowcrosser RegWe
timestamp 1386086759
transform 1 0 23883 0 1 778
box 0 0 48 799
use and2 g8285
timestamp 1386234845
transform 1 0 23931 0 1 778
box 0 0 120 799
use nand3 g8485
timestamp 1386234893
transform 1 0 24051 0 1 778
box 0 0 120 799
use inv g8204
timestamp 1386238110
transform 1 0 24171 0 1 778
box 0 0 120 799
use nand2 state_reg_91_0_93_
timestamp 1386234792
transform 1 0 24291 0 1 778
box 0 0 96 799
use scandtype g8302
timestamp 1386241841
transform 1 0 24387 0 1 778
box 0 0 624 799
use nand2 g8142
timestamp 1386234792
transform 1 0 25011 0 1 778
box 0 0 96 799
use nand2 g8441
timestamp 1386234792
transform 1 0 25107 0 1 778
box 0 0 96 799
use inv stateSub_reg_91_1_93_
timestamp 1386238110
transform 1 0 25203 0 1 778
box 0 0 120 799
use scandtype g8316
timestamp 1386241841
transform 1 0 25323 0 1 778
box 0 0 624 799
use and2 g8197
timestamp 1386234845
transform 1 0 25947 0 1 778
box 0 0 120 799
use nand2 g8364
timestamp 1386234792
transform 1 0 26067 0 1 778
box 0 0 96 799
use nand2 g8378
timestamp 1386234792
transform 1 0 26163 0 1 778
box 0 0 96 799
use nand2 g8291
timestamp 1386234792
transform 1 0 26259 0 1 778
box 0 0 96 799
use inv g8112
timestamp 1386238110
transform 1 0 26355 0 1 778
box 0 0 120 799
use nand3 g8448
timestamp 1386234893
transform 1 0 26475 0 1 778
box 0 0 120 799
use nand2 SysBus_91_1_93_
timestamp 1386234792
transform 1 0 26595 0 1 778
box 0 0 96 799
use rowcrosser nIRQ
timestamp 1386086759
transform 1 0 26691 0 1 778
box 0 0 48 799
use rowcrosser AluOR_91_0_93_
timestamp 1386086759
transform 1 0 26739 0 1 778
box 0 0 48 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 26787 0 1 778
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27267 0 1 778
box 0 0 320 799
<< labels >>
rlabel m2contact 26865 449 26865 449 8 AluOR[0]
rlabel m2contact 26865 65 26865 65 8 AluOR[0]
rlabel m2contact 26841 473 26841 473 8 ENB
rlabel m2contact 26841 17 26841 17 8 ENB
rlabel m2contact 26817 401 26817 401 8 AluOR[1]
rlabel m2contact 26817 41 26817 41 8 AluOR[1]
rlabel m2contact 26817 449 26817 449 8 AluOR[0]
rlabel m2contact 26769 425 26769 425 8 RegWe
rlabel m2contact 26721 401 26721 401 8 AluOR[1]
rlabel m2contact 26673 257 26673 257 8 n_9
rlabel m2contact 26385 497 26385 497 8 n_155
rlabel m2contact 26193 617 26193 617 8 n_111
rlabel m2contact 26121 665 26121 665 8 n_147
rlabel m2contact 24489 425 24489 425 8 n_289
rlabel m2contact 23985 569 23985 569 8 n_131
rlabel m2contact 23961 593 23961 593 8 n_233
rlabel metal2 23931 401 23931 401 8 SysBus[3]
rlabel m2contact 23913 401 23913 401 8 SysBus[3]
rlabel m2contact 23697 305 23697 305 8 n_142
rlabel m2contact 23673 449 23673 449 8 n_242
rlabel m2contact 23505 65 23505 65 8 nWE
rlabel m2contact 23409 401 23409 401 8 n_191
rlabel m2contact 23265 449 23265 449 8 n_242
rlabel m2contact 23145 521 23145 521 8 n_254
rlabel m2contact 23001 137 23001 137 8 n_244
rlabel m2contact 22905 545 22905 545 8 n_140
rlabel m2contact 22785 41 22785 41 8 n_83
rlabel m2contact 22665 449 22665 449 8 n_251
rlabel m2contact 22593 569 22593 569 8 n_131
rlabel m2contact 22137 473 22137 473 8 ENB
rlabel m2contact 22017 569 22017 569 8 n_78
rlabel m2contact 21969 473 21969 473 8 n_48
rlabel m2contact 21921 689 21921 689 8 n_105
rlabel m2contact 21393 593 21393 593 8 n_233
rlabel m2contact 21105 545 21105 545 8 n_140
rlabel m2contact 20601 209 20601 209 8 n_295
rlabel m2contact 20553 449 20553 449 8 n_251
rlabel m2contact 20457 89 20457 89 8 n_143
rlabel m2contact 20409 353 20409 353 8 n_106
rlabel m2contact 20361 737 20361 737 8 n_327
rlabel m2contact 20145 449 20145 449 8 n_97
rlabel m2contact 20049 593 20049 593 8 n_272
rlabel m2contact 19953 713 19953 713 8 n_41
rlabel m2contact 19665 641 19665 641 8 IRQ1
rlabel m2contact 19137 665 19137 665 8 n_147
rlabel m2contact 18609 281 18609 281 8 n_4
rlabel m2contact 18513 545 18513 545 8 n_353
rlabel m2contact 18177 161 18177 161 8 n_321
rlabel m2contact 18129 593 18129 593 8 n_272
rlabel m2contact 17865 377 17865 377 8 n_315
rlabel m2contact 17697 185 17697 185 8 n_318
rlabel m2contact 17649 593 17649 593 8 n_258
rlabel m2contact 16905 641 16905 641 8 IRQ1
rlabel m2contact 16785 593 16785 593 8 n_258
rlabel m2contact 16497 569 16497 569 8 n_78
rlabel m2contact 16089 569 16089 569 8 n_325
rlabel m2contact 16065 593 16065 593 8 n_333
rlabel m2contact 15921 473 15921 473 8 n_48
rlabel m2contact 15825 473 15825 473 8 n_51
rlabel m2contact 15705 233 15705 233 8 n_204
rlabel m2contact 15537 761 15537 761 8 n_110
rlabel m2contact 15369 521 15369 521 8 n_254
rlabel m2contact 15297 401 15297 401 8 n_191
rlabel m2contact 15153 401 15153 401 8 n_274
rlabel m2contact 15081 521 15081 521 8 n_197
rlabel m2contact 15033 521 15033 521 8 n_197
rlabel m2contact 15009 113 15009 113 8 n_45
rlabel m2contact 14961 449 14961 449 8 n_97
rlabel m2contact 14937 641 14937 641 8 n_79
rlabel m2contact 14433 17 14433 17 8 SysBus[2]
rlabel m2contact 14409 449 14409 449 8 n_50
rlabel m2contact 14217 521 14217 521 8 n_13
rlabel m2contact 14169 329 14169 329 8 n_73
rlabel m2contact 13833 641 13833 641 2 n_79
rlabel m2contact 13785 449 13785 449 2 n_50
rlabel m2contact 13713 449 13713 449 2 n_164
rlabel m2contact 13593 641 13593 641 2 n_220
rlabel m2contact 13257 761 13257 761 2 n_110
rlabel m2contact 12801 545 12801 545 2 n_353
rlabel m2contact 12609 545 12609 545 2 SysBus[0]
rlabel m2contact 11937 737 11937 737 2 n_327
rlabel m2contact 11889 185 11889 185 2 n_318
rlabel m2contact 11721 305 11721 305 2 n_142
rlabel m2contact 11649 185 11649 185 2 n_98
rlabel m2contact 11553 305 11553 305 2 n_385
rlabel m2contact 11529 713 11529 713 2 n_41
rlabel m2contact 11265 569 11265 569 2 n_325
rlabel metal2 11187 569 11187 569 2 SysBus[1]
rlabel m2contact 11169 569 11169 569 2 SysBus[1]
rlabel m2contact 11073 617 11073 617 2 n_111
rlabel m2contact 10881 401 10881 401 2 n_274
rlabel m2contact 10785 401 10785 401 2 n_203
rlabel m2contact 10665 569 10665 569 2 n_3
rlabel m2contact 10377 689 10377 689 2 n_105
rlabel m2contact 10281 665 10281 665 2 n_147
rlabel m2contact 10209 617 10209 617 2 n_111
rlabel m2contact 10017 593 10017 593 2 n_333
rlabel m2contact 9921 593 9921 593 2 n_5
rlabel m2contact 9705 641 9705 641 2 n_220
rlabel m2contact 9609 497 9609 497 2 n_155
rlabel m2contact 9441 497 9441 497 2 n_102
rlabel m2contact 9417 233 9417 233 2 n_204
rlabel m2contact 9009 617 9009 617 2 n_111
rlabel m2contact 8673 593 8673 593 2 n_5
rlabel m2contact 8553 329 8553 329 2 n_73
rlabel m2contact 8505 329 8505 329 2 n_16
rlabel m2contact 8481 569 8481 569 2 n_3
rlabel m2contact 7989 545 7989 545 2 SysBus[0]
rlabel m2contact 7881 521 7881 521 2 n_13
rlabel m2contact 7569 497 7569 497 2 n_102
rlabel m2contact 7521 473 7521 473 2 n_51
rlabel m2contact 7449 185 7449 185 2 n_98
rlabel m2contact 7329 425 7329 425 2 n_289
rlabel m2contact 7305 185 7305 185 2 n_238
rlabel m2contact 7137 425 7137 425 2 n_217
rlabel m2contact 7089 353 7089 353 2 n_106
rlabel m2contact 7041 353 7041 353 2 n_57
rlabel m2contact 6657 449 6657 449 2 n_164
rlabel m2contact 6609 377 6609 377 2 n_315
rlabel m2contact 6417 425 6417 425 2 n_217
rlabel m2contact 6273 401 6273 401 2 n_203
rlabel m2contact 5553 377 5553 377 2 n_315
rlabel m2contact 5265 353 5265 353 2 n_57
rlabel m2contact 5241 329 5241 329 2 n_16
rlabel m2contact 5025 257 5025 257 2 n_9
rlabel m2contact 4833 257 4833 257 2 n_53
rlabel m2contact 4737 305 4737 305 2 n_385
rlabel m2contact 4545 41 4545 41 2 n_83
rlabel m2contact 4473 281 4473 281 2 n_4
rlabel m2contact 4353 257 4353 257 2 n_53
rlabel m2contact 4329 233 4329 233 2 n_204
rlabel m2contact 4161 209 4161 209 2 n_295
rlabel m2contact 4065 185 4065 185 2 n_238
rlabel m2contact 3729 161 3729 161 2 n_321
rlabel m2contact 3705 137 3705 137 2 n_244
rlabel m2contact 3657 113 3657 113 2 n_45
rlabel m2contact 3561 17 3561 17 2 SysBus[2]
rlabel m2contact 2553 41 2553 41 2 n_83
rlabel m2contact 2241 41 2241 41 2 nIRQ
rlabel m2contact 1689 89 1689 89 2 n_143
rlabel m2contact 27321 4282 27321 4282 6 Rs1Sel[1]
rlabel m2contact 27321 1642 27321 1642 6 Rs1Sel[1]
rlabel m2contact 27297 1786 27297 1786 6 RwSel[0]
rlabel m2contact 27297 1618 27297 1618 6 RwSel[0]
rlabel m2contact 27273 4354 27273 4354 6 RwSel[1]
rlabel m2contact 27273 1594 27273 1594 6 RwSel[1]
rlabel m2contact 27249 1714 27249 1714 6 Flags[3]
rlabel m2contact 27201 3994 27201 3994 6 StatusRegEn
rlabel m2contact 27129 4042 27129 4042 6 n_74
rlabel m2contact 27081 6178 27081 6178 6 n_287
rlabel m2contact 27033 4066 27033 4066 6 n_141
rlabel m2contact 26985 3490 26985 3490 6 n_55
rlabel m2contact 26961 3130 26961 3130 6 n_104
rlabel m2contact 26937 7042 26937 7042 6 n_153
rlabel m2contact 26937 4330 26937 4330 6 n_153
rlabel m2contact 26913 6514 26913 6514 6 n_354
rlabel m2contact 26889 4402 26889 4402 6 n_128
rlabel m2contact 26889 1858 26889 1858 6 n_128
rlabel m2contact 26865 3682 26865 3682 6 n_135
rlabel m2contact 26841 3562 26841 3562 6 n_320
rlabel m2contact 26817 3154 26817 3154 6 AluOR[0]
rlabel m2contact 26793 4666 26793 4666 6 n_30
rlabel m2contact 26769 4378 26769 4378 6 n_6
rlabel m2contact 26769 3370 26769 3370 6 RegWe
rlabel m2contact 26745 5458 26745 5458 6 n_12
rlabel m2contact 26721 4114 26721 4114 6 AluOR[1]
rlabel m2contact 26697 5146 26697 5146 6 n_185
rlabel m2contact 26673 6154 26673 6154 6 n_176
rlabel m2contact 26649 1954 26649 1954 6 n_193
rlabel m2contact 26649 2122 26649 2122 6 n_184
rlabel m2contact 26625 1882 26625 1882 6 n_161
rlabel m2contact 26625 3850 26625 3850 6 n_202
rlabel m2contact 26601 5002 26601 5002 6 stateSub[1]
rlabel m2contact 26577 4450 26577 4450 6 n_370
rlabel m2contact 26553 7042 26553 7042 6 n_153
rlabel m2contact 26553 7018 26553 7018 6 n_266
rlabel m2contact 26529 4402 26529 4402 6 n_128
rlabel m2contact 26529 1930 26529 1930 6 n_330
rlabel m2contact 26505 2554 26505 2554 6 n_336
rlabel m2contact 26505 3658 26505 3658 6 n_114
rlabel m2contact 26481 4402 26481 4402 6 n_299
rlabel m2contact 26481 3538 26481 3538 6 n_299
rlabel m2contact 26457 3586 26457 3586 6 n_28
rlabel m2contact 26433 3994 26433 3994 6 StatusRegEn
rlabel m2contact 26433 4018 26433 4018 6 n_42
rlabel m2contact 26409 3826 26409 3826 6 n_138
rlabel m2contact 26385 4426 26385 4426 6 n_60
rlabel m2contact 26385 2842 26385 2842 6 n_60
rlabel m2contact 26361 4210 26361 4210 6 n_308
rlabel m2contact 26337 4234 26337 4234 6 n_101
rlabel m2contact 26337 6034 26337 6034 6 n_305
rlabel m2contact 26313 4402 26313 4402 6 n_299
rlabel m2contact 26313 3874 26313 3874 6 stateSub[0]
rlabel m2contact 26289 2602 26289 2602 6 n_56
rlabel m2contact 26265 3202 26265 3202 6 n_378
rlabel m2contact 26241 5026 26241 5026 6 n_24
rlabel m2contact 26241 4090 26241 4090 6 n_309
rlabel m2contact 26217 5506 26217 5506 6 n_323
rlabel m2contact 26217 3514 26217 3514 6 n_215
rlabel m2contact 26193 4234 26193 4234 6 n_101
rlabel m2contact 26169 4402 26169 4402 6 n_224
rlabel m2contact 26169 3442 26169 3442 6 n_224
rlabel m2contact 26145 4426 26145 4426 6 n_60
rlabel m2contact 26145 3610 26145 3610 6 n_344
rlabel m2contact 26121 3226 26121 3226 6 OpcodeCondIn[1]
rlabel m2contact 26097 6754 26097 6754 6 n_11
rlabel m2contact 26097 2962 26097 2962 6 n_294
rlabel m2contact 26073 6154 26073 6154 6 n_176
rlabel m2contact 26073 4306 26073 4306 6 n_176
rlabel m2contact 26049 4402 26049 4402 6 n_224
rlabel m2contact 26049 4138 26049 4138 6 n_219
rlabel m2contact 26025 1882 26025 1882 6 n_161
rlabel m2contact 26001 4306 26001 4306 6 n_176
rlabel m2contact 26001 5962 26001 5962 6 n_231
rlabel m2contact 25977 2098 25977 2098 6 n_145
rlabel m2contact 25953 6994 25953 6994 6 n_63
rlabel m2contact 25929 3706 25929 3706 6 n_222
rlabel m2contact 25905 1738 25905 1738 6 n_25
rlabel m2contact 25869 5050 25869 5050 6 n_228
rlabel m2contact 25869 2674 25869 2674 6 n_228
rlabel m2contact 25857 6538 25857 6538 6 n_151
rlabel m2contact 25833 5050 25833 5050 6 n_228
rlabel m2contact 25833 5002 25833 5002 6 stateSub[1]
rlabel m2contact 25809 3778 25809 3778 6 n_180
rlabel m2contact 25785 6034 25785 6034 6 n_305
rlabel m2contact 25761 6082 25761 6082 6 n_269
rlabel m2contact 25737 2650 25737 2650 6 n_178
rlabel m2contact 25713 6706 25713 6706 6 n_237
rlabel m2contact 25665 3466 25665 3466 6 n_313
rlabel m2contact 25641 4258 25641 4258 6 n_86
rlabel m2contact 25617 4402 25617 4402 6 n_277
rlabel m2contact 25569 5530 25569 5530 6 n_136
rlabel m2contact 25521 3082 25521 3082 6 OpcodeCondIn[5]
rlabel m2contact 25497 3634 25497 3634 6 OpcodeCondIn[6]
rlabel m2contact 25449 5818 25449 5818 6 OpcodeCondIn[5]
rlabel m2contact 25449 3082 25449 3082 6 OpcodeCondIn[5]
rlabel m2contact 25425 3202 25425 3202 6 n_378
rlabel m2contact 25425 3250 25425 3250 6 n_66
rlabel m2contact 25401 5074 25401 5074 6 StatusReg[0]
rlabel m2contact 25401 1666 25401 1666 6 StatusReg[0]
rlabel m2contact 25377 3034 25377 3034 6 n_31
rlabel m2contact 25353 6562 25353 6562 6 n_337
rlabel m2contact 25353 4738 25353 4738 6 n_337
rlabel m2contact 25329 2506 25329 2506 6 n_246
rlabel m2contact 25305 6058 25305 6058 6 n_166
rlabel m2contact 25281 5050 25281 5050 6 n_108
rlabel m2contact 25281 2698 25281 2698 6 n_10
rlabel m2contact 25245 5002 25245 5002 6 stateSub[1]
rlabel m2contact 25245 4306 25245 4306 6 stateSub[1]
rlabel m2contact 25233 2314 25233 2314 6 n_230
rlabel m2contact 25233 5410 25233 5410 6 n_133
rlabel m2contact 25209 6370 25209 6370 6 n_96
rlabel m2contact 25209 2050 25209 2050 6 n_96
rlabel m2contact 25185 5818 25185 5818 6 OpcodeCondIn[5]
rlabel m2contact 25185 5794 25185 5794 6 n_342
rlabel m2contact 25161 1666 25161 1666 6 StatusReg[0]
rlabel m2contact 25161 1690 25161 1690 6 n_64
rlabel m2contact 25137 5890 25137 5890 6 n_335
rlabel m2contact 25113 4354 25113 4354 6 RwSel[1]
rlabel m2contact 25089 6562 25089 6562 6 n_337
rlabel m2contact 25089 6490 25089 6490 6 n_119
rlabel m2contact 25065 4306 25065 4306 6 stateSub[1]
rlabel m2contact 25065 4354 25065 4354 6 n_374
rlabel m2contact 25041 2050 25041 2050 6 n_96
rlabel m2contact 25041 2074 25041 2074 6 n_214
rlabel m2contact 24993 2266 24993 2266 6 n_23
rlabel m2contact 24969 3898 24969 3898 6 n_14
rlabel m2contact 24945 5002 24945 5002 6 stateSub[1]
rlabel m2contact 24897 5842 24897 5842 6 n_249
rlabel m2contact 24897 4906 24897 4906 6 state[0]
rlabel m2contact 24873 4306 24873 4306 6 OpcodeCondIn[7]
rlabel m2contact 24849 5962 24849 5962 6 n_231
rlabel m2contact 24849 5650 24849 5650 6 n_21
rlabel m2contact 24801 5602 24801 5602 6 n_37
rlabel m2contact 24753 2842 24753 2842 6 n_60
rlabel m2contact 24729 5074 24729 5074 6 StatusReg[0]
rlabel m2contact 24681 4378 24681 4378 6 n_6
rlabel m2contact 24657 3082 24657 3082 6 OpcodeCondIn[5]
rlabel m2contact 24633 4906 24633 4906 6 state[0]
rlabel m2contact 24585 4426 24585 4426 6 n_194
rlabel m2contact 24561 3994 24561 3994 6 nWait
rlabel m2contact 24537 1906 24537 1906 6 n_168
rlabel m2contact 24513 4618 24513 4618 6 n_212
rlabel m2contact 24489 1954 24489 1954 6 n_193
rlabel m2contact 24453 4378 24453 4378 6 n_85
rlabel m2contact 24453 2794 24453 2794 6 n_85
rlabel m2contact 24441 4690 24441 4690 6 n_284
rlabel m2contact 24417 6010 24417 6010 6 SysBus[3]
rlabel m2contact 24417 1666 24417 1666 6 SysBus[3]
rlabel m2contact 24393 2482 24393 2482 6 n_235
rlabel m2contact 24369 4426 24369 4426 6 n_194
rlabel m2contact 24369 3538 24369 3538 6 n_299
rlabel m2contact 24345 6178 24345 6178 6 n_287
rlabel m2contact 24321 6562 24321 6562 6 n_32
rlabel m2contact 24321 4642 24321 4642 6 n_221
rlabel m2contact 24297 2458 24297 2458 6 n_498
rlabel m2contact 24273 3922 24273 3922 6 StatusReg[3]
rlabel m2contact 24249 1690 24249 1690 6 n_64
rlabel m2contact 24225 4402 24225 4402 6 n_277
rlabel m2contact 24201 6730 24201 6730 6 n_276
rlabel m2contact 24201 5098 24201 5098 6 OpcodeCondIn[4]
rlabel m2contact 24177 3394 24177 3394 6 n_248
rlabel m2contact 24153 1594 24153 1594 6 n_199
rlabel m2contact 24129 5098 24129 5098 6 OpcodeCondIn[4]
rlabel m2contact 24105 4378 24105 4378 6 n_85
rlabel m2contact 24105 2938 24105 2938 6 n_159
rlabel m2contact 24081 5290 24081 5290 6 n_362
rlabel m2contact 24081 1882 24081 1882 6 n_161
rlabel m2contact 24057 4930 24057 4930 6 n_319
rlabel m2contact 24033 4378 24033 4378 6 n_383
rlabel m2contact 24009 2242 24009 2242 6 n_91
rlabel m2contact 23985 4906 23985 4906 6 state[0]
rlabel m2contact 23961 6802 23961 6802 6 n_84
rlabel m2contact 23937 6154 23937 6154 6 n_176
rlabel m2contact 23937 4186 23937 4186 6 n_176
rlabel m2contact 23913 1666 23913 1666 6 SysBus[3]
rlabel m2contact 23913 1762 23913 1762 6 n_139
rlabel m2contact 23889 1882 23889 1882 6 n_161
rlabel m2contact 23865 4186 23865 4186 6 n_176
rlabel m2contact 23865 5674 23865 5674 6 n_103
rlabel m2contact 23817 6850 23817 6850 6 n_328
rlabel m2contact 23817 4306 23817 4306 6 OpcodeCondIn[7]
rlabel m2contact 23793 4498 23793 4498 6 n_232
rlabel m2contact 23769 6586 23769 6586 6 n_329
rlabel m2contact 23745 2170 23745 2170 6 n_285
rlabel m2contact 23721 4978 23721 4978 6 n_247
rlabel m2contact 23697 4858 23697 4858 6 n_137
rlabel m2contact 23673 3826 23673 3826 6 n_138
rlabel m2contact 23649 4906 23649 4906 6 state[0]
rlabel m2contact 23625 6418 23625 6418 6 n_109
rlabel m2contact 23601 5722 23601 5722 6 n_188
rlabel m2contact 23601 1978 23601 1978 6 n_188
rlabel m2contact 23577 5722 23577 5722 6 n_188
rlabel m2contact 23577 5698 23577 5698 6 OpcodeCondIn[3]
rlabel m2contact 23553 3826 23553 3826 6 n_138
rlabel m2contact 23529 6802 23529 6802 6 n_84
rlabel m2contact 23505 4402 23505 4402 6 n_64
rlabel m2contact 23505 1690 23505 1690 6 n_64
rlabel m2contact 23481 4210 23481 4210 6 n_308
rlabel m2contact 23457 4546 23457 4546 6 n_350
rlabel m2contact 23457 5986 23457 5986 6 n_243
rlabel m2contact 23433 5434 23433 5434 6 n_190
rlabel m2contact 23433 4210 23433 4210 6 n_190
rlabel m2contact 23409 3082 23409 3082 6 OpcodeCondIn[5]
rlabel m2contact 23385 1954 23385 1954 6 n_193
rlabel m2contact 23361 4162 23361 4162 6 n_65
rlabel m2contact 23361 3970 23361 3970 6 n_227
rlabel m2contact 23337 4402 23337 4402 6 n_64
rlabel m2contact 23337 3874 23337 3874 6 stateSub[0]
rlabel m2contact 23313 4210 23313 4210 6 n_190
rlabel m2contact 23313 4474 23313 4474 6 n_154
rlabel m2contact 23289 6106 23289 6106 6 n_268
rlabel m2contact 23289 5386 23289 5386 6 n_268
rlabel m2contact 23265 3946 23265 3946 6 n_322
rlabel m2contact 23241 2722 23241 2722 6 n_17
rlabel m2contact 23217 6106 23217 6106 6 n_268
rlabel m2contact 23217 6034 23217 6034 6 n_305
rlabel m2contact 23193 5938 23193 5938 6 n_95
rlabel m2contact 23193 4426 23193 4426 6 n_241
rlabel m2contact 23169 5746 23169 5746 6 n_29
rlabel m2contact 23145 6106 23145 6106 6 n_74
rlabel m2contact 23145 4042 23145 4042 6 n_74
rlabel m2contact 23121 4330 23121 4330 6 n_153
rlabel m2contact 23121 6442 23121 6442 6 n_92
rlabel m2contact 23097 3778 23097 3778 6 n_180
rlabel m2contact 23073 6034 23073 6034 6 n_305
rlabel m2contact 23073 3874 23073 3874 6 stateSub[0]
rlabel m2contact 23049 6106 23049 6106 6 n_74
rlabel m2contact 23049 6034 23049 6034 6 n_305
rlabel m2contact 23001 3802 23001 3802 6 n_263
rlabel m2contact 22977 6010 22977 6010 6 SysBus[3]
rlabel m2contact 22977 5986 22977 5986 6 n_243
rlabel m2contact 22953 3754 22953 3754 6 n_239
rlabel m2contact 22953 4714 22953 4714 6 n_265
rlabel m2contact 22929 4330 22929 4330 6 stateSub[2]
rlabel m2contact 22929 3106 22929 3106 6 stateSub[2]
rlabel m2contact 22905 4186 22905 4186 6 n_298
rlabel m2contact 22881 3274 22881 3274 6 n_100
rlabel m2contact 22881 4498 22881 4498 6 n_232
rlabel m2contact 22857 1762 22857 1762 6 n_139
rlabel m2contact 22857 6250 22857 6250 6 n_296
rlabel m2contact 22833 6346 22833 6346 6 n_297
rlabel m2contact 22809 5266 22809 5266 6 n_88
rlabel m2contact 22785 6946 22785 6946 6 n_38
rlabel m2contact 22761 4330 22761 4330 6 stateSub[2]
rlabel m2contact 22761 3826 22761 3826 6 n_138
rlabel m2contact 22737 2266 22737 2266 6 n_23
rlabel m2contact 22713 4738 22713 4738 6 n_337
rlabel m2contact 22689 6202 22689 6202 6 n_71
rlabel m2contact 22665 5914 22665 5914 6 n_69
rlabel m2contact 22641 2026 22641 2026 6 n_279
rlabel m2contact 22641 4210 22641 4210 6 n_70
rlabel m2contact 22617 4330 22617 4330 6 state[1]
rlabel m2contact 22617 3298 22617 3298 6 state[1]
rlabel m2contact 22593 2434 22593 2434 6 n_261
rlabel m2contact 22569 4330 22569 4330 6 state[1]
rlabel m2contact 22569 3730 22569 3730 6 n_130
rlabel m2contact 22545 4042 22545 4042 6 n_74
rlabel m2contact 22545 2938 22545 2938 6 n_159
rlabel m2contact 22497 5578 22497 5578 6 IrWe
rlabel m2contact 22449 4042 22449 4042 6 n_74
rlabel m2contact 22449 6346 22449 6346 6 n_297
rlabel m2contact 22425 6082 22425 6082 6 n_269
rlabel m2contact 22425 4330 22425 4330 6 n_311
rlabel m2contact 22353 2146 22353 2146 6 n_352
rlabel m2contact 22353 2866 22353 2866 6 n_61
rlabel m2contact 22305 3946 22305 3946 6 n_322
rlabel m2contact 22305 4402 22305 4402 6 n_58
rlabel m2contact 22269 4594 22269 4594 6 n_126
rlabel m2contact 22269 3946 22269 3946 6 n_126
rlabel m2contact 22257 6130 22257 6130 6 n_59
rlabel m2contact 22233 3946 22233 3946 6 n_126
rlabel m2contact 22233 4402 22233 4402 6 n_58
rlabel m2contact 22209 6298 22209 6298 6 n_33
rlabel m2contact 22185 6562 22185 6562 6 n_32
rlabel m2contact 22185 2746 22185 2746 6 n_125
rlabel m2contact 22149 4522 22149 4522 6 n_181
rlabel m2contact 22149 3946 22149 3946 6 n_181
rlabel m2contact 22137 6466 22137 6466 6 n_182
rlabel m2contact 22113 4018 22113 4018 6 n_42
rlabel m2contact 22089 4522 22089 4522 6 n_181
rlabel m2contact 22089 4330 22089 4330 6 n_311
rlabel m2contact 22065 5242 22065 5242 6 n_346
rlabel m2contact 21993 3586 21993 3586 6 n_28
rlabel m2contact 21945 5074 21945 5074 6 StatusReg[0]
rlabel m2contact 21897 2194 21897 2194 6 n_15
rlabel m2contact 21873 4162 21873 4162 6 n_65
rlabel m2contact 21825 5122 21825 5122 6 ImmSel
rlabel m2contact 21801 6826 21801 6826 6 n_373
rlabel m2contact 21777 6874 21777 6874 6 n_361
rlabel m2contact 21753 4378 21753 4378 6 n_383
rlabel m2contact 21705 6826 21705 6826 6 n_373
rlabel m2contact 21681 5698 21681 5698 6 OpcodeCondIn[3]
rlabel m2contact 21657 5218 21657 5218 6 n_250
rlabel m2contact 21633 4810 21633 4810 6 n_236
rlabel m2contact 21633 2218 21633 2218 6 n_236
rlabel m2contact 21609 6010 21609 6010 6 n_195
rlabel m2contact 21585 5482 21585 5482 6 n_179
rlabel m2contact 21585 3010 21585 3010 6 n_179
rlabel m2contact 21573 6610 21573 6610 6 n_372
rlabel m2contact 21573 5818 21573 5818 6 n_372
rlabel m2contact 21561 4570 21561 4570 6 n_127
rlabel m2contact 21537 6610 21537 6610 6 n_372
rlabel m2contact 21537 6538 21537 6538 6 n_151
rlabel m2contact 21501 5170 21501 5170 6 n_34
rlabel m2contact 21501 4762 21501 4762 6 n_34
rlabel m2contact 21489 4258 21489 4258 6 n_86
rlabel m2contact 21465 3298 21465 3298 6 state[1]
rlabel m2contact 21441 2794 21441 2794 6 n_85
rlabel m2contact 21417 4786 21417 4786 6 n_178
rlabel m2contact 21417 2650 21417 2650 6 n_178
rlabel m2contact 21393 2962 21393 2962 6 n_294
rlabel m2contact 21369 2314 21369 2314 6 n_230
rlabel m2contact 21345 6082 21345 6082 6 n_269
rlabel m2contact 21345 5962 21345 5962 6 n_231
rlabel m2contact 21321 4498 21321 4498 6 n_232
rlabel m2contact 21297 3418 21297 3418 6 n_306
rlabel m2contact 21273 6034 21273 6034 6 n_305
rlabel m2contact 21273 2626 21273 2626 6 n_156
rlabel m2contact 21249 1954 21249 1954 6 n_193
rlabel m2contact 21249 6106 21249 6106 6 n_262
rlabel m2contact 21225 2938 21225 2938 6 n_159
rlabel m2contact 21201 4402 21201 4402 6 n_58
rlabel m2contact 21201 4522 21201 4522 6 n_77
rlabel m2contact 21177 2314 21177 2314 6 n_230
rlabel m2contact 21153 5170 21153 5170 6 n_34
rlabel m2contact 21153 4954 21153 4954 6 n_163
rlabel m2contact 21129 4858 21129 4858 6 n_137
rlabel m2contact 21105 4834 21105 4834 6 n_158
rlabel m2contact 21081 6730 21081 6730 6 n_276
rlabel m2contact 21057 1858 21057 1858 6 n_128
rlabel m2contact 21057 4882 21057 4882 6 n_157
rlabel m2contact 21033 2914 21033 2914 6 n_115
rlabel m2contact 21009 6634 21009 6634 6 n_187
rlabel m2contact 21009 4498 21009 4498 6 n_232
rlabel m2contact 20985 3106 20985 3106 6 stateSub[2]
rlabel m2contact 20961 4834 20961 4834 6 n_158
rlabel m2contact 20937 3706 20937 3706 6 n_222
rlabel m2contact 20913 2986 20913 2986 6 n_288
rlabel m2contact 20889 6178 20889 6178 6 n_287
rlabel m2contact 20889 5698 20889 5698 6 OpcodeCondIn[3]
rlabel m2contact 20865 1810 20865 1810 6 n_275
rlabel m2contact 20841 3346 20841 3346 6 n_82
rlabel m2contact 20817 4810 20817 4810 6 n_236
rlabel m2contact 20817 2386 20817 2386 6 n_81
rlabel m2contact 20793 1762 20793 1762 6 n_139
rlabel m2contact 20793 5914 20793 5914 6 n_69
rlabel m2contact 20769 5674 20769 5674 6 n_103
rlabel m2contact 20745 3010 20745 3010 6 n_179
rlabel m2contact 20745 3106 20745 3106 6 stateSub[2]
rlabel m2contact 20721 3058 20721 3058 6 OpcodeCondIn[2]
rlabel m2contact 20721 4210 20721 4210 6 n_70
rlabel m2contact 20697 5698 20697 5698 6 OpcodeCondIn[3]
rlabel m2contact 20673 3754 20673 3754 6 n_239
rlabel m2contact 20649 5194 20649 5194 6 PcSel[0]
rlabel m2contact 20625 4786 20625 4786 6 n_178
rlabel m2contact 20625 3586 20625 3586 6 n_357
rlabel m2contact 20601 3946 20601 3946 6 n_181
rlabel m2contact 20553 4762 20553 4762 6 n_34
rlabel m2contact 20529 6562 20529 6562 6 n_32
rlabel m2contact 20529 6418 20529 6418 6 n_109
rlabel m2contact 20505 5218 20505 5218 6 n_250
rlabel m2contact 20505 6298 20505 6298 6 n_33
rlabel m2contact 20481 6922 20481 6922 6 n_1
rlabel m2contact 20481 2050 20481 2050 6 n_1
rlabel m2contact 20457 4786 20457 4786 6 n_236
rlabel m2contact 20457 2218 20457 2218 6 n_236
rlabel m2contact 20433 6922 20433 6922 6 n_1
rlabel m2contact 20433 6898 20433 6898 6 n_67
rlabel m2contact 20409 5986 20409 5986 6 n_243
rlabel m2contact 20409 3010 20409 3010 6 n_243
rlabel m2contact 20385 4258 20385 4258 6 nIRQ
rlabel m2contact 20361 4762 20361 4762 6 n_380
rlabel m2contact 20361 3202 20361 3202 6 n_380
rlabel m2contact 20337 6610 20337 6610 6 n_290
rlabel m2contact 20337 4834 20337 4834 6 n_367
rlabel m2contact 20313 4186 20313 4186 6 n_298
rlabel m2contact 20289 5170 20289 5170 6 n_172
rlabel m2contact 20265 4786 20265 4786 6 n_236
rlabel m2contact 20265 4186 20265 4186 6 n_22
rlabel m2contact 20241 5698 20241 5698 6 OpcodeCondIn[3]
rlabel m2contact 20217 3010 20217 3010 6 n_243
rlabel m2contact 20217 3178 20217 3178 6 Op2Sel[0]
rlabel m2contact 20193 5722 20193 5722 6 n_132
rlabel m2contact 20193 4162 20193 4162 6 n_132
rlabel m2contact 20169 4642 20169 4642 6 n_221
rlabel m2contact 20145 3322 20145 3322 6 n_349
rlabel m2contact 20121 2410 20121 2410 6 n_216
rlabel m2contact 20097 6370 20097 6370 6 n_96
rlabel m2contact 20073 2746 20073 2746 6 n_125
rlabel m2contact 20049 3730 20049 3730 6 n_130
rlabel m2contact 20025 3202 20025 3202 6 n_380
rlabel m2contact 20025 3826 20025 3826 6 n_138
rlabel m2contact 20001 3442 20001 3442 6 n_224
rlabel m2contact 19977 4546 19977 4546 6 n_350
rlabel m2contact 19953 3322 19953 3322 6 n_349
rlabel m2contact 19929 5242 19929 5242 6 n_346
rlabel m2contact 19929 5098 19929 5098 6 OpcodeCondIn[4]
rlabel m2contact 19905 5674 19905 5674 6 n_103
rlabel m2contact 19881 6778 19881 6778 6 n_334
rlabel m2contact 19857 4162 19857 4162 6 n_132
rlabel m2contact 19857 4642 19857 4642 6 StatusReg[2]
rlabel m2contact 19833 5890 19833 5890 6 n_335
rlabel m2contact 19833 4306 19833 4306 6 OpcodeCondIn[7]
rlabel m2contact 19809 2338 19809 2338 6 n_87
rlabel m2contact 19785 4546 19785 4546 6 n_332
rlabel m2contact 19737 6442 19737 6442 6 n_92
rlabel m2contact 19713 4786 19713 4786 6 n_307
rlabel m2contact 19665 4810 19665 4810 6 n_387
rlabel m2contact 19617 4738 19617 4738 6 n_337
rlabel m2contact 19593 1834 19593 1834 6 n_377
rlabel m2contact 19521 4738 19521 4738 6 n_94
rlabel m2contact 19473 2386 19473 2386 6 n_81
rlabel m2contact 19425 2002 19425 2002 6 Flags[0]
rlabel m2contact 19377 2530 19377 2530 6 n_200
rlabel m2contact 19353 6394 19353 6394 6 n_331
rlabel m2contact 19353 3442 19353 3442 6 n_331
rlabel m2contact 19329 3082 19329 3082 6 OpcodeCondIn[5]
rlabel m2contact 19305 1594 19305 1594 6 n_199
rlabel m2contact 19281 5410 19281 5410 6 n_133
rlabel m2contact 19281 3202 19281 3202 6 n_133
rlabel m2contact 19257 2050 19257 2050 6 n_1
rlabel m2contact 19257 2290 19257 2290 6 n_218
rlabel m2contact 19233 3706 19233 3706 6 n_222
rlabel m2contact 19209 4594 19209 4594 6 n_126
rlabel m2contact 19185 6034 19185 6034 6 n_305
rlabel m2contact 19161 4594 19161 4594 6 n_165
rlabel m2contact 19161 2578 19161 2578 6 n_165
rlabel m2contact 19137 4162 19137 4162 6 n_280
rlabel m2contact 19113 6346 19113 6346 6 n_297
rlabel m2contact 19089 6250 19089 6250 6 n_296
rlabel m2contact 19089 3058 19089 3058 6 OpcodeCondIn[2]
rlabel m2contact 19065 2842 19065 2842 6 n_60
rlabel m2contact 19041 5242 19041 5242 6 n_346
rlabel m2contact 19017 3442 19017 3442 6 n_331
rlabel m2contact 19017 6178 19017 6178 6 n_287
rlabel m2contact 18993 2002 18993 2002 6 Flags[0]
rlabel m2contact 18993 2050 18993 2050 6 n_282
rlabel m2contact 18969 6586 18969 6586 6 n_329
rlabel m2contact 18945 5218 18945 5218 6 n_250
rlabel m2contact 18921 3442 18921 3442 6 n_134
rlabel m2contact 18897 3202 18897 3202 6 n_133
rlabel m2contact 18897 4618 18897 4618 6 n_212
rlabel m2contact 18873 4594 18873 4594 6 n_165
rlabel m2contact 18873 2938 18873 2938 6 n_159
rlabel m2contact 18837 5674 18837 5674 6 n_103
rlabel m2contact 18837 3202 18837 3202 6 n_103
rlabel m2contact 18825 3130 18825 3130 6 n_104
rlabel m2contact 18825 6178 18825 6178 6 n_287
rlabel m2contact 18801 5650 18801 5650 6 n_21
rlabel m2contact 18777 3202 18777 3202 6 n_103
rlabel m2contact 18777 3826 18777 3826 6 n_138
rlabel m2contact 18753 3250 18753 3250 6 n_66
rlabel m2contact 18729 6682 18729 6682 6 n_317
rlabel m2contact 18729 6322 18729 6322 6 n_317
rlabel m2contact 18705 6682 18705 6682 6 n_317
rlabel m2contact 18705 6658 18705 6658 6 n_47
rlabel m2contact 18681 3298 18681 3298 6 state[1]
rlabel m2contact 18657 3010 18657 3010 6 n_46
rlabel m2contact 18633 4594 18633 4594 6 n_52
rlabel m2contact 18633 2770 18633 2770 6 n_52
rlabel m2contact 18609 3322 18609 3322 6 n_349
rlabel m2contact 18585 5650 18585 5650 6 n_21
rlabel m2contact 18585 3058 18585 3058 6 OpcodeCondIn[2]
rlabel m2contact 18561 3130 18561 3130 6 OpcodeCondIn[0]
rlabel m2contact 18537 5170 18537 5170 6 n_172
rlabel m2contact 18513 6154 18513 6154 6 n_176
rlabel m2contact 18489 4594 18489 4594 6 n_52
rlabel m2contact 18489 3322 18489 3322 6 n_349
rlabel m2contact 18465 2986 18465 2986 6 n_288
rlabel m2contact 18465 3106 18465 3106 6 stateSub[2]
rlabel m2contact 18441 3874 18441 3874 6 stateSub[0]
rlabel m2contact 18417 4762 18417 4762 6 n_380
rlabel m2contact 18393 2362 18393 2362 6 n_49
rlabel m2contact 18369 1882 18369 1882 6 n_161
rlabel m2contact 18369 2938 18369 2938 6 n_159
rlabel m2contact 18321 3634 18321 3634 6 OpcodeCondIn[6]
rlabel m2contact 18273 2002 18273 2002 6 n_40
rlabel m2contact 18249 5410 18249 5410 6 n_133
rlabel m2contact 18225 2362 18225 2362 6 n_49
rlabel m2contact 18153 5098 18153 5098 6 OpcodeCondIn[4]
rlabel m2contact 18105 3082 18105 3082 6 OpcodeCondIn[5]
rlabel m2contact 18057 3562 18057 3562 6 n_320
rlabel m2contact 18009 5098 18009 5098 6 OpcodeCondIn[4]
rlabel m2contact 17985 4162 17985 4162 6 n_280
rlabel m2contact 17913 6922 17913 6922 6 LrSel
rlabel m2contact 17817 4450 17817 4450 6 n_370
rlabel m2contact 17793 3730 17793 3730 6 n_130
rlabel m2contact 17769 6610 17769 6610 6 n_290
rlabel m2contact 17769 3562 17769 3562 6 n_290
rlabel m2contact 17745 5170 17745 5170 6 n_170
rlabel m2contact 17721 5242 17721 5242 6 OpcodeCondIn[2]
rlabel m2contact 17721 3058 17721 3058 6 OpcodeCondIn[2]
rlabel m2contact 17697 4162 17697 4162 6 n_234
rlabel m2contact 17673 3106 17673 3106 6 stateSub[2]
rlabel m2contact 17649 5218 17649 5218 6 n_175
rlabel m2contact 17625 6466 17625 6466 6 n_182
rlabel m2contact 17625 6322 17625 6322 6 n_317
rlabel m2contact 17601 6730 17601 6730 6 n_276
rlabel m2contact 17577 5314 17577 5314 6 n_93
rlabel m2contact 17553 2818 17553 2818 6 n_291
rlabel m2contact 17553 3322 17553 3322 6 n_349
rlabel m2contact 17529 6442 17529 6442 6 n_92
rlabel m2contact 17529 6322 17529 6322 6 n_317
rlabel m2contact 17505 4882 17505 4882 6 n_157
rlabel m2contact 17481 3562 17481 3562 6 n_290
rlabel m2contact 17481 5770 17481 5770 6 n_169
rlabel m2contact 17457 5242 17457 5242 6 OpcodeCondIn[2]
rlabel m2contact 17457 4978 17457 4978 6 n_247
rlabel m2contact 17433 1906 17433 1906 6 n_168
rlabel m2contact 17409 5434 17409 5434 6 n_190
rlabel m2contact 17337 4594 17337 4594 6 n_255
rlabel m2contact 17313 5626 17313 5626 6 IRQ2
rlabel m2contact 17289 5242 17289 5242 6 n_226
rlabel m2contact 17241 3202 17241 3202 6 n_206
rlabel m2contact 17217 6562 17217 6562 6 n_43
rlabel m2contact 17193 5362 17193 5362 6 n_207
rlabel m2contact 17145 4450 17145 4450 6 n_80
rlabel m2contact 17121 2914 17121 2914 6 n_115
rlabel m2contact 17097 4666 17097 4666 6 n_30
rlabel m2contact 17073 6970 17073 6970 6 n_201
rlabel m2contact 17073 2986 17073 2986 6 n_201
rlabel m2contact 17049 4666 17049 4666 6 n_301
rlabel m2contact 17025 3082 17025 3082 6 OpcodeCondIn[5]
rlabel m2contact 17001 5866 17001 5866 6 n_260
rlabel m2contact 16977 7042 16977 7042 6 n_20
rlabel m2contact 16977 3562 16977 3562 6 n_20
rlabel m2contact 16953 6226 16953 6226 6 n_68
rlabel m2contact 16929 5530 16929 5530 6 n_136
rlabel m2contact 16905 2650 16905 2650 6 n_178
rlabel m2contact 16869 6082 16869 6082 6 n_257
rlabel m2contact 16869 3250 16869 3250 6 n_257
rlabel m2contact 16857 6442 16857 6442 6 n_7
rlabel m2contact 16833 3130 16833 3130 6 OpcodeCondIn[0]
rlabel m2contact 16809 3226 16809 3226 6 OpcodeCondIn[1]
rlabel m2contact 16773 5338 16773 5338 6 n_58
rlabel m2contact 16773 4402 16773 4402 6 n_58
rlabel m2contact 16761 5458 16761 5458 6 n_12
rlabel m2contact 16737 2986 16737 2986 6 n_201
rlabel m2contact 16737 3634 16737 3634 6 OpcodeCondIn[6]
rlabel m2contact 16713 3250 16713 3250 6 n_257
rlabel m2contact 16713 3874 16713 3874 6 stateSub[0]
rlabel m2contact 16689 5698 16689 5698 6 OpcodeCondIn[3]
rlabel m2contact 16665 3490 16665 3490 6 n_55
rlabel m2contact 16641 3250 16641 3250 6 n_44
rlabel m2contact 16617 3874 16617 3874 6 stateSub[0]
rlabel m2contact 16593 3562 16593 3562 6 n_20
rlabel m2contact 16593 3634 16593 3634 6 OpcodeCondIn[6]
rlabel m2contact 16569 3826 16569 3826 6 n_138
rlabel m2contact 16545 6466 16545 6466 6 n_118
rlabel m2contact 16521 5338 16521 5338 6 n_58
rlabel m2contact 16521 5002 16521 5002 6 stateSub[1]
rlabel m2contact 16497 5362 16497 5362 6 n_207
rlabel m2contact 16497 1666 16497 1666 6 n_207
rlabel m2contact 16473 3226 16473 3226 6 OpcodeCondIn[1]
rlabel m2contact 16449 6754 16449 6754 6 n_11
rlabel m2contact 16449 3490 16449 3490 6 n_35
rlabel m2contact 16425 1954 16425 1954 6 n_193
rlabel m2contact 16401 3562 16401 3562 6 n_121
rlabel m2contact 16401 2842 16401 2842 6 n_60
rlabel m2contact 16377 5458 16377 5458 6 n_62
rlabel m2contact 16353 5674 16353 5674 6 n_103
rlabel m2contact 16329 1666 16329 1666 6 n_207
rlabel m2contact 16329 5002 16329 5002 6 stateSub[1]
rlabel m2contact 16305 5554 16305 5554 6 n_89
rlabel m2contact 16305 2986 16305 2986 6 n_89
rlabel m2contact 16281 5050 16281 5050 6 n_108
rlabel m2contact 16281 4762 16281 4762 6 n_380
rlabel m2contact 16257 4498 16257 4498 6 n_232
rlabel m2contact 16233 2986 16233 2986 6 n_89
rlabel m2contact 16233 3514 16233 3514 6 n_215
rlabel m2contact 16209 3058 16209 3058 6 OpcodeCondIn[2]
rlabel m2contact 16185 2986 16185 2986 6 AluWe
rlabel m2contact 16185 2098 16185 2098 6 n_145
rlabel m2contact 16137 5338 16137 5338 6 n_369
rlabel m2contact 16113 3802 16113 3802 6 n_263
rlabel m2contact 16041 3106 16041 3106 6 stateSub[2]
rlabel m2contact 16017 1738 16017 1738 6 n_25
rlabel m2contact 15993 3802 15993 3802 6 n_8
rlabel m2contact 15993 3826 15993 3826 6 n_138
rlabel m2contact 15969 5026 15969 5026 6 n_24
rlabel m2contact 15897 3130 15897 3130 6 OpcodeCondIn[0]
rlabel m2contact 15873 3250 15873 3250 6 n_44
rlabel m2contact 15777 3706 15777 3706 6 n_222
rlabel m2contact 15753 5674 15753 5674 6 n_103
rlabel m2contact 15657 1762 15657 1762 6 n_139
rlabel m2contact 15633 3562 15633 3562 6 n_121
rlabel m2contact 15633 6682 15633 6682 6 n_293
rlabel m2contact 15585 2410 15585 2410 6 n_216
rlabel m2contact 15561 2746 15561 2746 6 n_125
rlabel m2contact 15537 5650 15537 5650 6 n_21
rlabel m2contact 15537 3562 15537 3562 6 n_21
rlabel m2contact 15513 2746 15513 2746 6 n_198
rlabel m2contact 15489 2722 15489 2722 6 n_17
rlabel m2contact 15489 4618 15489 4618 6 n_212
rlabel m2contact 15465 3562 15465 3562 6 n_21
rlabel m2contact 15465 3826 15465 3826 6 n_138
rlabel m2contact 15441 3874 15441 3874 6 stateSub[0]
rlabel m2contact 15417 3562 15417 3562 6 PcSel[1]
rlabel m2contact 15393 2986 15393 2986 6 AluWe
rlabel m2contact 15345 4378 15345 4378 6 n_383
rlabel m2contact 15321 4354 15321 4354 6 n_374
rlabel m2contact 15273 3922 15273 3922 6 StatusReg[3]
rlabel m2contact 15249 5050 15249 5050 6 n_240
rlabel m2contact 15225 3082 15225 3082 6 OpcodeCondIn[5]
rlabel m2contact 15225 6274 15225 6274 6 n_499
rlabel m2contact 15201 3754 15201 3754 6 n_239
rlabel m2contact 15105 4738 15105 4738 6 n_94
rlabel m2contact 14985 4066 14985 4066 6 n_141
rlabel m2contact 14889 3754 14889 3754 6 n_209
rlabel m2contact 14865 5338 14865 5338 6 n_369
rlabel m2contact 14841 6154 14841 6154 6 n_176
rlabel m2contact 14817 2578 14817 2578 6 n_165
rlabel m2contact 14745 6898 14745 6898 6 n_67
rlabel m2contact 14745 6730 14745 6730 6 n_276
rlabel m2contact 14721 6034 14721 6034 6 n_305
rlabel m2contact 14697 2266 14697 2266 6 n_23
rlabel m2contact 14697 2602 14697 2602 6 n_56
rlabel m2contact 14649 4330 14649 4330 6 n_311
rlabel m2contact 14625 5290 14625 5290 6 n_362
rlabel m2contact 14601 3322 14601 3322 6 n_349
rlabel m2contact 14577 2674 14577 2674 6 n_228
rlabel m2contact 14577 5338 14577 5338 6 n_356
rlabel m2contact 14553 5290 14553 5290 6 n_267
rlabel m2contact 14553 2986 14553 2986 6 n_267
rlabel m2contact 14529 5818 14529 5818 6 n_372
rlabel m2contact 14529 3082 14529 3082 6 n_286
rlabel m2contact 14505 5290 14505 5290 6 n_267
rlabel m2contact 14505 5098 14505 5098 6 OpcodeCondIn[4]
rlabel m2contact 14481 6394 14481 6394 6 n_331
rlabel m2contact 14481 5818 14481 5818 6 n_186
rlabel m2contact 14457 5794 14457 5794 6 n_342
rlabel m2contact 14457 5530 14457 5530 6 n_136
rlabel m2contact 14433 5290 14433 5290 6 n_145
rlabel m2contact 14433 2098 14433 2098 6 n_145
rlabel m2contact 14409 5194 14409 5194 6 PcSel[0]
rlabel m2contact 14373 6394 14373 6394 6 n_271
rlabel m2contact 14373 2722 14373 2722 6 n_271
rlabel m2contact 14361 2362 14361 2362 6 n_49
rlabel m2contact 14337 4930 14337 4930 6 n_319
rlabel m2contact 14337 3826 14337 3826 6 n_138
rlabel m2contact 14313 5794 14313 5794 6 IntStatus
rlabel m2contact 14313 1666 14313 1666 6 IntStatus
rlabel m2contact 14289 6586 14289 6586 6 n_329
rlabel m2contact 14289 4930 14289 4930 6 n_99
rlabel m2contact 14265 5986 14265 5986 6 n_243
rlabel m2contact 14241 5290 14241 5290 6 n_145
rlabel m2contact 14241 5194 14241 5194 6 n_54
rlabel m2contact 14217 6586 14217 6586 6 n_329
rlabel m2contact 14217 4066 14217 4066 6 n_329
rlabel m2contact 14193 2314 14193 2314 6 n_230
rlabel m2contact 14169 6418 14169 6418 6 n_109
rlabel m2contact 14145 2866 14145 2866 6 n_61
rlabel m2contact 14121 4786 14121 4786 6 n_307
rlabel m2contact 14121 2842 14121 2842 6 n_60
rlabel m2contact 14097 7066 14097 7066 6 n_219
rlabel m2contact 14097 4138 14097 4138 6 n_219
rlabel m2contact 14073 2722 14073 2722 6 n_271
rlabel m2contact 14073 3322 14073 3322 6 n_349
rlabel m2contact 14049 2266 14049 2266 6 n_259
rlabel m2contact 14025 1738 14025 1738 4 n_90
rlabel m2contact 14001 4786 14001 4786 4 n_213
rlabel m2contact 14001 4858 14001 4858 4 n_137
rlabel m2contact 13977 6706 13977 6706 4 n_237
rlabel m2contact 13977 1618 13977 1618 4 n_237
rlabel m2contact 13953 5626 13953 5626 4 IRQ2
rlabel m2contact 13953 5290 13953 5290 4 n_256
rlabel m2contact 13929 5794 13929 5794 4 IntStatus
rlabel m2contact 13929 5698 13929 5698 4 OpcodeCondIn[3]
rlabel m2contact 13905 3754 13905 3754 4 n_209
rlabel m2contact 13881 2314 13881 2314 4 n_230
rlabel m2contact 13881 5794 13881 5794 4 n_144
rlabel m2contact 13857 5698 13857 5698 4 OpcodeCondIn[3]
rlabel m2contact 13833 2938 13833 2938 4 n_159
rlabel m2contact 13809 6898 13809 6898 4 n_193
rlabel m2contact 13809 1954 13809 1954 4 n_193
rlabel m2contact 13785 5626 13785 5626 4 n_19
rlabel m2contact 13761 1762 13761 1762 4 n_39
rlabel m2contact 13761 3130 13761 3130 4 OpcodeCondIn[0]
rlabel m2contact 13737 5074 13737 5074 4 StatusReg[0]
rlabel m2contact 13713 3226 13713 3226 4 OpcodeCondIn[1]
rlabel m2contact 13689 5434 13689 5434 4 n_190
rlabel m2contact 13665 4786 13665 4786 4 n_213
rlabel m2contact 13665 3778 13665 3778 4 n_180
rlabel m2contact 13641 6418 13641 6418 4 n_109
rlabel m2contact 13641 1642 13641 1642 4 n_109
rlabel m2contact 13617 4066 13617 4066 4 n_329
rlabel m2contact 13617 4618 13617 4618 4 n_212
rlabel m2contact 13593 5962 13593 5962 4 n_231
rlabel m2contact 13569 4162 13569 4162 4 n_234
rlabel m2contact 13545 1594 13545 1594 4 n_199
rlabel m2contact 13545 2050 13545 2050 4 n_282
rlabel m2contact 13521 4786 13521 4786 4 n_304
rlabel m2contact 13497 2722 13497 2722 4 n_273
rlabel m2contact 13473 7066 13473 7066 4 n_219
rlabel m2contact 13473 5074 13473 5074 4 n_245
rlabel m2contact 13449 1690 13449 1690 4 n_64
rlabel m2contact 13425 1618 13425 1618 4 n_237
rlabel m2contact 13425 4066 13425 4066 4 n_281
rlabel m2contact 13401 4162 13401 4162 4 n_210
rlabel m2contact 13377 6250 13377 6250 4 n_296
rlabel m2contact 13377 4786 13377 4786 4 n_304
rlabel m2contact 13353 5986 13353 5986 4 n_243
rlabel m2contact 13329 7042 13329 7042 4 n_20
rlabel m2contact 13329 2938 13329 2938 4 n_159
rlabel m2contact 13305 6898 13305 6898 4 n_193
rlabel m2contact 13305 2650 13305 2650 4 n_178
rlabel m2contact 13281 3826 13281 3826 4 n_138
rlabel m2contact 13257 1882 13257 1882 4 n_161
rlabel m2contact 13233 4498 13233 4498 4 n_232
rlabel m2contact 13209 1642 13209 1642 4 n_109
rlabel m2contact 13209 3970 13209 3970 4 n_227
rlabel m2contact 13161 3682 13161 3682 4 n_135
rlabel m2contact 13161 3850 13161 3850 4 n_202
rlabel m2contact 13137 6418 13137 6418 4 n_109
rlabel m2contact 13113 4930 13113 4930 4 n_99
rlabel m2contact 13089 2938 13089 2938 4 n_159
rlabel m2contact 13017 1954 13017 1954 4 n_193
rlabel m2contact 12969 3682 12969 3682 4 MemEn
rlabel m2contact 12969 3058 12969 3058 4 OpcodeCondIn[2]
rlabel m2contact 12921 6370 12921 6370 4 n_96
rlabel m2contact 12921 4570 12921 4570 4 n_127
rlabel m2contact 12897 6178 12897 6178 4 n_287
rlabel m2contact 12897 1882 12897 1882 4 n_161
rlabel m2contact 12873 6418 12873 6418 4 n_27
rlabel m2contact 12873 3730 12873 3730 4 n_130
rlabel m2contact 12825 3682 12825 3682 4 MemEn
rlabel m2contact 12825 6898 12825 6898 4 n_211
rlabel m2contact 12801 4162 12801 4162 4 n_210
rlabel m2contact 12777 5146 12777 5146 4 n_185
rlabel m2contact 12777 5962 12777 5962 4 n_231
rlabel m2contact 12753 3682 12753 3682 4 n_312
rlabel m2contact 12729 6370 12729 6370 4 n_340
rlabel m2contact 12705 5146 12705 5146 4 n_252
rlabel m2contact 12681 1954 12681 1954 4 n_193
rlabel m2contact 12681 6178 12681 6178 4 n_177
rlabel m2contact 12657 4138 12657 4138 4 n_219
rlabel m2contact 12657 5290 12657 5290 4 n_256
rlabel m2contact 12609 4138 12609 4138 4 SysBus[0]
rlabel m2contact 12609 5290 12609 5290 4 n_278
rlabel m2contact 12585 3970 12585 3970 4 n_227
rlabel m2contact 12561 2506 12561 2506 4 n_246
rlabel m2contact 12513 2506 12513 2506 4 LrWe
rlabel m2contact 12465 1666 12465 1666 4 IntStatus
rlabel m2contact 12465 1762 12465 1762 4 n_39
rlabel m2contact 12417 1882 12417 1882 4 n_161
rlabel m2contact 12393 3010 12393 3010 4 n_46
rlabel m2contact 12345 2794 12345 2794 4 n_85
rlabel m2contact 12321 6730 12321 6730 4 n_276
rlabel m2contact 12297 4042 12297 4042 4 n_74
rlabel m2contact 12249 2986 12249 2986 4 n_267
rlabel m2contact 12225 4138 12225 4138 4 SysBus[0]
rlabel m2contact 12201 4714 12201 4714 4 n_265
rlabel m2contact 12153 4138 12153 4138 4 n_174
rlabel m2contact 12105 5530 12105 5530 4 n_136
rlabel m2contact 12081 2938 12081 2938 4 n_159
rlabel m2contact 12033 1882 12033 1882 4 WdSel
rlabel m2contact 11985 7018 11985 7018 4 n_266
rlabel m2contact 11961 1762 11961 1762 4 SysBus[1]
rlabel m2contact 11937 4714 11937 4714 4 n_265
rlabel m2contact 11889 2986 11889 2986 4 n_167
rlabel m2contact 11865 4162 11865 4162 4 n_210
rlabel m2contact 11841 1882 11841 1882 4 WdSel
rlabel m2contact 11841 1906 11841 1906 4 n_168
rlabel m2contact 11817 7018 11817 7018 4 n_122
rlabel m2contact 11817 2794 11817 2794 4 n_122
rlabel m2contact 11793 7018 11793 7018 4 n_122
rlabel m2contact 11793 5482 11793 5482 4 n_179
rlabel m2contact 11769 6994 11769 6994 4 n_63
rlabel m2contact 11769 6010 11769 6010 4 n_195
rlabel m2contact 11745 4450 11745 4450 4 n_80
rlabel m2contact 11721 6994 11721 6994 4 n_228
rlabel m2contact 11721 2674 11721 2674 4 n_228
rlabel m2contact 11697 4450 11697 4450 4 n_292
rlabel m2contact 11673 6994 11673 6994 4 n_228
rlabel m2contact 11673 5170 11673 5170 4 n_170
rlabel m2contact 11649 1882 11649 1882 4 n_253
rlabel m2contact 11625 3850 11625 3850 4 n_202
rlabel m2contact 11601 2890 11601 2890 4 Rs1Sel[0]
rlabel m2contact 11577 6970 11577 6970 4 n_201
rlabel m2contact 11577 6322 11577 6322 4 n_317
rlabel m2contact 11553 2890 11553 2890 4 n_149
rlabel m2contact 11529 4906 11529 4906 4 state[0]
rlabel m2contact 11505 6946 11505 6946 4 n_38
rlabel m2contact 11481 6922 11481 6922 4 LrSel
rlabel m2contact 11481 5098 11481 5098 4 OpcodeCondIn[4]
rlabel m2contact 11481 1666 11481 1666 4 OpcodeCondIn[4]
rlabel m2contact 11457 5194 11457 5194 4 n_54
rlabel m2contact 11433 1666 11433 1666 4 OpcodeCondIn[4]
rlabel m2contact 11433 4354 11433 4354 4 n_374
rlabel m2contact 11409 3706 11409 3706 4 n_222
rlabel m2contact 11385 4834 11385 4834 4 n_367
rlabel m2contact 11361 6898 11361 6898 4 n_211
rlabel m2contact 11361 4018 11361 4018 4 n_42
rlabel m2contact 11337 5986 11337 5986 4 n_243
rlabel m2contact 11313 1690 11313 1690 4 n_64
rlabel m2contact 11313 3010 11313 3010 4 n_46
rlabel m2contact 11265 5650 11265 5650 4 n_21
rlabel m2contact 11241 1714 11241 1714 4 Flags[3]
rlabel m2contact 11241 3826 11241 3826 4 n_138
rlabel m2contact 11217 6586 11217 6586 4 n_329
rlabel m2contact 11193 1738 11193 1738 4 n_90
rlabel m2contact 11169 1762 11169 1762 4 SysBus[1]
rlabel m2contact 11169 6898 11169 6898 4 n_261
rlabel m2contact 11169 2434 11169 2434 4 n_261
rlabel m2contact 11145 5002 11145 5002 4 stateSub[1]
rlabel m2contact 11121 6898 11121 6898 4 n_261
rlabel m2contact 11121 3586 11121 3586 4 n_357
rlabel m2contact 11097 6730 11097 6730 4 n_276
rlabel m2contact 11037 6898 11037 6898 4 n_357
rlabel m2contact 11037 3586 11037 3586 4 n_357
rlabel m2contact 11025 1810 11025 1810 4 n_275
rlabel m2contact 11001 6898 11001 6898 4 n_357
rlabel m2contact 11001 3706 11001 3706 4 n_222
rlabel m2contact 10977 2722 10977 2722 4 n_273
rlabel m2contact 10953 6082 10953 6082 4 n_257
rlabel m2contact 10953 1810 10953 1810 4 n_257
rlabel m2contact 10929 1786 10929 1786 4 RwSel[0]
rlabel m2contact 10929 5962 10929 5962 4 n_231
rlabel m2contact 10905 5002 10905 5002 4 stateSub[1]
rlabel m2contact 10881 5794 10881 5794 4 n_144
rlabel m2contact 10857 6322 10857 6322 4 n_317
rlabel m2contact 10833 1810 10833 1810 4 n_257
rlabel m2contact 10833 2578 10833 2578 4 n_165
rlabel m2contact 10785 6730 10785 6730 4 n_276
rlabel m2contact 10761 3850 10761 3850 4 n_202
rlabel m2contact 10737 2410 10737 2410 4 n_216
rlabel m2contact 10713 5122 10713 5122 4 ImmSel
rlabel m2contact 10677 5122 10677 5122 4 n_188
rlabel m2contact 10677 1978 10677 1978 4 n_188
rlabel m2contact 10665 6322 10665 6322 4 n_107
rlabel m2contact 10641 4042 10641 4042 4 n_74
rlabel m2contact 10617 5122 10617 5122 4 n_188
rlabel m2contact 10617 3994 10617 3994 4 nWait
rlabel m2contact 10545 6874 10545 6874 4 n_361
rlabel m2contact 10545 5434 10545 5434 4 n_190
rlabel m2contact 10497 1858 10497 1858 4 n_128
rlabel m2contact 10497 5122 10497 5122 4 n_351
rlabel m2contact 10473 4042 10473 4042 4 n_184
rlabel m2contact 10473 2122 10473 2122 4 n_184
rlabel m2contact 10449 2482 10449 2482 4 n_235
rlabel m2contact 10425 4042 10425 4042 4 n_184
rlabel m2contact 10425 3634 10425 3634 4 OpcodeCondIn[6]
rlabel m2contact 10401 5962 10401 5962 4 n_231
rlabel m2contact 10377 5554 10377 5554 4 n_89
rlabel m2contact 10353 6154 10353 6154 4 n_176
rlabel m2contact 10353 4042 10353 4042 4 n_176
rlabel m2contact 10329 2890 10329 2890 4 n_149
rlabel m2contact 10329 5938 10329 5938 4 n_95
rlabel m2contact 10305 4042 10305 4042 4 n_176
rlabel m2contact 10305 6034 10305 6034 4 n_305
rlabel m2contact 10281 4738 10281 4738 4 n_94
rlabel m2contact 10233 5170 10233 5170 4 n_170
rlabel m2contact 10209 4042 10209 4042 4 n_72
rlabel m2contact 10185 2914 10185 2914 4 n_115
rlabel m2contact 10161 2434 10161 2434 4 n_261
rlabel m2contact 10137 1906 10137 1906 4 n_168
rlabel m2contact 10113 2482 10113 2482 4 n_326
rlabel m2contact 10089 2890 10089 2890 4 n_208
rlabel m2contact 10089 5002 10089 5002 4 stateSub[1]
rlabel m2contact 10065 3418 10065 3418 4 n_306
rlabel m2contact 10065 3970 10065 3970 4 n_227
rlabel m2contact 10041 5986 10041 5986 4 n_243
rlabel m2contact 10041 1858 10041 1858 4 n_243
rlabel m2contact 10017 5938 10017 5938 4 n_371
rlabel m2contact 9993 3922 9993 3922 4 StatusReg[3]
rlabel m2contact 9993 4738 9993 4738 4 n_264
rlabel m2contact 9969 6850 9969 6850 4 n_328
rlabel m2contact 9969 5890 9969 5890 4 n_335
rlabel m2contact 9945 6778 9945 6778 4 n_334
rlabel m2contact 9921 6850 9921 6850 4 n_165
rlabel m2contact 9921 2578 9921 2578 4 n_165
rlabel m2contact 9897 3298 9897 3298 4 state[1]
rlabel m2contact 9873 6754 9873 6754 4 n_11
rlabel m2contact 9873 4906 9873 4906 4 state[0]
rlabel m2contact 9849 6154 9849 6154 4 n_176
rlabel m2contact 9849 3922 9849 3922 4 n_176
rlabel m2contact 9825 1834 9825 1834 4 n_377
rlabel m2contact 9825 3130 9825 3130 4 OpcodeCondIn[0]
rlabel m2contact 9801 6778 9801 6778 4 n_349
rlabel m2contact 9801 3322 9801 3322 4 n_349
rlabel m2contact 9777 2530 9777 2530 4 n_200
rlabel m2contact 9777 5578 9777 5578 4 IrWe
rlabel m2contact 9753 3418 9753 3418 4 n_355
rlabel m2contact 9729 2938 9729 2938 4 n_159
rlabel m2contact 9705 6754 9705 6754 4 n_229
rlabel m2contact 9705 2530 9705 2530 4 n_229
rlabel m2contact 9681 1858 9681 1858 4 n_243
rlabel m2contact 9681 3106 9681 3106 4 stateSub[2]
rlabel m2contact 9657 6850 9657 6850 4 n_165
rlabel m2contact 9657 5362 9657 5362 4 n_207
rlabel m2contact 9633 5578 9633 5578 4 OpcodeCondIn[2]
rlabel m2contact 9633 3058 9633 3058 4 OpcodeCondIn[2]
rlabel m2contact 9609 4282 9609 4282 4 Rs1Sel[1]
rlabel m2contact 9585 6826 9585 6826 4 n_373
rlabel m2contact 9585 4474 9585 4474 4 n_154
rlabel m2contact 9561 1906 9561 1906 4 n_168
rlabel m2contact 9561 4354 9561 4354 4 n_374
rlabel m2contact 9537 3922 9537 3922 4 n_176
rlabel m2contact 9537 4282 9537 4282 4 n_324
rlabel m2contact 9513 6370 9513 6370 4 n_340
rlabel m2contact 9489 3922 9489 3922 4 nME
rlabel m2contact 9465 4114 9465 4114 4 AluOR[1]
rlabel m2contact 9465 2386 9465 2386 4 n_81
rlabel m2contact 9441 2026 9441 2026 4 n_279
rlabel m2contact 9417 4114 9417 4114 4 n_359
rlabel m2contact 9393 4834 9393 4834 4 n_367
rlabel m2contact 9369 1906 9369 1906 4 n_120
rlabel m2contact 9345 6802 9345 6802 4 n_84
rlabel m2contact 9345 4858 9345 4858 4 n_137
rlabel m2contact 9321 6778 9321 6778 4 n_349
rlabel m2contact 9321 3826 9321 3826 4 n_138
rlabel m2contact 9297 6730 9297 6730 4 n_276
rlabel m2contact 9273 6082 9273 6082 4 n_257
rlabel m2contact 9249 6754 9249 6754 4 n_229
rlabel m2contact 9249 3706 9249 3706 4 n_222
rlabel m2contact 9225 5578 9225 5578 4 OpcodeCondIn[2]
rlabel m2contact 9225 4906 9225 4906 4 state[0]
rlabel m2contact 9201 3970 9201 3970 4 n_227
rlabel m2contact 9177 2674 9177 2674 4 n_228
rlabel m2contact 9153 1882 9153 1882 4 n_253
rlabel m2contact 9153 4618 9153 4618 4 n_212
rlabel m2contact 9105 5242 9105 5242 4 n_226
rlabel m2contact 9105 5146 9105 5146 4 n_252
rlabel m2contact 9081 2002 9081 2002 4 n_40
rlabel m2contact 9057 5578 9057 5578 4 n_116
rlabel m2contact 9057 5242 9057 5242 4 n_112
rlabel m2contact 9033 5266 9033 5266 4 n_88
rlabel m2contact 9033 5002 9033 5002 4 stateSub[1]
rlabel m2contact 9009 5722 9009 5722 4 n_132
rlabel m2contact 8985 5266 8985 5266 4 n_302
rlabel m2contact 8985 2002 8985 2002 4 n_302
rlabel m2contact 8961 2002 8961 2002 4 n_302
rlabel m2contact 8961 4834 8961 4834 4 n_367
rlabel m2contact 8937 1978 8937 1978 4 n_188
rlabel m2contact 8937 5650 8937 5650 4 n_21
rlabel m2contact 8913 6730 8913 6730 4 n_276
rlabel m2contact 8913 5722 8913 5722 4 n_270
rlabel m2contact 8889 3106 8889 3106 4 stateSub[2]
rlabel m2contact 8865 3298 8865 3298 4 state[1]
rlabel m2contact 8841 2914 8841 2914 4 n_115
rlabel m2contact 8817 2002 8817 2002 4 n_160
rlabel m2contact 8793 4906 8793 4906 4 state[0]
rlabel m2contact 8793 4306 8793 4306 4 OpcodeCondIn[7]
rlabel m2contact 8769 1906 8769 1906 4 n_120
rlabel m2contact 8745 2602 8745 2602 4 n_56
rlabel m2contact 8721 6706 8721 6706 4 n_237
rlabel m2contact 8697 3826 8697 3826 4 n_138
rlabel m2contact 8673 4306 8673 4306 4 OpcodeCondIn[7]
rlabel m2contact 8649 4138 8649 4138 4 n_174
rlabel m2contact 8625 6346 8625 6346 4 n_297
rlabel m2contact 8601 1930 8601 1930 4 n_330
rlabel m2contact 8577 1954 8577 1954 4 n_193
rlabel m2contact 8553 6586 8553 6586 4 n_329
rlabel m2contact 8505 5386 8505 5386 4 n_268
rlabel m2contact 8481 5986 8481 5986 4 n_243
rlabel m2contact 8457 5386 8457 5386 4 n_225
rlabel m2contact 8457 3322 8457 3322 4 n_349
rlabel m2contact 8409 6682 8409 6682 4 n_293
rlabel m2contact 8409 6586 8409 6586 4 n_189
rlabel m2contact 8385 6658 8385 6658 4 n_47
rlabel m2contact 8385 1978 8385 1978 4 n_188
rlabel m2contact 8361 2002 8361 2002 4 n_160
rlabel m2contact 8361 6634 8361 6634 4 n_187
rlabel m2contact 8337 6610 8337 6610 4 n_290
rlabel m2contact 8313 6586 8313 6586 4 n_189
rlabel m2contact 8313 2026 8313 2026 4 n_279
rlabel m2contact 8289 2098 8289 2098 4 n_145
rlabel m2contact 8265 6562 8265 6562 4 n_43
rlabel m2contact 8265 3754 8265 3754 4 n_209
rlabel m2contact 8241 4018 8241 4018 4 n_42
rlabel m2contact 8217 3850 8217 3850 4 n_202
rlabel m2contact 8217 4186 8217 4186 4 n_22
rlabel m2contact 8193 5650 8193 5650 4 n_21
rlabel m2contact 8193 2098 8193 2098 4 n_21
rlabel m2contact 8169 2098 8169 2098 4 n_21
rlabel m2contact 8169 4714 8169 4714 4 n_265
rlabel m2contact 8145 3298 8145 3298 4 state[1]
rlabel m2contact 8121 3754 8121 3754 4 n_209
rlabel m2contact 8097 2122 8097 2122 4 n_184
rlabel m2contact 8073 3754 8073 3754 4 n_283
rlabel m2contact 8037 5434 8037 5434 4 n_190
rlabel m2contact 8037 2098 8037 2098 4 n_190
rlabel m2contact 8025 6538 8025 6538 4 n_151
rlabel m2contact 8025 2050 8025 2050 4 n_282
rlabel m2contact 8013 5098 8013 5098 4 OpcodeCondIn[4]
rlabel m2contact 8013 2122 8013 2122 4 OpcodeCondIn[4]
rlabel m2contact 8001 6514 8001 6514 4 n_354
rlabel m2contact 7977 2074 7977 2074 4 n_214
rlabel m2contact 7977 4762 7977 4762 4 n_380
rlabel m2contact 7953 2098 7953 2098 4 n_190
rlabel m2contact 7953 3586 7953 3586 4 n_357
rlabel m2contact 7929 5962 7929 5962 4 n_231
rlabel m2contact 7905 6514 7905 6514 4 n_26
rlabel m2contact 7881 5530 7881 5530 4 n_136
rlabel m2contact 7857 2122 7857 2122 4 OpcodeCondIn[4]
rlabel m2contact 7857 4906 7857 4906 4 state[0]
rlabel m2contact 7833 2914 7833 2914 4 n_115
rlabel m2contact 7809 5530 7809 5530 4 n_379
rlabel m2contact 7785 6514 7785 6514 4 n_26
rlabel m2contact 7785 4474 7785 4474 4 n_154
rlabel m2contact 7761 2146 7761 2146 4 n_352
rlabel m2contact 7737 6490 7737 6490 4 n_119
rlabel m2contact 7737 3058 7737 3058 4 OpcodeCondIn[2]
rlabel m2contact 7713 6466 7713 6466 4 n_118
rlabel m2contact 7713 6442 7713 6442 4 n_7
rlabel m2contact 7665 6418 7665 6418 4 n_27
rlabel m2contact 7641 2914 7641 2914 4 n_115
rlabel m2contact 7641 4834 7641 4834 4 n_367
rlabel m2contact 7617 6394 7617 6394 4 n_271
rlabel m2contact 7617 3250 7617 3250 4 n_44
rlabel m2contact 7593 6370 7593 6370 4 n_340
rlabel m2contact 7569 2170 7569 2170 4 n_285
rlabel m2contact 7521 2194 7521 2194 4 n_15
rlabel m2contact 7497 5986 7497 5986 4 n_243
rlabel m2contact 7497 4234 7497 4234 4 n_101
rlabel m2contact 7473 2914 7473 2914 4 n_115
rlabel m2contact 7449 6034 7449 6034 4 n_305
rlabel m2contact 7449 2194 7449 2194 4 n_305
rlabel m2contact 7425 2194 7425 2194 4 n_305
rlabel m2contact 7425 4234 7425 4234 4 n_310
rlabel m2contact 7401 3778 7401 3778 4 n_180
rlabel m2contact 7401 4090 7401 4090 4 n_309
rlabel m2contact 7377 5986 7377 5986 4 n_192
rlabel m2contact 7377 3874 7377 3874 4 stateSub[0]
rlabel m2contact 7353 5290 7353 5290 4 n_278
rlabel m2contact 7305 5290 7305 5290 4 n_303
rlabel m2contact 7281 2218 7281 2218 4 n_236
rlabel m2contact 7281 4042 7281 4042 4 n_72
rlabel m2contact 7257 2242 7257 2242 4 n_91
rlabel m2contact 7257 6250 7257 6250 4 n_296
rlabel m2contact 7233 6346 7233 6346 4 n_297
rlabel m2contact 7233 6322 7233 6322 4 n_107
rlabel m2contact 7185 2266 7185 2266 4 n_259
rlabel m2contact 7185 6298 7185 6298 4 n_33
rlabel m2contact 7161 2290 7161 2290 4 n_218
rlabel m2contact 7161 6274 7161 6274 4 n_499
rlabel m2contact 7137 4642 7137 4642 4 StatusReg[2]
rlabel m2contact 7065 6250 7065 6250 4 n_296
rlabel m2contact 7065 3874 7065 3874 4 stateSub[0]
rlabel m2contact 7017 5842 7017 5842 4 n_249
rlabel m2contact 6993 2314 6993 2314 4 n_230
rlabel m2contact 6969 2338 6969 2338 4 n_87
rlabel m2contact 6945 6226 6945 6226 4 n_68
rlabel m2contact 6945 3130 6945 3130 4 OpcodeCondIn[0]
rlabel m2contact 6921 6202 6921 6202 4 n_71
rlabel m2contact 6921 3226 6921 3226 4 OpcodeCondIn[1]
rlabel m2contact 6873 2362 6873 2362 4 n_49
rlabel m2contact 6873 6178 6873 6178 4 n_177
rlabel m2contact 6849 6154 6849 6154 4 n_176
rlabel m2contact 6825 3970 6825 3970 4 n_227
rlabel m2contact 6825 3634 6825 3634 4 OpcodeCondIn[6]
rlabel m2contact 6801 6034 6801 6034 4 n_305
rlabel m2contact 6801 2914 6801 2914 4 n_115
rlabel m2contact 6753 5722 6753 5722 4 n_270
rlabel m2contact 6753 3970 6753 3970 4 nOE
rlabel m2contact 6729 2434 6729 2434 4 n_261
rlabel m2contact 6729 2746 6729 2746 4 n_198
rlabel m2contact 6705 5146 6705 5146 4 n_252
rlabel m2contact 6705 4546 6705 4546 4 n_332
rlabel m2contact 6681 2986 6681 2986 4 n_167
rlabel m2contact 6657 5146 6657 5146 4 n_113
rlabel m2contact 6633 4498 6633 4498 4 n_232
rlabel m2contact 6609 5722 6609 5722 4 n_36
rlabel m2contact 6585 4474 6585 4474 4 n_154
rlabel m2contact 6561 2962 6561 2962 4 n_294
rlabel m2contact 6561 2986 6561 2986 4 n_162
rlabel m2contact 6537 5626 6537 5626 4 n_19
rlabel m2contact 6513 2386 6513 2386 4 n_81
rlabel m2contact 6513 4546 6513 4546 4 n_117
rlabel m2contact 6489 5626 6489 5626 4 n_76
rlabel m2contact 6489 4018 6489 4018 4 n_42
rlabel m2contact 6465 6130 6465 6130 4 n_59
rlabel m2contact 6465 4906 6465 4906 4 state[0]
rlabel m2contact 6417 3514 6417 3514 4 n_215
rlabel m2contact 6393 3514 6393 3514 4 n_215
rlabel m2contact 6369 2410 6369 2410 4 n_216
rlabel m2contact 6369 6034 6369 6034 4 n_305
rlabel m2contact 6345 3898 6345 3898 4 n_14
rlabel m2contact 6321 6106 6321 6106 4 n_262
rlabel m2contact 6297 2434 6297 2434 4 n_261
rlabel m2contact 6273 2770 6273 2770 4 n_52
rlabel m2contact 6225 6082 6225 6082 4 n_257
rlabel m2contact 6177 6058 6177 6058 4 n_166
rlabel m2contact 6153 4618 6153 4618 4 n_212
rlabel m2contact 6129 6034 6129 6034 4 n_305
rlabel m2contact 6129 4642 6129 4642 4 StatusReg[2]
rlabel m2contact 6081 2458 6081 2458 4 n_498
rlabel m2contact 6081 4642 6081 4642 4 n_223
rlabel m2contact 6057 3706 6057 3706 4 n_222
rlabel m2contact 6033 6010 6033 6010 4 n_195
rlabel m2contact 5985 5986 5985 5986 4 n_192
rlabel m2contact 5961 3730 5961 3730 4 n_130
rlabel m2contact 5937 5962 5937 5962 4 n_231
rlabel m2contact 5889 3034 5889 3034 4 n_31
rlabel m2contact 5841 4402 5841 4402 4 n_58
rlabel m2contact 5817 3034 5817 3034 4 n_18
rlabel m2contact 5769 4402 5769 4402 4 n_364
rlabel m2contact 5721 5938 5721 5938 4 n_371
rlabel m2contact 5697 2482 5697 2482 4 n_326
rlabel m2contact 5649 5914 5649 5914 4 n_69
rlabel m2contact 5601 2506 5601 2506 4 LrWe
rlabel m2contact 5601 3634 5601 3634 4 OpcodeCondIn[6]
rlabel m2contact 5577 2530 5577 2530 4 n_229
rlabel m2contact 5577 5098 5577 5098 4 OpcodeCondIn[4]
rlabel m2contact 5529 5098 5529 5098 4 n_129
rlabel m2contact 5505 3730 5505 3730 4 n_130
rlabel m2contact 5481 2674 5481 2674 4 n_228
rlabel m2contact 5481 3778 5481 3778 4 n_180
rlabel m2contact 5457 3514 5457 3514 4 n_215
rlabel m2contact 5433 5026 5433 5026 4 n_24
rlabel m2contact 5409 2554 5409 2554 4 n_336
rlabel m2contact 5385 5890 5385 5890 4 n_335
rlabel m2contact 5361 5890 5361 5890 4 n_335
rlabel m2contact 5361 5170 5361 5170 4 n_170
rlabel m2contact 5337 4594 5337 4594 4 n_255
rlabel m2contact 5313 2578 5313 2578 4 n_165
rlabel m2contact 5313 5866 5313 5866 4 n_260
rlabel m2contact 5289 4594 5289 4594 4 n_183
rlabel m2contact 5265 5842 5265 5842 4 n_249
rlabel m2contact 5217 5818 5217 5818 4 n_186
rlabel m2contact 5217 2602 5217 2602 4 n_56
rlabel m2contact 5193 5794 5193 5794 4 n_144
rlabel m2contact 5169 2626 5169 2626 4 n_156
rlabel m2contact 5145 2650 5145 2650 4 n_178
rlabel m2contact 5097 5770 5097 5770 4 n_169
rlabel m2contact 5097 5194 5097 5194 4 n_54
rlabel m2contact 5073 3610 5073 3610 4 n_344
rlabel m2contact 5049 5746 5049 5746 4 n_29
rlabel m2contact 5025 5722 5025 5722 4 n_36
rlabel m2contact 5001 2674 5001 2674 4 n_228
rlabel m2contact 5001 5698 5001 5698 4 OpcodeCondIn[3]
rlabel m2contact 4977 2698 4977 2698 4 n_10
rlabel m2contact 4929 5674 4929 5674 4 n_103
rlabel m2contact 4929 2722 4929 2722 4 n_273
rlabel m2contact 4881 2746 4881 2746 4 n_198
rlabel m2contact 4881 2914 4881 2914 4 n_115
rlabel m2contact 4857 5650 4857 5650 4 n_21
rlabel m2contact 4809 5626 4809 5626 4 n_76
rlabel m2contact 4809 3898 4809 3898 4 n_14
rlabel m2contact 4785 2770 4785 2770 4 n_52
rlabel m2contact 4785 3058 4785 3058 4 OpcodeCondIn[2]
rlabel m2contact 4761 5602 4761 5602 4 n_37
rlabel m2contact 4713 5578 4713 5578 4 n_116
rlabel m2contact 4689 2794 4689 2794 4 n_122
rlabel m2contact 4689 4498 4689 4498 4 n_232
rlabel m2contact 4665 5554 4665 5554 4 n_89
rlabel m2contact 4665 5530 4665 5530 4 n_379
rlabel m2contact 4617 5506 4617 5506 4 n_323
rlabel m2contact 4593 5002 4593 5002 4 stateSub[1]
rlabel m2contact 4593 4498 4593 4498 4 n_232
rlabel m2contact 4569 2818 4569 2818 4 n_291
rlabel m2contact 4521 4426 4521 4426 4 n_241
rlabel m2contact 4497 5482 4497 5482 4 n_179
rlabel m2contact 4497 5458 4497 5458 4 n_62
rlabel m2contact 4473 3778 4473 3778 4 n_180
rlabel m2contact 4449 5434 4449 5434 4 n_190
rlabel m2contact 4449 2842 4449 2842 4 n_60
rlabel m2contact 4425 2866 4425 2866 4 n_61
rlabel m2contact 4401 2890 4401 2890 4 n_208
rlabel m2contact 4377 5410 4377 5410 4 n_133
rlabel m2contact 4377 5386 4377 5386 4 n_225
rlabel m2contact 4353 5362 4353 5362 4 n_207
rlabel m2contact 4305 5338 4305 5338 4 n_356
rlabel m2contact 4281 5314 4281 5314 4 n_93
rlabel m2contact 4281 3946 4281 3946 4 n_181
rlabel m2contact 4257 5290 4257 5290 4 n_303
rlabel m2contact 4233 5266 4233 5266 4 n_302
rlabel m2contact 4233 2914 4233 2914 4 n_115
rlabel m2contact 4209 5242 4209 5242 4 n_112
rlabel m2contact 4209 2938 4209 2938 4 n_159
rlabel m2contact 4161 5218 4161 5218 4 n_175
rlabel m2contact 4137 5194 4137 5194 4 n_54
rlabel m2contact 4137 2962 4137 2962 4 n_294
rlabel m2contact 4113 2986 4113 2986 4 n_162
rlabel m2contact 4113 4138 4113 4138 4 n_174
rlabel m2contact 4065 4138 4065 4138 4 n_171
rlabel m2contact 4041 5170 4041 5170 4 n_170
rlabel m2contact 4041 4138 4041 4138 4 n_171
rlabel m2contact 4017 3010 4017 3010 4 n_46
rlabel m2contact 4017 5146 4017 5146 4 n_113
rlabel m2contact 3993 4138 3993 4138 4 n_124
rlabel m2contact 3945 3034 3945 3034 4 n_18
rlabel m2contact 3945 5122 3945 5122 4 n_351
rlabel m2contact 3921 3058 3921 3058 4 OpcodeCondIn[2]
rlabel m2contact 3921 5098 3921 5098 4 n_129
rlabel m2contact 3897 3082 3897 3082 4 n_286
rlabel m2contact 3873 5074 3873 5074 4 n_245
rlabel m2contact 3873 3106 3873 3106 4 stateSub[2]
rlabel m2contact 3849 5050 3849 5050 4 n_240
rlabel m2contact 3849 3130 3849 3130 4 OpcodeCondIn[0]
rlabel m2contact 3801 3154 3801 3154 4 AluOR[0]
rlabel m2contact 3777 3178 3777 3178 4 Op2Sel[0]
rlabel m2contact 3777 4834 3777 4834 4 n_367
rlabel m2contact 3753 3202 3753 3202 4 n_206
rlabel m2contact 3753 4114 3753 4114 4 n_359
rlabel m2contact 3705 5026 3705 5026 4 n_24
rlabel m2contact 3681 3874 3681 3874 4 stateSub[0]
rlabel m2contact 3657 5002 3657 5002 4 stateSub[1]
rlabel m2contact 3633 3226 3633 3226 4 OpcodeCondIn[1]
rlabel m2contact 3609 3250 3609 3250 4 n_44
rlabel m2contact 3609 3394 3609 3394 4 n_248
rlabel m2contact 3585 4978 3585 4978 4 n_247
rlabel m2contact 3561 4954 3561 4954 4 n_163
rlabel m2contact 3561 3394 3561 3394 4 SysBus[2]
rlabel m2contact 3513 3274 3513 3274 4 n_100
rlabel m2contact 3489 4930 3489 4930 4 n_99
rlabel m2contact 3465 4906 3465 4906 4 state[0]
rlabel m2contact 3417 3298 3417 3298 4 state[1]
rlabel m2contact 3417 4882 3417 4882 4 n_157
rlabel m2contact 3393 4858 3393 4858 4 n_137
rlabel m2contact 3369 3322 3369 3322 4 n_349
rlabel m2contact 3369 3346 3369 3346 4 n_82
rlabel m2contact 3321 3370 3321 3370 4 RegWe
rlabel m2contact 3297 4834 3297 4834 4 n_367
rlabel m2contact 3273 4810 3273 4810 4 n_387
rlabel m2contact 3249 4786 3249 4786 4 n_304
rlabel m2contact 3225 4762 3225 4762 4 n_380
rlabel m2contact 3177 4738 3177 4738 4 n_264
rlabel m2contact 3153 3394 3153 3394 4 SysBus[2]
rlabel m2contact 3129 4714 3129 4714 4 n_265
rlabel m2contact 3081 3418 3081 3418 4 n_355
rlabel m2contact 3057 3442 3057 3442 4 n_134
rlabel m2contact 3033 4690 3033 4690 4 n_284
rlabel m2contact 3009 3466 3009 3466 4 n_313
rlabel m2contact 3009 4666 3009 4666 4 n_301
rlabel m2contact 2985 4642 2985 4642 4 n_223
rlabel m2contact 2913 4618 2913 4618 4 n_212
rlabel m2contact 2889 4594 2889 4594 4 n_183
rlabel m2contact 2865 4570 2865 4570 4 n_127
rlabel m2contact 2865 3706 2865 3706 4 n_222
rlabel m2contact 2841 3946 2841 3946 4 n_181
rlabel m2contact 2817 4546 2817 4546 4 n_117
rlabel m2contact 2793 3946 2793 3946 4 ALE
rlabel m2contact 2769 3490 2769 3490 4 n_35
rlabel m2contact 2745 3514 2745 3514 4 n_215
rlabel m2contact 2745 4522 2745 4522 4 n_77
rlabel m2contact 2721 3538 2721 3538 4 n_299
rlabel m2contact 2697 4138 2697 4138 4 n_124
rlabel m2contact 2673 3562 2673 3562 4 PcSel[1]
rlabel m2contact 2673 4498 2673 4498 4 n_232
rlabel m2contact 2649 3586 2649 3586 4 n_357
rlabel m2contact 2649 4474 2649 4474 4 n_154
rlabel m2contact 2625 3610 2625 3610 4 n_344
rlabel m2contact 2601 4450 2601 4450 4 n_292
rlabel m2contact 2577 4426 2577 4426 4 n_241
rlabel m2contact 2553 4402 2553 4402 4 n_364
rlabel m2contact 2529 3634 2529 3634 4 OpcodeCondIn[6]
rlabel m2contact 2529 4378 2529 4378 4 n_383
rlabel m2contact 2505 4354 2505 4354 4 n_374
rlabel m2contact 2505 4042 2505 4042 4 n_72
rlabel m2contact 2457 3658 2457 3658 4 n_114
rlabel m2contact 2457 3682 2457 3682 4 n_312
rlabel m2contact 2433 3706 2433 3706 4 n_222
rlabel m2contact 2433 4330 2433 4330 4 n_311
rlabel m2contact 2409 3730 2409 3730 4 n_130
rlabel m2contact 2409 3754 2409 3754 4 n_283
rlabel m2contact 2361 3778 2361 3778 4 n_180
rlabel m2contact 2361 3802 2361 3802 4 n_8
rlabel m2contact 2337 4306 2337 4306 4 OpcodeCondIn[7]
rlabel m2contact 2313 3826 2313 3826 4 n_138
rlabel m2contact 2313 3874 2313 3874 4 stateSub[0]
rlabel m2contact 2289 3850 2289 3850 4 n_202
rlabel m2contact 2241 4282 2241 4282 4 n_324
rlabel m2contact 2241 4258 2241 4258 4 nIRQ
rlabel m2contact 2193 4234 2193 4234 4 n_310
rlabel m2contact 2121 4210 2121 4210 4 n_70
rlabel m2contact 2097 3874 2097 3874 4 stateSub[0]
rlabel m2contact 2073 4186 2073 4186 4 n_22
rlabel m2contact 2049 3898 2049 3898 4 n_14
rlabel m2contact 2001 4162 2001 4162 4 n_210
rlabel m2contact 1953 4138 1953 4138 4 n_124
rlabel m2contact 1905 4114 1905 4114 4 n_359
rlabel m2contact 1857 4090 1857 4090 4 n_309
rlabel m2contact 1833 4066 1833 4066 4 n_281
rlabel m2contact 1785 3922 1785 3922 4 nME
rlabel m2contact 1737 3946 1737 3946 4 ALE
rlabel m2contact 1665 4042 1665 4042 4 n_72
rlabel m2contact 1617 4018 1617 4018 4 n_42
rlabel m2contact 27321 8043 27321 8043 6 Flags[2]
rlabel m2contact 27321 7947 27321 7947 6 Flags[2]
rlabel m2contact 27297 7947 27297 7947 6 Flags[0]
rlabel m2contact 27297 7899 27297 7899 6 Flags[0]
rlabel m2contact 27273 8019 27273 8019 6 Flags[3]
rlabel m2contact 27273 7971 27273 7971 6 Flags[3]
rlabel m2contact 27273 7923 27273 7923 6 Flags[1]
rlabel m2contact 27273 7899 27273 7899 6 Flags[1]
rlabel m2contact 27249 8019 27249 8019 6 Flags[3]
rlabel metal2 27219 8019 27219 8019 6 StatusRegEn
rlabel m2contact 27201 8019 27201 8019 6 StatusRegEn
rlabel m2contact 25629 8019 25629 8019 6 StatusReg[3]
rlabel m2contact 24777 7923 24777 7923 6 StatusReg[2]
rlabel m2contact 24729 8067 24729 8067 6 StatusReg[0]
rlabel m2contact 24273 8019 24273 8019 6 StatusReg[3]
rlabel m2contact 24129 8091 24129 8091 6 PcEn
rlabel m2contact 23925 8019 23925 8019 6 StatusReg[1]
rlabel m2contact 23901 8067 23901 8067 6 StatusReg[0]
rlabel m2contact 23793 8043 23793 8043 6 Flags[2]
rlabel m2contact 22497 8115 22497 8115 6 Op1Sel
rlabel m2contact 22221 8067 22221 8067 6 AluEn
rlabel m2contact 21369 8043 21369 8043 6 AluWe
rlabel m2contact 20517 7971 20517 7971 6 Op2Sel[1]
rlabel metal2 20235 8139 20235 8139 6 Op2Sel[0]
rlabel m2contact 20217 8139 20217 8139 6 Op2Sel[0]
rlabel m2contact 19857 7923 19857 7923 6 StatusReg[2]
rlabel m2contact 19425 7947 19425 7947 6 Flags[0]
rlabel m2contact 18813 8115 18813 8115 6 Op1Sel
rlabel m2contact 18789 8091 18789 8091 6 PcEn
rlabel m2contact 18225 7995 18225 7995 6 CFlag
rlabel m2contact 17109 8163 17109 8163 6 WdSel
rlabel m2contact 17025 7947 17025 7947 6 OpcodeCondIn[5]
rlabel m2contact 16257 8139 16257 8139 6 PcWe
rlabel m2contact 16185 8043 16185 8043 6 AluWe
rlabel m2contact 15417 8043 15417 8043 6 PcSel[1]
rlabel m2contact 15405 8091 15405 8091 6 PcSel[2]
rlabel m2contact 15381 8043 15381 8043 6 PcSel[1]
rlabel metal2 14427 8043 14427 8043 6 PcSel[0]
rlabel m2contact 14409 8043 14409 8043 6 PcSel[0]
rlabel m2contact 13713 8043 13713 8043 4 OpcodeCondIn[1]
rlabel m2contact 13065 8019 13065 8019 4 StatusReg[1]
rlabel m2contact 13017 7995 13017 7995 4 CFlag
rlabel m2contact 12969 7923 12969 7923 4 MemEn
rlabel m2contact 12837 8019 12837 8019 4 LrEn
rlabel metal2 12531 8187 12531 8187 4 LrWe
rlabel m2contact 12513 8187 12513 8187 4 LrWe
rlabel m2contact 12033 8163 12033 8163 4 WdSel
rlabel metal2 11499 8163 11499 8163 4 LrSel
rlabel m2contact 11481 8163 11481 8163 4 LrSel
rlabel m2contact 11049 8091 11049 8091 4 PcSel[2]
rlabel metal2 10731 8091 10731 8091 4 ImmSel
rlabel m2contact 10713 8091 10713 8091 4 ImmSel
rlabel m2contact 9825 8091 9825 8091 4 OpcodeCondIn[0]
rlabel metal2 9795 8163 9795 8163 4 IrWe
rlabel m2contact 9777 8163 9777 8163 4 IrWe
rlabel m2contact 9345 7923 9345 7923 4 MemEn
rlabel m2contact 8673 7923 8673 7923 4 OpcodeCondIn[7]
rlabel m2contact 8577 7899 8577 7899 4 Flags[1]
rlabel m2contact 8481 7923 8481 7923 4 OpcodeCondIn[7]
rlabel m2contact 8049 8139 8049 8139 4 PcWe
rlabel m2contact 7665 7971 7665 7971 4 Op2Sel[1]
rlabel m2contact 6789 7971 6789 7971 4 OpcodeCondIn[6]
rlabel m2contact 6753 7947 6753 7947 4 OpcodeCondIn[5]
rlabel m2contact 5721 8115 5721 8115 4 Op1Sel
rlabel m2contact 5601 7971 5601 7971 4 OpcodeCondIn[6]
rlabel metal2 5595 8115 5595 8115 4 OpcodeCondIn[4]
rlabel m2contact 5577 8115 5577 8115 4 OpcodeCondIn[4]
rlabel m2contact 5385 7995 5385 7995 4 CFlag
rlabel m2contact 5121 8019 5121 8019 4 LrEn
rlabel metal2 5019 8019 5019 8019 4 OpcodeCondIn[3]
rlabel m2contact 5001 8019 5001 8019 4 OpcodeCondIn[3]
rlabel m2contact 4785 8019 4785 8019 4 OpcodeCondIn[2]
rlabel m2contact 4161 8019 4161 8019 4 OpcodeCondIn[2]
rlabel m2contact 3297 8043 3297 8043 4 OpcodeCondIn[1]
rlabel m2contact 2601 8067 2601 8067 4 AluEn
rlabel m2contact 2433 8091 2433 8091 4 OpcodeCondIn[0]
rlabel m2contact 1785 8067 1785 8067 4 nME
rlabel m2contact 1737 8091 1737 8091 4 ALE
rlabel metal2 27207 8204 27219 8204 6 StatusRegEn
rlabel metal2 25623 8204 25635 8204 6 StatusReg[3]
rlabel metal2 24771 8204 24783 8204 6 StatusReg[2]
rlabel metal2 23919 8204 23931 8204 6 StatusReg[1]
rlabel metal2 23895 8204 23907 8204 6 StatusReg[0]
rlabel metal2 22215 8204 22227 8204 6 AluEn
rlabel metal2 21363 8204 21375 8204 6 AluWe
rlabel metal2 20511 8204 20523 8204 6 Op2Sel[1]
rlabel metal2 20223 8204 20235 8204 6 Op2Sel[0]
rlabel metal2 18807 8204 18819 8204 6 Op1Sel
rlabel metal2 18783 8204 18795 8204 6 PcEn
rlabel metal2 17103 8204 17115 8204 6 WdSel
rlabel metal2 16251 8204 16263 8204 6 PcWe
rlabel metal2 15399 8204 15411 8204 6 PcSel[2]
rlabel metal2 15375 8204 15387 8204 6 PcSel[1]
rlabel metal2 14415 8204 14427 8204 6 PcSel[0]
rlabel metal2 12831 8204 12843 8204 4 LrEn
rlabel metal2 12519 8204 12531 8204 4 LrWe
rlabel metal2 11487 8204 11499 8204 4 LrSel
rlabel metal2 10719 8204 10731 8204 4 ImmSel
rlabel metal2 9783 8204 9795 8204 4 IrWe
rlabel metal2 9339 8204 9351 8204 4 MemEn
rlabel metal2 8475 8204 8487 8204 4 OpcodeCondIn[7]
rlabel metal2 6783 8204 6795 8204 4 OpcodeCondIn[6]
rlabel metal2 6747 8204 6759 8204 4 OpcodeCondIn[5]
rlabel metal2 5583 8204 5595 8204 4 OpcodeCondIn[4]
rlabel metal2 5007 8204 5019 8204 4 OpcodeCondIn[3]
rlabel metal2 4155 8204 4167 8204 4 OpcodeCondIn[2]
rlabel metal2 3291 8204 3303 8204 4 OpcodeCondIn[1]
rlabel metal2 2427 8204 2439 8204 4 OpcodeCondIn[0]
rlabel metal2 23919 0 23931 0 8 SysBus[3]
rlabel metal2 14427 0 14439 0 8 SysBus[2]
rlabel metal2 11175 0 11187 0 2 SysBus[1]
rlabel metal2 7983 0 7995 0 2 SysBus[0]
rlabel metal2 27735 419 27735 431 8 RegWe
rlabel metal2 27735 59 27735 71 8 AluOR[0]
rlabel metal2 27735 35 27735 47 8 AluOR[1]
rlabel metal2 27735 11 27735 23 8 ENB
rlabel metal2 27735 2884 27735 2896 6 Rs1Sel[0]
rlabel metal2 27735 1636 27735 1648 6 Rs1Sel[1]
rlabel metal2 27735 1612 27735 1624 6 RwSel[0]
rlabel metal2 27735 1588 27735 1600 6 RwSel[1]
rlabel metal2 27735 7989 27735 8001 6 CFlag
rlabel metal2 27735 7965 27735 7977 6 Flags[3]
rlabel metal2 27735 7941 27735 7953 6 Flags[2]
rlabel metal2 27735 7917 27735 7929 6 Flags[1]
rlabel metal2 27735 7893 27735 7905 6 Flags[0]
rlabel metal2 0 59 0 71 2 nWE
rlabel metal2 0 35 0 47 2 nIRQ
rlabel metal2 0 3988 0 4000 4 nWait
rlabel metal2 0 3964 0 3976 4 nOE
rlabel metal2 0 8085 0 8097 4 ALE
rlabel metal2 0 8061 0 8073 4 nME
rlabel metal2 123 8204 323 8204 5 Vdd!
rlabel metal2 411 8204 423 8204 5 nReset
rlabel metal2 387 8204 399 8204 5 Clock
rlabel metal2 363 8204 375 8204 5 Test
rlabel metal2 339 8204 351 8204 5 SDO
rlabel metal2 27387 0 27587 0 1 GND!
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 339 0 351 0 1 SDI
rlabel space 123 0 324 0 1 Vdd!
rlabel metal2 27387 8204 27587 8204 5 GND!
<< end >>
