magic
tech c035u
timestamp 1394103428
<< error_ps >>
rect 2416 1680 2422 1690
rect 2426 1485 2432 1680
<< metal1 >>
rect 12588 6553 13145 6563
rect 12588 6368 12598 6553
rect 13105 6508 13145 6518
rect 12997 6488 13145 6498
rect 12875 6463 13145 6473
rect 12718 6430 13145 6442
rect 12811 6406 13145 6416
rect 12655 6379 13145 6390
rect 12442 6358 12598 6368
rect 12202 6328 13145 6338
rect 11963 6303 13092 6313
rect 11723 6280 12981 6290
rect 10235 6256 11538 6266
rect 11557 6256 11780 6266
rect 11794 6256 12020 6266
rect 12034 6256 12260 6266
rect 10522 6231 10627 6241
rect 10642 6231 11108 6241
rect 11122 6231 11588 6241
rect 11602 6231 12068 6241
rect 10356 6205 11084 6215
rect 11098 6205 11324 6215
rect 11338 6205 12044 6215
rect 12058 6205 12284 6215
rect 17911 6202 18468 6212
rect 10283 6170 10580 6180
rect 10594 6170 10820 6180
rect 10834 6170 11060 6180
rect 11074 6170 11296 6180
rect 11483 6168 12861 6178
rect 10475 6148 10867 6158
rect 11244 6146 12703 6156
rect 10402 6119 10603 6130
rect 10619 6119 10844 6130
rect 10858 6119 11564 6130
rect 11578 6119 11804 6130
rect 11003 6094 12795 6104
rect 10926 6071 11348 6081
rect 11363 6071 11828 6081
rect 11842 6071 12308 6081
rect 10762 6049 12641 6060
rect 17911 6017 17921 6202
rect 18428 6157 18468 6167
rect 18320 6137 18468 6147
rect 18198 6112 18468 6122
rect 18041 6079 18468 6091
rect 18134 6055 18468 6065
rect 17978 6028 18468 6039
rect 17765 6007 17921 6017
rect 17525 5977 18468 5987
rect 10666 5947 10700 5957
rect 10906 5948 10940 5958
rect 11146 5948 11180 5958
rect 11387 5953 11420 5963
rect 11626 5953 11660 5963
rect 11866 5953 11900 5963
rect 12106 5953 12140 5963
rect 12347 5953 12379 5963
rect 17286 5952 18415 5962
rect 17046 5929 18304 5939
rect 6259 5914 6816 5924
rect 6259 5729 6269 5914
rect 15558 5905 16861 5915
rect 16880 5905 17103 5915
rect 17117 5905 17343 5915
rect 17357 5905 17583 5915
rect 6776 5869 6816 5879
rect 10172 5863 10197 5888
rect 15845 5880 15950 5890
rect 15965 5880 16431 5890
rect 16445 5880 16911 5890
rect 16925 5880 17391 5890
rect 6668 5849 6816 5859
rect 15679 5854 16407 5864
rect 16421 5854 16647 5864
rect 16661 5854 17367 5864
rect 17381 5854 17607 5864
rect 6546 5824 6816 5834
rect 15606 5819 15903 5829
rect 15917 5819 16143 5829
rect 16157 5819 16383 5829
rect 16397 5819 16619 5829
rect 16806 5817 18184 5827
rect 6389 5791 6816 5803
rect 15798 5797 16190 5807
rect 16567 5795 18026 5805
rect 6482 5767 6816 5777
rect 15725 5768 15926 5779
rect 15942 5768 16167 5779
rect 16181 5768 16887 5779
rect 16901 5768 17127 5779
rect 6326 5740 6816 5751
rect 16326 5743 18118 5753
rect 6113 5719 6269 5729
rect 16249 5720 16671 5730
rect 16686 5720 17151 5730
rect 17165 5720 17631 5730
rect 5873 5689 6816 5699
rect 16085 5698 17964 5709
rect 5634 5664 6763 5674
rect 5394 5641 6652 5651
rect 3906 5617 5209 5627
rect 5228 5617 5451 5627
rect 5465 5617 5691 5627
rect 5705 5617 5931 5627
rect 4193 5592 4298 5602
rect 4313 5592 4779 5602
rect 4793 5592 5259 5602
rect 5273 5592 5739 5602
rect 15989 5596 16023 5606
rect 16229 5597 16263 5607
rect 16469 5597 16503 5607
rect 16710 5602 16743 5612
rect 16949 5602 16983 5612
rect 17189 5602 17223 5612
rect 17429 5602 17463 5612
rect 17670 5602 17702 5612
rect 4027 5566 4755 5576
rect 4769 5566 4995 5576
rect 5009 5566 5715 5576
rect 5729 5566 5955 5576
rect 3954 5531 4251 5541
rect 4265 5531 4491 5541
rect 4505 5531 4731 5541
rect 4745 5531 4967 5541
rect 5154 5529 6532 5539
rect 4146 5509 4538 5519
rect 4915 5507 6374 5517
rect 15495 5512 15520 5537
rect 4073 5480 4274 5491
rect 4290 5480 4515 5491
rect 4529 5480 5235 5491
rect 5249 5480 5475 5491
rect 4674 5455 6466 5465
rect 4597 5432 5019 5442
rect 5034 5432 5499 5442
rect 5513 5432 5979 5442
rect 4433 5410 6312 5421
rect 4337 5308 4371 5318
rect 4577 5309 4611 5319
rect 4817 5309 4851 5319
rect 5058 5314 5091 5324
rect 5297 5314 5331 5324
rect 5537 5314 5571 5324
rect 5777 5314 5811 5324
rect 6018 5314 6050 5324
rect 3843 5224 3868 5249
rect 10172 5218 10197 5243
rect 10172 5195 10197 5205
rect 10172 5149 10197 5159
rect 15495 4867 15520 4892
rect 15495 4844 15520 4854
rect 15495 4798 15520 4808
rect 3843 4579 3868 4604
rect 3843 4556 3868 4566
rect 3843 4510 3868 4520
rect 13455 1865 14528 1875
rect 12303 1837 14528 1847
rect 3133 1785 6670 1795
rect 9998 1781 14330 1791
rect 11150 1717 14246 1727
rect 2422 1680 14400 1690
rect 2422 1485 2426 1680
rect 3091 1655 13248 1665
rect 2933 1635 12096 1645
rect 2825 1615 10944 1625
rect 2703 1590 9792 1600
rect 2546 1557 8639 1569
rect 8847 1567 14528 1577
rect 2639 1533 7487 1543
rect 2483 1506 6335 1517
rect 6005 1485 14184 1495
rect 2422 1455 3078 1465
rect 6005 1455 13031 1465
rect 2422 1430 2920 1440
rect 6005 1430 11880 1440
rect 14261 1430 14516 1440
rect 2422 1407 2809 1417
rect 6006 1407 10728 1417
rect 14344 1407 14516 1417
rect 7695 1340 13937 1350
rect 2422 1295 2689 1305
rect 6006 1295 9574 1305
rect 2422 1273 2531 1283
rect 6006 1273 8424 1283
rect 6543 1250 7428 1260
rect 2422 1221 2623 1231
rect 6006 1221 7272 1231
rect 7418 1231 7428 1250
rect 7418 1221 14516 1231
rect 2422 1176 2469 1187
rect 6006 1176 6120 1187
rect 6690 1180 14516 1190
rect 13951 1151 14516 1161
rect 3638 1107 3753 1117
rect 6006 1107 6048 1117
rect 6062 1107 6264 1117
rect 7069 1094 7200 1104
rect 7214 1094 7416 1104
rect 8221 1094 8352 1104
rect 8366 1094 8568 1104
rect 9373 1094 9504 1104
rect 9518 1094 9720 1104
rect 10525 1094 10656 1104
rect 10670 1094 10872 1104
rect 11677 1094 11808 1104
rect 11822 1094 12024 1104
rect 12829 1094 12960 1104
rect 12974 1094 13176 1104
rect 13981 1094 14112 1104
rect 14126 1094 14328 1104
rect 0 75 2328 85
rect 2342 75 16815 85
rect 0 40 6191 50
rect 6206 40 7343 50
rect 7358 40 8495 50
rect 8510 40 9648 50
rect 9663 40 10798 50
rect 10816 40 11950 50
rect 11968 40 13102 50
rect 13120 40 14256 50
rect 14270 40 16815 50
rect 0 5 6408 15
rect 6422 5 7560 15
rect 7574 5 8712 15
rect 8726 5 9864 15
rect 9879 5 11015 15
rect 11033 5 12167 15
rect 12185 5 13319 15
rect 13337 5 14472 15
rect 14486 5 16815 15
<< m2contact >>
rect 12428 6357 12442 6371
rect 13090 6508 13105 6522
rect 12980 6486 12997 6500
rect 12860 6460 12875 6475
rect 12702 6427 12718 6443
rect 12797 6405 12811 6419
rect 12641 6378 12655 6392
rect 12188 6326 12202 6340
rect 11948 6301 11963 6315
rect 13092 6302 13106 6316
rect 11707 6277 11723 6292
rect 12981 6278 12995 6292
rect 10221 6255 10235 6269
rect 11538 6254 11557 6270
rect 11780 6253 11794 6267
rect 12020 6255 12034 6269
rect 12260 6255 12275 6269
rect 10508 6230 10522 6244
rect 10627 6230 10642 6244
rect 11108 6230 11122 6244
rect 11588 6230 11602 6244
rect 12068 6229 12083 6243
rect 10339 6203 10356 6217
rect 11084 6205 11098 6219
rect 11324 6204 11338 6218
rect 12044 6204 12058 6218
rect 12284 6203 12299 6217
rect 10268 6168 10283 6182
rect 10580 6168 10594 6182
rect 10820 6169 10834 6183
rect 11060 6169 11074 6183
rect 11296 6168 11313 6185
rect 11466 6166 11483 6180
rect 12861 6167 12875 6181
rect 10460 6146 10475 6160
rect 10867 6142 10883 6160
rect 11227 6143 11244 6158
rect 12703 6144 12717 6158
rect 10388 6118 10402 6132
rect 10603 6117 10619 6131
rect 10844 6118 10858 6132
rect 11564 6118 11578 6132
rect 11804 6118 11818 6132
rect 10987 6092 11003 6106
rect 12795 6093 12809 6107
rect 10912 6070 10926 6084
rect 11348 6070 11363 6084
rect 11828 6070 11842 6084
rect 12308 6070 12322 6084
rect 10748 6049 10762 6063
rect 12641 6048 12655 6062
rect 17751 6006 17765 6020
rect 18413 6157 18428 6171
rect 18303 6135 18320 6149
rect 18183 6109 18198 6124
rect 18025 6076 18041 6092
rect 18120 6054 18134 6068
rect 17964 6027 17978 6041
rect 17511 5975 17525 5989
rect 10652 5944 10666 5958
rect 10700 5944 10714 5958
rect 10892 5947 10906 5961
rect 10940 5946 10954 5960
rect 11132 5947 11146 5961
rect 11180 5947 11194 5961
rect 11372 5951 11387 5965
rect 11420 5951 11435 5965
rect 11611 5951 11626 5965
rect 11660 5951 11675 5965
rect 11852 5952 11866 5966
rect 11900 5951 11914 5965
rect 12092 5952 12106 5966
rect 12140 5951 12154 5965
rect 12332 5951 12347 5965
rect 12379 5951 12394 5965
rect 17271 5950 17286 5964
rect 18415 5951 18429 5965
rect 17030 5926 17046 5941
rect 18304 5927 18318 5941
rect 6099 5718 6113 5732
rect 15544 5904 15558 5918
rect 16861 5903 16880 5919
rect 17103 5902 17117 5916
rect 17343 5904 17357 5918
rect 17583 5904 17598 5918
rect 6761 5869 6776 5883
rect 15831 5879 15845 5893
rect 15950 5879 15965 5893
rect 16431 5879 16445 5893
rect 16911 5879 16925 5893
rect 17391 5878 17406 5892
rect 6651 5847 6668 5861
rect 15662 5852 15679 5866
rect 16407 5854 16421 5868
rect 16647 5853 16661 5867
rect 17367 5853 17381 5867
rect 17607 5852 17622 5866
rect 6531 5821 6546 5836
rect 15591 5817 15606 5831
rect 15903 5817 15917 5831
rect 16143 5818 16157 5832
rect 16383 5818 16397 5832
rect 16619 5817 16636 5834
rect 16789 5815 16806 5829
rect 18184 5816 18198 5830
rect 6373 5788 6389 5804
rect 15783 5795 15798 5809
rect 16190 5791 16206 5809
rect 16550 5792 16567 5807
rect 18026 5793 18040 5807
rect 6468 5766 6482 5780
rect 15711 5767 15725 5781
rect 15926 5766 15942 5780
rect 16167 5767 16181 5781
rect 16887 5767 16901 5781
rect 17127 5767 17141 5781
rect 6312 5739 6326 5753
rect 16310 5741 16326 5755
rect 18118 5742 18132 5756
rect 16235 5719 16249 5733
rect 16671 5719 16686 5733
rect 17151 5719 17165 5733
rect 17631 5719 17645 5733
rect 5859 5687 5873 5701
rect 16071 5698 16085 5712
rect 17964 5697 17978 5711
rect 5619 5662 5634 5676
rect 6763 5663 6777 5677
rect 5378 5638 5394 5653
rect 6652 5639 6666 5653
rect 3892 5616 3906 5630
rect 5209 5615 5228 5631
rect 5451 5614 5465 5628
rect 5691 5616 5705 5630
rect 5931 5616 5946 5630
rect 4179 5591 4193 5605
rect 4298 5591 4313 5605
rect 4779 5591 4793 5605
rect 5259 5591 5273 5605
rect 5739 5590 5754 5604
rect 15975 5593 15989 5607
rect 16023 5593 16037 5607
rect 16215 5596 16229 5610
rect 16263 5595 16277 5609
rect 16455 5596 16469 5610
rect 16503 5596 16517 5610
rect 16695 5600 16710 5614
rect 16743 5600 16758 5614
rect 16934 5600 16949 5614
rect 16983 5600 16998 5614
rect 17175 5601 17189 5615
rect 17223 5600 17237 5614
rect 17415 5601 17429 5615
rect 17463 5600 17477 5614
rect 17655 5600 17670 5614
rect 17702 5600 17717 5614
rect 4010 5564 4027 5578
rect 4755 5566 4769 5580
rect 4995 5565 5009 5579
rect 5715 5565 5729 5579
rect 5955 5564 5970 5578
rect 3939 5529 3954 5543
rect 4251 5529 4265 5543
rect 4491 5530 4505 5544
rect 4731 5530 4745 5544
rect 4967 5529 4984 5546
rect 5137 5527 5154 5541
rect 6532 5528 6546 5542
rect 4131 5507 4146 5521
rect 4538 5503 4554 5521
rect 4898 5504 4915 5519
rect 6374 5505 6388 5519
rect 4059 5479 4073 5493
rect 4274 5478 4290 5492
rect 4515 5479 4529 5493
rect 5235 5479 5249 5493
rect 5475 5479 5489 5493
rect 4658 5453 4674 5467
rect 6466 5454 6480 5468
rect 4583 5431 4597 5445
rect 5019 5431 5034 5445
rect 5499 5431 5513 5445
rect 5979 5431 5993 5445
rect 4419 5410 4433 5424
rect 6312 5409 6326 5423
rect 4323 5305 4337 5319
rect 4371 5305 4385 5319
rect 4563 5308 4577 5322
rect 4611 5307 4625 5321
rect 4803 5308 4817 5322
rect 4851 5308 4865 5322
rect 5043 5312 5058 5326
rect 5091 5312 5106 5326
rect 5282 5312 5297 5326
rect 5331 5312 5346 5326
rect 5523 5313 5537 5327
rect 5571 5312 5585 5326
rect 5763 5313 5777 5327
rect 5811 5312 5825 5326
rect 6003 5312 6018 5326
rect 6050 5312 6065 5326
rect 13440 1863 13455 1877
rect 12288 1835 12303 1849
rect 3118 1784 3133 1798
rect 6670 1776 6691 1799
rect 9982 1779 9998 1793
rect 14330 1779 14345 1793
rect 11136 1716 11150 1730
rect 14246 1716 14260 1730
rect 14400 1679 14414 1693
rect 3075 1655 3091 1669
rect 13248 1654 13262 1668
rect 2918 1635 2933 1649
rect 12096 1631 12110 1645
rect 2808 1613 2825 1627
rect 10944 1611 10958 1625
rect 2688 1587 2703 1602
rect 9792 1589 9806 1603
rect 2530 1554 2546 1570
rect 8639 1555 8657 1570
rect 8829 1564 8847 1580
rect 2625 1532 2639 1546
rect 7487 1531 7502 1545
rect 2469 1505 2483 1519
rect 6335 1505 6350 1519
rect 14184 1484 14198 1498
rect 3078 1454 3092 1468
rect 13031 1453 13047 1467
rect 2920 1429 2934 1443
rect 11880 1429 11894 1443
rect 14247 1428 14261 1442
rect 2809 1405 2823 1419
rect 10728 1405 10742 1419
rect 14330 1405 14344 1419
rect 7681 1339 7695 1353
rect 13937 1338 13952 1352
rect 2689 1294 2703 1308
rect 9574 1293 9593 1310
rect 2531 1271 2545 1285
rect 8424 1271 8438 1285
rect 6528 1248 6543 1262
rect 2623 1220 2637 1234
rect 7272 1220 7287 1234
rect 2469 1175 2483 1189
rect 6120 1175 6134 1189
rect 6674 1177 6690 1193
rect 13937 1150 13951 1164
rect 3624 1105 3638 1119
rect 6048 1105 6062 1119
rect 6264 1104 6278 1118
rect 7055 1092 7069 1106
rect 7200 1091 7214 1105
rect 7416 1092 7430 1106
rect 8207 1092 8221 1106
rect 8352 1091 8366 1105
rect 8568 1092 8582 1106
rect 9359 1092 9373 1106
rect 9504 1091 9518 1105
rect 9720 1092 9734 1106
rect 10511 1092 10525 1106
rect 10656 1091 10670 1105
rect 10872 1092 10886 1106
rect 11663 1092 11677 1106
rect 11808 1091 11822 1105
rect 12024 1092 12038 1106
rect 12815 1092 12829 1106
rect 12960 1091 12974 1105
rect 13176 1092 13190 1106
rect 13967 1092 13981 1106
rect 14112 1091 14126 1105
rect 14328 1092 14342 1106
rect 2328 74 2342 88
rect 6191 38 6206 52
rect 7343 38 7358 52
rect 8495 38 8510 52
rect 9648 38 9663 53
rect 10798 38 10816 53
rect 11950 38 11968 53
rect 13102 38 13120 53
rect 14256 37 14270 52
rect 6408 4 6422 18
rect 7560 4 7574 18
rect 8712 4 8726 18
rect 9864 3 9879 18
rect 11015 0 11033 15
rect 12167 0 12185 15
rect 13319 0 13337 15
rect 14472 3 14486 18
<< metal2 >>
rect 10221 6269 10233 6768
rect 3892 5630 3904 6129
rect 3892 5302 3904 5616
rect 4012 5578 4024 6129
rect 3940 5302 3952 5529
rect 4012 5302 4024 5564
rect 4132 5521 4144 6129
rect 10221 5941 10233 6255
rect 10341 6217 10353 6768
rect 10269 5941 10281 6168
rect 10341 5941 10353 6203
rect 10461 6160 10473 6768
rect 10389 5941 10401 6118
rect 10461 5941 10473 6146
rect 10509 5941 10521 6230
rect 10581 5941 10593 6168
rect 10605 5941 10617 6117
rect 10629 5941 10641 6230
rect 10653 5941 10665 5944
rect 10701 5941 10713 5944
rect 10749 5941 10761 6049
rect 10821 5941 10833 6169
rect 10883 6146 10924 6158
rect 10845 5941 10857 6118
rect 10869 5941 10881 6142
rect 10912 6084 10924 6146
rect 10893 5941 10905 5947
rect 10941 5941 10953 5946
rect 10989 5941 11001 6092
rect 11061 5941 11073 6169
rect 11085 5941 11097 6205
rect 11109 5941 11121 6230
rect 11133 5941 11145 5947
rect 11181 5941 11193 5947
rect 11229 5941 11241 6143
rect 11301 5941 11313 6168
rect 11325 5941 11337 6204
rect 11349 5941 11361 6070
rect 11373 5941 11385 5951
rect 11421 5941 11433 5951
rect 11469 5941 11481 6166
rect 11541 5941 11553 6254
rect 11565 5941 11577 6118
rect 11589 5941 11601 6230
rect 11613 5941 11625 5951
rect 11661 5941 11673 5951
rect 11709 5941 11721 6277
rect 11781 5941 11793 6253
rect 11805 5941 11817 6118
rect 11829 5941 11841 6070
rect 11853 5941 11865 5952
rect 11901 5941 11913 5951
rect 11949 5941 11961 6301
rect 12021 5941 12033 6255
rect 12045 5941 12057 6204
rect 12069 5941 12081 6229
rect 12093 5941 12105 5952
rect 12141 5941 12153 5951
rect 12189 5941 12201 6326
rect 12261 5941 12273 6255
rect 12285 5941 12297 6203
rect 12309 5941 12321 6070
rect 12333 5941 12345 5951
rect 12381 5941 12393 5951
rect 12429 5941 12441 6357
rect 12642 6062 12654 6378
rect 12704 6158 12716 6427
rect 12797 6107 12809 6405
rect 12862 6181 12874 6460
rect 12982 6292 12994 6486
rect 13092 6316 13104 6508
rect 15544 5918 15556 6417
rect 4060 5302 4072 5479
rect 4132 5302 4144 5507
rect 4180 5302 4192 5591
rect 4252 5302 4264 5529
rect 4276 5302 4288 5478
rect 4300 5302 4312 5591
rect 4324 5302 4336 5305
rect 4372 5302 4384 5305
rect 4420 5302 4432 5410
rect 4492 5302 4504 5530
rect 4554 5507 4595 5519
rect 4516 5302 4528 5479
rect 4540 5302 4552 5503
rect 4583 5445 4595 5507
rect 4564 5302 4576 5308
rect 4612 5302 4624 5307
rect 4660 5302 4672 5453
rect 4732 5302 4744 5530
rect 4756 5302 4768 5566
rect 4780 5302 4792 5591
rect 4804 5302 4816 5308
rect 4852 5302 4864 5308
rect 4900 5302 4912 5504
rect 4972 5302 4984 5529
rect 4996 5302 5008 5565
rect 5020 5302 5032 5431
rect 5044 5302 5056 5312
rect 5092 5302 5104 5312
rect 5140 5302 5152 5527
rect 5212 5302 5224 5615
rect 5236 5302 5248 5479
rect 5260 5302 5272 5591
rect 5284 5302 5296 5312
rect 5332 5302 5344 5312
rect 5380 5302 5392 5638
rect 5452 5302 5464 5614
rect 5476 5302 5488 5479
rect 5500 5302 5512 5431
rect 5524 5302 5536 5313
rect 5572 5302 5584 5312
rect 5620 5302 5632 5662
rect 5692 5302 5704 5616
rect 5716 5302 5728 5565
rect 5740 5302 5752 5590
rect 5764 5302 5776 5313
rect 5812 5302 5824 5312
rect 5860 5302 5872 5687
rect 5932 5302 5944 5616
rect 5956 5302 5968 5564
rect 5980 5302 5992 5431
rect 6004 5302 6016 5312
rect 6052 5302 6064 5312
rect 6100 5302 6112 5718
rect 6313 5423 6325 5739
rect 6375 5519 6387 5788
rect 6468 5468 6480 5766
rect 6533 5542 6545 5821
rect 6653 5653 6665 5847
rect 6763 5677 6775 5869
rect 15544 5590 15556 5904
rect 15664 5866 15676 6417
rect 15592 5590 15604 5817
rect 15664 5590 15676 5852
rect 15784 5809 15796 6417
rect 15712 5590 15724 5767
rect 15784 5590 15796 5795
rect 15832 5590 15844 5879
rect 15904 5590 15916 5817
rect 15928 5590 15940 5766
rect 15952 5590 15964 5879
rect 15976 5590 15988 5593
rect 16024 5590 16036 5593
rect 16072 5590 16084 5698
rect 16144 5590 16156 5818
rect 16206 5795 16247 5807
rect 16168 5590 16180 5767
rect 16192 5590 16204 5791
rect 16235 5733 16247 5795
rect 16216 5590 16228 5596
rect 16264 5590 16276 5595
rect 16312 5590 16324 5741
rect 16384 5590 16396 5818
rect 16408 5590 16420 5854
rect 16432 5590 16444 5879
rect 16456 5590 16468 5596
rect 16504 5590 16516 5596
rect 16552 5590 16564 5792
rect 16624 5590 16636 5817
rect 16648 5590 16660 5853
rect 16672 5590 16684 5719
rect 16696 5590 16708 5600
rect 16744 5590 16756 5600
rect 16792 5590 16804 5815
rect 16864 5590 16876 5903
rect 16888 5590 16900 5767
rect 16912 5590 16924 5879
rect 16936 5590 16948 5600
rect 16984 5590 16996 5600
rect 17032 5590 17044 5926
rect 17104 5590 17116 5902
rect 17128 5590 17140 5767
rect 17152 5590 17164 5719
rect 17176 5590 17188 5601
rect 17224 5590 17236 5600
rect 17272 5590 17284 5950
rect 17344 5590 17356 5904
rect 17368 5590 17380 5853
rect 17392 5590 17404 5878
rect 17416 5590 17428 5601
rect 17464 5590 17476 5600
rect 17512 5590 17524 5975
rect 17584 5590 17596 5904
rect 17608 5590 17620 5852
rect 17632 5590 17644 5719
rect 17656 5590 17668 5600
rect 17704 5590 17716 5600
rect 17752 5590 17764 6006
rect 17965 5711 17977 6027
rect 18027 5807 18039 6076
rect 18120 5756 18132 6054
rect 18185 5830 18197 6109
rect 18305 5941 18317 6135
rect 18415 5965 18427 6157
rect 12501 5072 12513 5142
rect 17824 4721 17836 4791
rect 6172 4433 6184 4503
rect 3119 1798 3131 1895
rect 2470 1189 2482 1505
rect 2532 1285 2544 1554
rect 2625 1234 2637 1532
rect 2690 1308 2702 1587
rect 2810 1419 2822 1613
rect 2920 1443 2932 1635
rect 3079 1468 3091 1655
rect 3119 1223 3131 1784
rect 3769 1428 3781 1895
rect 3889 1428 3901 1895
rect 4009 1428 4021 1895
rect 3097 1211 3131 1223
rect 3097 1068 3109 1211
rect 3625 1068 3637 1105
rect 6049 1068 6061 1105
rect 6121 1068 6133 1175
rect 6265 1068 6277 1104
rect 6337 1068 6349 1505
rect 6529 1068 6541 1248
rect 6675 1193 6687 1776
rect 7057 1068 7069 1092
rect 7201 1068 7213 1091
rect 7273 1068 7285 1220
rect 7417 1068 7429 1092
rect 7489 1068 7501 1531
rect 7681 1068 7693 1339
rect 8209 1068 8221 1092
rect 8353 1068 8365 1091
rect 8425 1068 8437 1271
rect 8569 1068 8581 1092
rect 8641 1068 8653 1555
rect 8833 1068 8845 1564
rect 9361 1068 9373 1092
rect 9505 1068 9517 1091
rect 9577 1068 9589 1293
rect 9721 1068 9733 1092
rect 9793 1068 9805 1589
rect 9985 1068 9997 1779
rect 10513 1068 10525 1092
rect 10657 1068 10669 1091
rect 10729 1068 10741 1405
rect 10873 1068 10885 1092
rect 10945 1068 10957 1611
rect 11137 1068 11149 1716
rect 11665 1068 11677 1092
rect 11809 1068 11821 1091
rect 11881 1068 11893 1429
rect 12025 1068 12037 1092
rect 12097 1068 12109 1631
rect 12289 1068 12301 1835
rect 12817 1068 12829 1092
rect 12961 1068 12973 1091
rect 13033 1068 13045 1453
rect 13177 1068 13189 1092
rect 13249 1068 13261 1654
rect 13441 1068 13453 1863
rect 13938 1164 13950 1338
rect 13969 1068 13981 1092
rect 14113 1068 14125 1091
rect 14185 1068 14197 1484
rect 14247 1442 14259 1716
rect 14331 1419 14343 1779
rect 14329 1068 14341 1092
rect 14401 1068 14413 1679
rect 2329 88 2341 269
rect 6193 52 6205 269
rect 6409 18 6421 269
rect 7345 52 7357 269
rect 7561 18 7573 269
rect 8497 52 8509 269
rect 8713 18 8725 269
rect 9649 53 9661 269
rect 9865 18 9877 269
rect 10801 53 10813 269
rect 11017 15 11029 269
rect 11953 53 11965 269
rect 12169 15 12181 269
rect 13105 53 13117 269
rect 13321 15 13333 269
rect 14257 52 14269 269
rect 14473 18 14485 269
use inv inv_33
timestamp 1386238110
transform 1 0 3868 0 1 4503
box 0 0 120 799
use inv inv_34
timestamp 1386238110
transform 1 0 3988 0 1 4503
box 0 0 120 799
use inv inv_35
timestamp 1386238110
transform 1 0 4108 0 1 4503
box 0 0 120 799
use nand3 nand3_24
timestamp 1386234893
transform 1 0 4228 0 1 4503
box 0 0 120 799
use inv inv_36
timestamp 1386238110
transform 1 0 4348 0 1 4503
box 0 0 120 799
use nand3 nand3_25
timestamp 1386234893
transform 1 0 4468 0 1 4503
box 0 0 120 799
use inv inv_37
timestamp 1386238110
transform 1 0 4588 0 1 4503
box 0 0 120 799
use nand3 nand3_26
timestamp 1386234893
transform 1 0 4708 0 1 4503
box 0 0 120 799
use inv inv_38
timestamp 1386238110
transform 1 0 4828 0 1 4503
box 0 0 120 799
use nand3 nand3_27
timestamp 1386234893
transform 1 0 4948 0 1 4503
box 0 0 120 799
use inv inv_39
timestamp 1386238110
transform 1 0 5068 0 1 4503
box 0 0 120 799
use nand3 nand3_28
timestamp 1386234893
transform 1 0 5188 0 1 4503
box 0 0 120 799
use inv inv_40
timestamp 1386238110
transform 1 0 5308 0 1 4503
box 0 0 120 799
use nand3 nand3_29
timestamp 1386234893
transform 1 0 5428 0 1 4503
box 0 0 120 799
use inv inv_41
timestamp 1386238110
transform 1 0 5548 0 1 4503
box 0 0 120 799
use nand3 nand3_30
timestamp 1386234893
transform 1 0 5668 0 1 4503
box 0 0 120 799
use inv inv_42
timestamp 1386238110
transform 1 0 5788 0 1 4503
box 0 0 120 799
use nand3 nand3_31
timestamp 1386234893
transform 1 0 5908 0 1 4503
box 0 0 120 799
use inv inv_43
timestamp 1386238110
transform 1 0 6028 0 1 4503
box 0 0 120 799
use inv inv_44
timestamp 1386238110
transform 1 0 10197 0 1 5142
box 0 0 120 799
use inv inv_45
timestamp 1386238110
transform 1 0 10317 0 1 5142
box 0 0 120 799
use inv inv_46
timestamp 1386238110
transform 1 0 10437 0 1 5142
box 0 0 120 799
use nand3 nand3_32
timestamp 1386234893
transform 1 0 10557 0 1 5142
box 0 0 120 799
use inv inv_47
timestamp 1386238110
transform 1 0 10677 0 1 5142
box 0 0 120 799
use nand3 nand3_33
timestamp 1386234893
transform 1 0 10797 0 1 5142
box 0 0 120 799
use inv inv_48
timestamp 1386238110
transform 1 0 10917 0 1 5142
box 0 0 120 799
use nand3 nand3_34
timestamp 1386234893
transform 1 0 11037 0 1 5142
box 0 0 120 799
use inv inv_49
timestamp 1386238110
transform 1 0 11157 0 1 5142
box 0 0 120 799
use nand3 nand3_35
timestamp 1386234893
transform 1 0 11277 0 1 5142
box 0 0 120 799
use inv inv_50
timestamp 1386238110
transform 1 0 11397 0 1 5142
box 0 0 120 799
use nand3 nand3_36
timestamp 1386234893
transform 1 0 11517 0 1 5142
box 0 0 120 799
use inv inv_51
timestamp 1386238110
transform 1 0 11637 0 1 5142
box 0 0 120 799
use nand3 nand3_37
timestamp 1386234893
transform 1 0 11757 0 1 5142
box 0 0 120 799
use inv inv_52
timestamp 1386238110
transform 1 0 11877 0 1 5142
box 0 0 120 799
use nand3 nand3_38
timestamp 1386234893
transform 1 0 11997 0 1 5142
box 0 0 120 799
use inv inv_53
timestamp 1386238110
transform 1 0 12117 0 1 5142
box 0 0 120 799
use nand3 nand3_39
timestamp 1386234893
transform 1 0 12237 0 1 5142
box 0 0 120 799
use inv inv_54
timestamp 1386238110
transform 1 0 12357 0 1 5142
box 0 0 120 799
use inv inv_55
timestamp 1386238110
transform 1 0 15520 0 1 4791
box 0 0 120 799
use inv inv_56
timestamp 1386238110
transform 1 0 15640 0 1 4791
box 0 0 120 799
use inv inv_57
timestamp 1386238110
transform 1 0 15760 0 1 4791
box 0 0 120 799
use nand3 nand3_40
timestamp 1386234893
transform 1 0 15880 0 1 4791
box 0 0 120 799
use inv inv_58
timestamp 1386238110
transform 1 0 16000 0 1 4791
box 0 0 120 799
use nand3 nand3_41
timestamp 1386234893
transform 1 0 16120 0 1 4791
box 0 0 120 799
use inv inv_59
timestamp 1386238110
transform 1 0 16240 0 1 4791
box 0 0 120 799
use nand3 nand3_42
timestamp 1386234893
transform 1 0 16360 0 1 4791
box 0 0 120 799
use inv inv_60
timestamp 1386238110
transform 1 0 16480 0 1 4791
box 0 0 120 799
use nand3 nand3_43
timestamp 1386234893
transform 1 0 16600 0 1 4791
box 0 0 120 799
use inv inv_61
timestamp 1386238110
transform 1 0 16720 0 1 4791
box 0 0 120 799
use nand3 nand3_44
timestamp 1386234893
transform 1 0 16840 0 1 4791
box 0 0 120 799
use inv inv_62
timestamp 1386238110
transform 1 0 16960 0 1 4791
box 0 0 120 799
use nand3 nand3_45
timestamp 1386234893
transform 1 0 17080 0 1 4791
box 0 0 120 799
use inv inv_63
timestamp 1386238110
transform 1 0 17200 0 1 4791
box 0 0 120 799
use nand3 nand3_46
timestamp 1386234893
transform 1 0 17320 0 1 4791
box 0 0 120 799
use inv inv_64
timestamp 1386238110
transform 1 0 17440 0 1 4791
box 0 0 120 799
use nand3 nand3_47
timestamp 1386234893
transform 1 0 17560 0 1 4791
box 0 0 120 799
use inv inv_65
timestamp 1386238110
transform 1 0 17680 0 1 4791
box 0 0 120 799
use scanreg scanreg_1
timestamp 1386241447
transform 1 0 3025 0 1 269
box 0 0 720 799
use trisbuf trisbuf_0
timestamp 1386237216
transform 1 0 6025 0 1 269
box 0 0 216 799
use trisbuf trisbuf_1
timestamp 1386237216
transform 1 0 6241 0 1 269
box 0 0 216 799
use scanreg scanreg_2
timestamp 1386241447
transform 1 0 6457 0 1 269
box 0 0 720 799
use trisbuf trisbuf_2
timestamp 1386237216
transform 1 0 7177 0 1 269
box 0 0 216 799
use trisbuf trisbuf_3
timestamp 1386237216
transform 1 0 7393 0 1 269
box 0 0 216 799
use scanreg scanreg_3
timestamp 1386241447
transform 1 0 7609 0 1 269
box 0 0 720 799
use trisbuf trisbuf_4
timestamp 1386237216
transform 1 0 8329 0 1 269
box 0 0 216 799
use trisbuf trisbuf_5
timestamp 1386237216
transform 1 0 8545 0 1 269
box 0 0 216 799
use scanreg scanreg_4
timestamp 1386241447
transform 1 0 8761 0 1 269
box 0 0 720 799
use trisbuf trisbuf_6
timestamp 1386237216
transform 1 0 9481 0 1 269
box 0 0 216 799
use trisbuf trisbuf_7
timestamp 1386237216
transform 1 0 9697 0 1 269
box 0 0 216 799
use scanreg scanreg_5
timestamp 1386241447
transform 1 0 9913 0 1 269
box 0 0 720 799
use trisbuf trisbuf_8
timestamp 1386237216
transform 1 0 10633 0 1 269
box 0 0 216 799
use trisbuf trisbuf_9
timestamp 1386237216
transform 1 0 10849 0 1 269
box 0 0 216 799
use scanreg scanreg_6
timestamp 1386241447
transform 1 0 11065 0 1 269
box 0 0 720 799
use trisbuf trisbuf_10
timestamp 1386237216
transform 1 0 11785 0 1 269
box 0 0 216 799
use trisbuf trisbuf_11
timestamp 1386237216
transform 1 0 12001 0 1 269
box 0 0 216 799
use scanreg scanreg_7
timestamp 1386241447
transform 1 0 12217 0 1 269
box 0 0 720 799
use trisbuf trisbuf_12
timestamp 1386237216
transform 1 0 12937 0 1 269
box 0 0 216 799
use trisbuf trisbuf_13
timestamp 1386237216
transform 1 0 13153 0 1 269
box 0 0 216 799
use scanreg scanreg_8
timestamp 1386241447
transform 1 0 13369 0 1 269
box 0 0 720 799
use trisbuf trisbuf_14
timestamp 1386237216
transform 1 0 14089 0 1 269
box 0 0 216 799
use trisbuf trisbuf_15
timestamp 1386237216
transform 1 0 14305 0 1 269
box 0 0 216 799
<< labels >>
rlabel metal2 3769 1895 3781 1895 5 Rs1[0]
rlabel metal2 3889 1895 3901 1895 5 Rs1[1]
rlabel metal2 4009 1895 4021 1895 5 Rs1[2]
rlabel metal2 3119 1895 3131 1895 5 WData[0]
rlabel metal1 0 75 0 85 3 Databus
rlabel metal1 0 40 0 50 3 Rd1[0]
rlabel metal1 0 5 0 15 3 Rd2[0]
rlabel metal1 16815 75 16815 85 7 Databus
rlabel metal1 16815 40 16815 50 7 Rd1[0]
rlabel metal1 16815 5 16815 15 7 Rd2[0]
rlabel metal2 10221 6768 10233 6768 5 Rs2[0]
rlabel metal2 10341 6768 10353 6768 5 Rs2[1]
rlabel metal2 10461 6768 10473 6768 5 Rs2[2]
rlabel metal1 10172 5863 10172 5888 3 Vdd!
rlabel metal1 10172 5218 10172 5243 3 GND!
rlabel metal1 10172 5195 10172 5205 3 Clock
rlabel metal1 10172 5149 10172 5159 3 nReset
rlabel metal2 15544 6417 15556 6417 5 Rs2[0]
rlabel metal2 15664 6417 15676 6417 5 Rs2[1]
rlabel metal2 15784 6417 15796 6417 5 Rs2[2]
rlabel metal1 15495 5512 15495 5537 3 Vdd!
rlabel metal1 15495 4867 15495 4892 3 GND!
rlabel metal1 15495 4844 15495 4854 3 Clock
rlabel metal1 15495 4798 15495 4808 3 nReset
rlabel metal2 3892 6129 3904 6129 5 Rs2[0]
rlabel metal2 4012 6129 4024 6129 5 Rs2[1]
rlabel metal2 4132 6129 4144 6129 5 Rs2[2]
rlabel metal1 3843 5224 3843 5249 3 Vdd!
rlabel metal1 3843 4579 3843 4604 3 GND!
rlabel metal1 3843 4556 3843 4566 3 Clock
rlabel metal1 3843 4510 3843 4520 3 nReset
<< end >>
