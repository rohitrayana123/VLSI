magic
tech c035u
timestamp 1394833348
<< checkpaint >>
rect 11084 3405 17801 3898
rect 4724 771 17801 3405
rect 4724 -813 16540 771
<< nwell >>
rect 1416 1428 3432 1826
rect 15240 1428 15864 1826
rect 23518 1428 24288 1826
<< pwell >>
rect 1416 1027 3432 1428
rect 15240 1034 15864 1428
rect 23518 1027 24288 1428
<< pohmic >>
rect 1416 1103 1422 1113
rect 3426 1103 3432 1113
rect 15240 1103 15246 1113
rect 15858 1103 15864 1113
rect 23518 1103 23524 1113
rect 24282 1103 24288 1113
<< nohmic >>
rect 1416 1763 1422 1773
rect 3426 1763 3432 1773
rect 15240 1763 15246 1773
rect 15858 1763 15864 1773
rect 23518 1763 23524 1773
rect 24282 1763 24288 1773
<< psubstratetap >>
rect 1422 1103 3426 1119
rect 15246 1103 15858 1119
rect 23524 1103 24282 1119
<< nsubstratetap >>
rect 1422 1757 3426 1773
rect 15246 1757 15858 1773
rect 23524 1757 24282 1773
<< metal1 >>
rect 3829 2221 6359 2231
rect 13453 2227 16487 2237
rect 4261 2199 6335 2209
rect 13261 2205 16367 2215
rect 4693 2177 6311 2187
rect 13069 2183 16247 2193
rect 5125 2154 6095 2164
rect 12877 2161 16127 2171
rect 5557 2133 6071 2143
rect 12685 2139 16007 2149
rect 5989 2111 6047 2121
rect 12493 2117 15887 2127
rect 4381 2007 5711 2017
rect 4429 1985 5663 1995
rect 3997 1963 5231 1973
rect 3949 1941 5279 1951
rect 3564 1919 4799 1929
rect 3517 1897 4847 1907
rect 3493 1875 3911 1885
rect 3925 1875 4343 1885
rect 4789 1875 5207 1885
rect 5221 1875 5639 1885
rect 3733 1853 4151 1863
rect 4165 1853 4583 1863
rect 5029 1853 5447 1863
rect 5461 1853 5879 1863
rect 3589 1831 3743 1841
rect 4021 1831 4175 1841
rect 4453 1831 4607 1841
rect 4885 1831 5039 1841
rect 5317 1831 5471 1841
rect 5749 1831 5903 1841
rect 1416 1809 3432 1819
rect 15240 1809 15864 1819
rect 23518 1809 24288 1819
rect 1416 1786 3432 1796
rect 15240 1786 15864 1796
rect 23518 1786 24288 1796
rect 1416 1757 1422 1773
rect 3426 1757 3432 1773
rect 1416 1748 3432 1757
rect 15240 1757 15246 1773
rect 15858 1757 15864 1773
rect 15240 1748 15864 1757
rect 23518 1757 23524 1773
rect 24282 1757 24288 1773
rect 23518 1748 24288 1757
rect 1416 1119 3432 1128
rect 1416 1103 1422 1119
rect 3426 1103 3432 1119
rect 15240 1119 15864 1128
rect 15240 1103 15246 1119
rect 15858 1103 15864 1119
rect 23518 1119 24288 1128
rect 23518 1103 23524 1119
rect 24282 1103 24288 1119
rect 1416 1080 3432 1090
rect 15240 1080 15864 1090
rect 1416 1057 3432 1067
rect 15240 1057 15864 1067
rect 1416 1034 3432 1044
rect 15240 1034 15864 1044
rect 21301 28 21335 38
rect 21349 28 21383 38
rect 21397 28 21431 38
rect 21445 28 21479 38
rect 21493 28 21527 38
rect 21541 28 21575 38
rect 21589 28 21623 38
rect 21637 28 21935 38
rect 21949 28 21983 38
rect 21997 28 22031 38
rect 22045 28 22079 38
rect 22093 28 22391 38
rect 22405 28 22439 38
rect 22453 28 22751 38
<< m2contact >>
rect 3815 2219 3829 2233
rect 6359 2219 6373 2233
rect 13439 2226 13453 2240
rect 16487 2225 16501 2239
rect 4247 2197 4261 2211
rect 6335 2197 6349 2211
rect 13247 2203 13261 2217
rect 16367 2203 16381 2217
rect 4679 2175 4693 2189
rect 6311 2175 6325 2189
rect 13055 2181 13069 2195
rect 16247 2181 16261 2195
rect 5111 2152 5125 2166
rect 6095 2152 6109 2166
rect 12863 2159 12877 2173
rect 16127 2159 16141 2173
rect 5543 2130 5557 2144
rect 6071 2130 6085 2144
rect 12671 2137 12685 2151
rect 16007 2137 16021 2151
rect 5975 2109 5989 2123
rect 6047 2108 6061 2122
rect 12479 2115 12493 2129
rect 15887 2115 15901 2129
rect 4367 2005 4381 2019
rect 5711 2005 5725 2019
rect 4415 1983 4429 1997
rect 5663 1983 5677 1997
rect 3983 1961 3997 1975
rect 5231 1961 5245 1975
rect 3935 1939 3949 1953
rect 5279 1939 5293 1953
rect 3550 1917 3564 1931
rect 4799 1917 4813 1931
rect 3503 1895 3517 1909
rect 4847 1895 4861 1909
rect 3479 1873 3493 1887
rect 3911 1873 3925 1887
rect 4343 1873 4357 1887
rect 4775 1873 4789 1887
rect 5207 1873 5221 1887
rect 5639 1873 5653 1887
rect 3719 1851 3733 1865
rect 4151 1851 4165 1865
rect 4583 1851 4597 1865
rect 5015 1851 5029 1865
rect 5447 1851 5461 1865
rect 5879 1851 5893 1865
rect 3575 1829 3589 1843
rect 3743 1829 3757 1843
rect 4007 1829 4021 1843
rect 4175 1829 4189 1843
rect 4439 1829 4453 1843
rect 4607 1829 4621 1843
rect 4871 1829 4885 1843
rect 5039 1829 5053 1843
rect 5303 1829 5317 1843
rect 5471 1829 5485 1843
rect 5735 1829 5749 1843
rect 5903 1829 5917 1843
rect 21287 26 21301 40
rect 21335 26 21349 40
rect 21383 26 21397 40
rect 21431 26 21445 40
rect 21479 26 21493 40
rect 21527 26 21541 40
rect 21575 26 21589 40
rect 21623 26 21637 40
rect 21935 25 21949 39
rect 21983 25 21997 39
rect 22031 25 22045 39
rect 22079 25 22093 39
rect 22391 26 22405 40
rect 22439 26 22453 40
rect 22751 26 22765 40
<< metal2 >>
rect -48 1826 152 2783
rect 168 1826 180 2783
rect 192 1826 204 2783
rect 216 1826 228 2783
rect 240 1826 252 2783
rect 3480 1887 3492 2783
rect 3504 1909 3516 2783
rect 3552 1931 3564 2783
rect 3480 1826 3492 1873
rect 3504 1826 3516 1895
rect 3552 1826 3564 1917
rect 3720 1865 3732 2783
rect 3576 1826 3588 1829
rect 3720 1826 3732 1851
rect 3744 1826 3756 1829
rect 3816 1826 3828 2219
rect 3936 1953 3948 2783
rect 3984 1975 3996 2783
rect 3912 1826 3924 1873
rect 3936 1826 3948 1939
rect 3984 1826 3996 1961
rect 4008 1826 4020 1829
rect 4152 1826 4164 1851
rect 4176 1826 4188 1829
rect 4248 1826 4260 2197
rect 4368 2019 4380 2783
rect 4344 1826 4356 1873
rect 4368 1826 4380 2005
rect 4416 1997 4428 2783
rect 4416 1826 4428 1983
rect 4440 1826 4452 1829
rect 4584 1826 4596 1851
rect 4608 1826 4620 1829
rect 4680 1826 4692 2175
rect 4776 1887 4788 2783
rect 4776 1826 4788 1873
rect 4800 1826 4812 1917
rect 4848 1826 4860 1895
rect 5016 1865 5028 2783
rect 4872 1826 4884 1829
rect 5016 1826 5028 1851
rect 5040 1826 5052 1829
rect 5112 1826 5124 2152
rect 5208 1826 5220 1873
rect 5232 1826 5244 1961
rect 5280 1826 5292 1939
rect 5304 1826 5316 1829
rect 5448 1826 5460 1851
rect 5472 1826 5484 1829
rect 5544 1826 5556 2130
rect 5640 1826 5652 1873
rect 5664 1826 5676 1983
rect 5712 1826 5724 2005
rect 5736 1826 5748 1829
rect 5880 1826 5892 1851
rect 5904 1826 5916 1829
rect 5976 1826 5988 2109
rect 6048 2105 6060 2108
rect 6072 2105 6084 2130
rect 6096 2105 6108 2152
rect 6146 2105 6158 2783
rect 6312 2105 6324 2175
rect 6336 2105 6348 2197
rect 6360 2105 6372 2219
rect 6456 2105 6468 2783
rect 6480 2105 6492 2783
rect 6504 2105 6516 2783
rect 12384 2105 12396 2783
rect 12408 2105 12420 2783
rect 12480 2105 12492 2115
rect 12600 2105 12612 2783
rect 12648 2105 12660 2783
rect 12672 2105 12684 2137
rect 12792 2105 12804 2783
rect 12864 2105 12876 2159
rect 12984 2105 12996 2783
rect 13056 2105 13068 2181
rect 13176 2105 13188 2783
rect 13248 2105 13260 2203
rect 13368 2105 13380 2783
rect 13440 2105 13452 2226
rect 15888 1999 15900 2115
rect 16008 1997 16020 2137
rect 16128 2002 16140 2159
rect 16248 2002 16260 2181
rect 16368 2002 16380 2203
rect 16488 2001 16500 2225
rect 16920 2002 16932 2783
rect 17112 2002 17124 2783
rect 17184 2002 17196 2783
rect 17280 2002 17292 2783
rect 21936 2002 21948 2783
rect 22128 2002 22140 2783
rect 22248 2002 22260 2783
rect 22368 2002 22380 2783
rect 24408 1826 24608 2783
rect -48 0 152 1027
rect 168 0 180 1027
rect 192 0 204 1027
rect 216 0 228 1027
rect 240 0 252 1027
rect 3648 1017 3660 1027
rect 3792 1017 3804 1027
rect 3648 1005 3804 1017
rect 4080 1017 4092 1027
rect 4224 1017 4236 1027
rect 4080 1005 4236 1017
rect 4512 1017 4524 1027
rect 4656 1017 4668 1027
rect 4512 1005 4668 1017
rect 4944 1017 4956 1027
rect 5088 1017 5100 1027
rect 4944 1005 5100 1017
rect 5376 1017 5388 1027
rect 5520 1017 5532 1027
rect 5376 1005 5532 1017
rect 5808 1017 5820 1027
rect 5952 1017 5964 1027
rect 5808 1005 5964 1017
rect 6096 0 6108 487
rect 6840 0 6852 487
rect 7056 0 7068 487
rect 7248 0 7260 487
rect 7992 0 8004 487
rect 8208 0 8220 487
rect 8400 0 8412 487
rect 9144 0 9156 487
rect 9360 0 9372 487
rect 9552 0 9564 487
rect 10296 0 10308 487
rect 10512 0 10524 487
rect 10704 0 10716 487
rect 11448 0 11460 487
rect 11664 0 11676 487
rect 11856 0 11868 487
rect 12600 0 12612 487
rect 12816 0 12828 487
rect 13008 0 13020 487
rect 13752 0 13764 487
rect 13968 0 13980 487
rect 14160 0 14172 487
rect 14904 0 14916 487
rect 15120 0 15132 487
rect 15936 0 15948 763
rect 16200 0 16212 763
rect 16368 0 16380 763
rect 16536 0 16548 763
rect 16560 0 16572 763
rect 16632 0 16644 763
rect 16848 0 16860 763
rect 16992 0 17004 763
rect 17328 0 17340 763
rect 17688 0 17700 763
rect 18096 0 18108 763
rect 18432 0 18444 763
rect 18744 0 18756 763
rect 19080 0 19092 763
rect 19200 0 19212 763
rect 19248 0 19260 763
rect 19416 0 19428 763
rect 21216 0 21228 763
rect 21241 0 21253 763
rect 21528 40 21540 763
rect 21288 0 21300 26
rect 21336 0 21348 26
rect 21384 0 21396 26
rect 21432 0 21444 26
rect 21480 0 21492 26
rect 21528 0 21540 26
rect 21576 0 21588 26
rect 21624 0 21636 26
rect 21864 0 21876 763
rect 21936 0 21948 25
rect 21984 0 21996 25
rect 22032 0 22044 25
rect 22080 0 22092 25
rect 22320 0 22332 763
rect 22392 0 22404 26
rect 22440 0 22452 26
rect 22680 0 22692 763
rect 22752 0 22764 26
rect 23040 0 23052 763
rect 23208 0 23220 763
rect 23448 73 23460 763
rect 23448 61 24180 73
rect 24168 0 24180 61
rect 24408 0 24608 1027
use leftbuf  leftbuf_1
timestamp 1386242881
transform 1 0 -48 0 1 1027
box 0 0 1464 799
use mux2  mux2_6
timestamp 1386235218
transform 1 0 3432 0 1 1027
box 0 0 192 799
use tiehigh  tiehigh_3
timestamp 1386086759
transform 1 0 3624 0 1 1027
box 0 0 48 799
use mux2  mux2_7
timestamp 1386235218
transform 1 0 3672 0 1 1027
box 0 0 192 799
use mux2  mux2_8
timestamp 1386235218
transform 1 0 3864 0 1 1027
box 0 0 192 799
use tiehigh  tiehigh_4
timestamp 1386086759
transform 1 0 4056 0 1 1027
box 0 0 48 799
use mux2  mux2_9
timestamp 1386235218
transform 1 0 4104 0 1 1027
box 0 0 192 799
use mux2  mux2_10
timestamp 1386235218
transform 1 0 4296 0 1 1027
box 0 0 192 799
use tiehigh  tiehigh_5
timestamp 1386086759
transform 1 0 4488 0 1 1027
box 0 0 48 799
use mux2  mux2_11
timestamp 1386235218
transform 1 0 4536 0 1 1027
box 0 0 192 799
use mux2  mux2_4
timestamp 1386235218
transform 1 0 4728 0 1 1027
box 0 0 192 799
use tiehigh  tiehigh_2
timestamp 1386086759
transform 1 0 4920 0 1 1027
box 0 0 48 799
use mux2  mux2_5
timestamp 1386235218
transform 1 0 4968 0 1 1027
box 0 0 192 799
use mux2  mux2_2
timestamp 1386235218
transform 1 0 5160 0 1 1027
box 0 0 192 799
use tiehigh  tiehigh_1
timestamp 1386086759
transform 1 0 5352 0 1 1027
box 0 0 48 799
use mux2  mux2_3
timestamp 1386235218
transform 1 0 5400 0 1 1027
box 0 0 192 799
use mux2  mux2_1
timestamp 1386235218
transform 1 0 5592 0 1 1027
box 0 0 192 799
use tiehigh  tiehigh_0
timestamp 1386086759
transform 1 0 5784 0 1 1027
box 0 0 48 799
use mux2  mux2_0
timestamp 1386235218
transform 1 0 5832 0 1 1027
box 0 0 192 799
use regBlock_decoder  regBlock_decoder_0
timestamp 1394802642
transform 1 0 6024 0 1 487
box 0 0 9216 1618
use ALUDecoder_new  ALUDecoder_new_0
timestamp 1394755051
transform 1 0 15864 0 1 763
box 0 0 7654 1239
use rightend  rightend_0
timestamp 1386235834
transform 1 0 24288 0 1 1027
box 0 0 320 799
<< labels >>
rlabel metal2 21216 0 21228 0 1 Sh8
rlabel metal2 16632 0 16644 0 1 Flags[3]
rlabel metal2 15936 0 15948 0 1 ZeroA
rlabel metal2 23208 0 23220 0 1 LLI
rlabel metal2 23040 0 23052 0 1 ShOut
rlabel metal2 22320 0 22332 0 1 Sh2
rlabel metal2 21241 0 21253 0 1 ShR
rlabel metal2 22680 0 22692 0 1 Sh1
rlabel metal2 21864 0 21876 0 1 Sh4
rlabel metal2 19080 0 19092 0 1 NOR
rlabel metal2 19248 0 19260 0 1 ShB
rlabel metal2 19200 0 19212 0 1 ASign
rlabel metal2 19416 0 19428 0 1 ShL
rlabel metal2 18432 0 18444 0 1 NOT
rlabel metal2 18096 0 18108 0 1 XOR
rlabel metal2 17688 0 17700 0 1 OR
rlabel metal2 17328 0 17340 0 1 AND
rlabel metal2 16992 0 17004 0 1 FAOut
rlabel metal2 16848 0 16860 0 1 nZ
rlabel metal2 16560 0 16572 0 1 COut
rlabel metal2 16536 0 16548 0 1 LastCIn
rlabel metal2 16368 0 16380 0 1 CIn_slice
rlabel metal2 16200 0 16212 0 1 SUB
rlabel metal2 18744 0 18756 0 1 NAND
rlabel metal2 21576 0 21588 0 5 Sh8G_R
rlabel metal2 21528 0 21540 0 5 Sh8F_R
rlabel metal2 21480 0 21492 0 5 Sh8E_R
rlabel metal2 21432 0 21444 0 5 Sh8D_R
rlabel metal2 21288 0 21300 0 5 Sh8A_R
rlabel metal2 21336 0 21348 0 5 Sh8B_R
rlabel metal2 21384 0 21396 0 5 Sh8C_R
rlabel metal2 21624 0 21636 0 5 Sh8H_R
rlabel metal2 21984 0 21996 0 5 Sh4A_R
rlabel metal2 22032 0 22044 0 5 Sh4B_R
rlabel metal2 22080 0 22092 0 5 Sh4C_R
rlabel metal2 21936 0 21948 0 5 Sh4Z_R
rlabel metal2 22392 0 22404 0 5 Sh2A_R
rlabel metal2 22440 0 22452 0 5 Sh2B_R
rlabel metal2 22752 0 22764 0 1 Sh1_R_In
rlabel metal2 24168 0 24180 0 1 OutEn
rlabel metal2 24410 0 24608 0 1 GND!
rlabel metal2 5016 2783 5028 2783 5 RwSel[1]
rlabel metal2 4368 2783 4380 2783 5 Ir[8]
rlabel metal2 4416 2783 4428 2783 5 Ir[5]
rlabel metal2 3984 2783 3996 2783 5 Ir[6]
rlabel metal2 3936 2783 3948 2783 5 Ir[9]
rlabel metal2 3552 2783 3564 2783 5 Ir[7]
rlabel metal2 3504 2783 3516 2783 5 Ir[10]
rlabel metal2 3720 2783 3732 2783 5 Rs1Sel[1]
rlabel metal2 3480 2783 3492 2783 5 Rs1Sel[0]
rlabel metal2 6146 2783 6158 2783 5 RegWe
rlabel metal2 6504 2783 6516 2783 5 Ir[4]
rlabel metal2 6480 2783 6492 2783 5 Ir[3]
rlabel metal2 6456 2783 6468 2783 5 Ir[2]
rlabel metal2 4776 2783 4788 2783 5 RwSel[0]
rlabel metal2 6096 0 6108 0 1 Rw[0]
rlabel metal2 6840 0 6852 0 1 Rs1[0]
rlabel metal2 7056 0 7068 0 1 Rs2[0]
rlabel metal2 8208 0 8220 0 1 Rs2[1]
rlabel metal2 8400 0 8412 0 1 Rw[2]
rlabel metal2 9144 0 9156 0 1 Rs1[2]
rlabel metal2 9360 0 9372 0 1 Rs2[2]
rlabel metal2 9552 0 9564 0 1 Rw[3]
rlabel metal2 10296 0 10308 0 1 Rs1[3]
rlabel metal2 10704 0 10716 0 1 Rw[4]
rlabel metal2 11448 0 11460 0 1 Rs1[4]
rlabel metal2 11664 0 11676 0 1 Rs2[4]
rlabel metal2 11856 0 11868 0 1 Rw[5]
rlabel metal2 12600 0 12612 0 1 Rs1[5]
rlabel metal2 12816 0 12828 0 1 Rs2[5]
rlabel metal2 13008 0 13020 0 1 Rw[6]
rlabel metal2 13752 0 13764 0 1 Rs1[6]
rlabel metal2 13968 0 13980 0 1 Rs2[6]
rlabel metal2 14160 0 14172 0 1 Rw[7]
rlabel metal2 14904 0 14916 0 1 Rs1[7]
rlabel metal2 15120 0 15132 0 1 Rs2[7]
rlabel metal2 7248 0 7260 0 1 Rw[1]
rlabel metal2 7992 0 8004 0 1 Rs1[1]
rlabel metal2 10512 0 10524 0 1 Rs2[3]
rlabel metal1 6021 2116 6021 2116 1 Rw0
rlabel metal1 6020 2137 6020 2137 1 Rw1
rlabel metal1 6014 2159 6014 2159 1 Rw2
rlabel metal1 6016 2181 6016 2181 1 Rs10
rlabel metal1 6016 2204 6016 2204 1 Rs11
rlabel metal1 6017 2224 6017 2224 1 Rs12
rlabel metal2 192 2783 204 2783 1 Test
rlabel metal2 216 2783 228 2783 1 Clock
rlabel metal2 240 2783 252 2783 1 nReset
rlabel metal2 -48 2783 152 2783 5 Vdd!
rlabel metal2 168 2783 180 2783 5 SDO
rlabel metal2 168 0 180 0 1 SDI
rlabel metal2 192 0 204 0 1 Test
rlabel metal2 216 0 228 0 1 Clock
rlabel metal2 240 0 252 0 1 nReset
rlabel metal2 -48 0 152 0 1 Vdd!
rlabel metal2 24408 2783 24608 2783 1 GND!
rlabel metal2 17280 2783 17292 2783 5 Flagss[0]
rlabel metal2 17184 2783 17196 2783 5 Flags[3]
rlabel metal2 17112 2783 17124 2783 5 Flags[1]
rlabel metal2 16920 2783 16932 2783 5 Flags[2]
rlabel metal2 21936 2783 21948 2783 5 Ir[3]
rlabel metal2 22128 2783 22140 2783 5 Ir[2]
rlabel metal2 22248 2783 22260 2783 5 Ir[1]
rlabel metal2 22368 2783 22380 2783 5 Ir[0]
rlabel metal2 12384 2783 12396 2783 1 AluOR[1]
rlabel metal2 12408 2783 12420 2783 5 Ir[15]
rlabel metal2 12600 2783 12612 2783 5 Ir[14]
rlabel metal2 12648 2783 12660 2783 1 AluOR[0]
rlabel metal2 12792 2783 12804 2783 5 Ir[13]
rlabel metal2 12984 2783 12996 2783 5 Ir[12]
rlabel metal2 13176 2783 13188 2783 5 Ir[11]
rlabel metal2 13368 2783 13380 2783 5 Cin
<< end >>
