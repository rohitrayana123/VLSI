../../../Design/Implementation/verilog/behavioural/demux_bus.sv