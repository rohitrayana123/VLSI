../../../Design/Implementation/verilog/behavioural/system.sv