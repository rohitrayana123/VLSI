magic
tech c035u
timestamp 1395422108
<< nwell >>
rect 27435 1534 27795 1932
<< pwell >>
rect 27435 1133 27795 1534
<< metal1 >>
rect 18832 8777 24734 8787
rect 16936 8753 23198 8763
rect 13384 8729 20126 8739
rect 13048 8705 17054 8715
rect 18688 8705 27842 8715
rect 12256 8679 12274 8693
rect 12688 8681 21662 8691
rect 7144 8655 7162 8669
rect 10864 8657 18866 8667
rect 20116 8657 23834 8667
rect 84 8633 25778 8643
rect 84 8609 1706 8619
rect 2872 8609 4694 8619
rect 6952 8609 27866 8619
rect 84 8585 1754 8595
rect 3124 8585 9218 8595
rect 10360 8585 27818 8595
rect 27856 8585 28227 8595
rect 4672 8561 7826 8571
rect 8752 8559 8770 8573
rect 11104 8561 26270 8571
rect 27736 8561 28227 8571
rect 7096 8537 27842 8547
rect 27880 8537 28227 8547
rect 13960 8513 23186 8523
rect 27784 8513 27794 8523
rect 27856 8513 28227 8523
rect 15508 8489 25562 8499
rect 27808 8489 28227 8499
rect 16840 8465 27794 8475
rect 27832 8465 28227 8475
rect 17044 8441 22850 8451
rect 27808 8441 28227 8451
rect 13120 7608 13778 7618
rect 12208 7584 12962 7594
rect 13096 7584 13250 7594
rect 13840 7584 21362 7594
rect 12112 7560 12650 7570
rect 12784 7560 15890 7570
rect 11800 7536 24266 7546
rect 11728 7512 24362 7522
rect 11656 7488 23426 7498
rect 25576 7488 25778 7498
rect 11272 7464 11306 7474
rect 11584 7464 11786 7474
rect 11896 7464 25562 7474
rect 11248 7440 23714 7450
rect 11200 7416 24218 7426
rect 11080 7392 17066 7402
rect 10720 7368 21266 7378
rect 10576 7344 22298 7354
rect 10552 7320 17474 7330
rect 10288 7296 17306 7306
rect 17632 7296 17642 7306
rect 10024 7272 10658 7282
rect 10672 7272 12482 7282
rect 12760 7272 12794 7282
rect 12856 7272 21314 7282
rect 9952 7248 9986 7258
rect 10072 7248 16514 7258
rect 16528 7248 20858 7258
rect 20872 7248 22058 7258
rect 9928 7224 17618 7234
rect 9880 7200 24194 7210
rect 9856 7176 21386 7186
rect 9832 7152 13130 7162
rect 13672 7152 17858 7162
rect 9472 7128 12962 7138
rect 13048 7128 13154 7138
rect 13480 7128 25490 7138
rect 25504 7128 26858 7138
rect 9112 7104 11138 7114
rect 11152 7104 13226 7114
rect 13240 7104 13706 7114
rect 13720 7104 17978 7114
rect 9064 7080 19490 7090
rect 19504 7080 24986 7090
rect 25000 7080 27290 7090
rect 8992 7056 9086 7066
rect 9448 7056 13802 7066
rect 13816 7056 25682 7066
rect 8296 7032 8306 7042
rect 8440 7032 9458 7042
rect 9472 7032 12722 7042
rect 12736 7032 16730 7042
rect 16744 7032 19322 7042
rect 19336 7032 22250 7042
rect 8224 7008 10298 7018
rect 10504 7008 21146 7018
rect 8200 6984 10922 6994
rect 10936 6984 12722 6994
rect 12736 6984 21098 6994
rect 21112 6984 22562 6994
rect 8176 6960 11714 6970
rect 11728 6960 13226 6970
rect 13240 6960 19106 6970
rect 19120 6960 19946 6970
rect 8152 6936 14714 6946
rect 8128 6912 8258 6922
rect 8272 6912 9410 6922
rect 9424 6912 12050 6922
rect 12064 6912 12266 6922
rect 12280 6912 18146 6922
rect 18160 6912 24650 6922
rect 8104 6888 27458 6898
rect 8008 6864 19778 6874
rect 19792 6864 24986 6874
rect 7888 6840 11690 6850
rect 11704 6840 12338 6850
rect 12352 6840 19706 6850
rect 19720 6840 23666 6850
rect 7816 6816 18170 6826
rect 18184 6816 22826 6826
rect 22840 6816 23186 6826
rect 23200 6816 25202 6826
rect 7792 6792 9026 6802
rect 9040 6792 17738 6802
rect 7768 6768 19082 6778
rect 7720 6744 20546 6754
rect 7624 6720 20378 6730
rect 7600 6696 7610 6706
rect 7672 6696 7874 6706
rect 7888 6696 9122 6706
rect 9136 6696 9746 6706
rect 9760 6696 13538 6706
rect 13552 6696 18146 6706
rect 7504 6672 13274 6682
rect 13336 6672 13826 6682
rect 7384 6648 15074 6658
rect 7360 6624 25922 6634
rect 7336 6600 25442 6610
rect 7312 6576 17402 6586
rect 7288 6552 26018 6562
rect 7192 6528 8930 6538
rect 8944 6528 27074 6538
rect 7048 6504 23738 6514
rect 7000 6480 13130 6490
rect 13144 6480 21434 6490
rect 23800 6480 23834 6490
rect 6856 6456 7538 6466
rect 7552 6456 13334 6466
rect 13348 6456 14426 6466
rect 14440 6456 14618 6466
rect 14632 6456 19826 6466
rect 19840 6456 23282 6466
rect 23296 6456 27002 6466
rect 27016 6456 27218 6466
rect 6784 6432 10394 6442
rect 10456 6432 10682 6442
rect 10960 6432 18674 6442
rect 18688 6432 23786 6442
rect 6664 6408 9554 6418
rect 9568 6408 15962 6418
rect 18040 6408 20330 6418
rect 20800 6408 20954 6418
rect 6616 6384 21938 6394
rect 6544 6360 17426 6370
rect 17440 6360 27866 6370
rect 6472 6336 10946 6346
rect 10960 6336 14690 6346
rect 14704 6336 23858 6346
rect 23872 6336 26498 6346
rect 6400 6312 20786 6322
rect 20800 6312 21122 6322
rect 21136 6312 22706 6322
rect 6328 6288 17090 6298
rect 17944 6288 19226 6298
rect 6136 6264 25178 6274
rect 6112 6240 21842 6250
rect 21856 6240 22442 6250
rect 6040 6216 19394 6226
rect 5872 6192 21602 6202
rect 21616 6192 27434 6202
rect 5824 6168 20666 6178
rect 5776 6144 6626 6154
rect 6640 6144 6746 6154
rect 6760 6144 11522 6154
rect 11536 6144 12530 6154
rect 12544 6144 16010 6154
rect 16024 6144 23498 6154
rect 5728 6120 13922 6130
rect 14848 6120 19178 6130
rect 5680 6096 11354 6106
rect 11368 6096 15122 6106
rect 15136 6096 18122 6106
rect 18136 6096 20642 6106
rect 20656 6096 21626 6106
rect 5488 6072 8978 6082
rect 8992 6072 18218 6082
rect 5464 6048 6986 6058
rect 7000 6048 19730 6058
rect 5440 6024 5570 6034
rect 5584 6024 11930 6034
rect 11944 6024 19922 6034
rect 19936 6024 27314 6034
rect 5392 6000 14810 6010
rect 15880 6000 22610 6010
rect 5344 5976 10826 5986
rect 10840 5976 11162 5986
rect 11176 5976 13442 5986
rect 13456 5976 14570 5986
rect 14584 5976 16586 5986
rect 16600 5976 17810 5986
rect 17824 5976 24674 5986
rect 5320 5952 10850 5962
rect 10864 5952 19898 5962
rect 5248 5928 9698 5938
rect 9712 5928 25514 5938
rect 5152 5904 20642 5914
rect 20656 5904 24194 5914
rect 5104 5880 21626 5890
rect 21640 5880 26786 5890
rect 26800 5880 27338 5890
rect 5080 5856 15938 5866
rect 16048 5856 16106 5866
rect 16192 5856 21866 5866
rect 5032 5832 5210 5842
rect 5224 5832 7514 5842
rect 7528 5832 8666 5842
rect 8680 5832 11426 5842
rect 11440 5832 14042 5842
rect 14056 5832 14330 5842
rect 14344 5832 17786 5842
rect 17800 5832 21914 5842
rect 21928 5832 26402 5842
rect 4936 5808 5714 5818
rect 5728 5808 12074 5818
rect 12088 5808 13106 5818
rect 13120 5808 20234 5818
rect 4888 5784 13970 5794
rect 13984 5784 21434 5794
rect 4864 5760 20306 5770
rect 20704 5760 25754 5770
rect 4696 5736 5354 5746
rect 5368 5736 17450 5746
rect 17464 5736 18482 5746
rect 18496 5736 21722 5746
rect 21736 5736 24002 5746
rect 24016 5736 25898 5746
rect 4672 5712 22658 5722
rect 4648 5688 13034 5698
rect 13048 5688 16490 5698
rect 16504 5688 20690 5698
rect 20704 5688 25826 5698
rect 4576 5664 13634 5674
rect 13648 5664 15986 5674
rect 16000 5664 22130 5674
rect 22144 5664 24554 5674
rect 4504 5640 7898 5650
rect 7912 5640 9338 5650
rect 9352 5640 14450 5650
rect 14464 5640 23474 5650
rect 4432 5616 10874 5626
rect 10984 5616 17450 5626
rect 17920 5616 18194 5626
rect 20488 5616 20714 5626
rect 4384 5592 20138 5602
rect 20464 5592 20618 5602
rect 26920 5592 26930 5602
rect 4312 5568 18914 5578
rect 19000 5568 26906 5578
rect 4264 5544 7250 5554
rect 7264 5544 22154 5554
rect 4216 5520 19274 5530
rect 19528 5520 20810 5530
rect 20824 5520 25010 5530
rect 4192 5496 4466 5506
rect 4480 5496 4538 5506
rect 4552 5496 5282 5506
rect 5296 5496 7970 5506
rect 7984 5496 9938 5506
rect 9952 5496 10346 5506
rect 10360 5496 11258 5506
rect 11272 5496 14834 5506
rect 14848 5496 18038 5506
rect 18052 5496 22178 5506
rect 22192 5496 24698 5506
rect 4048 5472 8786 5482
rect 8800 5472 14258 5482
rect 15688 5472 20762 5482
rect 4000 5448 7418 5458
rect 7432 5448 16346 5458
rect 17728 5448 21050 5458
rect 3976 5424 17042 5434
rect 17056 5424 21158 5434
rect 21172 5424 22034 5434
rect 22048 5424 25850 5434
rect 3880 5400 14546 5410
rect 14920 5400 14978 5410
rect 15208 5400 20066 5410
rect 20368 5400 20498 5410
rect 21256 5400 25130 5410
rect 3856 5376 7682 5386
rect 7696 5376 13418 5386
rect 13432 5376 13754 5386
rect 13768 5376 14066 5386
rect 14080 5376 16178 5386
rect 16192 5376 18098 5386
rect 18112 5376 23378 5386
rect 25240 5376 25250 5386
rect 3832 5352 12506 5362
rect 12520 5352 18890 5362
rect 18904 5352 20282 5362
rect 20296 5352 24506 5362
rect 24520 5352 25226 5362
rect 25240 5352 26642 5362
rect 3784 5328 21458 5338
rect 21760 5328 24410 5338
rect 3760 5304 10154 5314
rect 10168 5304 10202 5314
rect 10216 5304 11378 5314
rect 11392 5304 15050 5314
rect 15064 5304 19994 5314
rect 20272 5304 23810 5314
rect 3736 5280 3938 5290
rect 3952 5280 5858 5290
rect 5872 5280 10010 5290
rect 10024 5280 11546 5290
rect 11560 5280 12290 5290
rect 12304 5280 13082 5290
rect 13096 5280 17138 5290
rect 17152 5280 20882 5290
rect 20896 5280 23474 5290
rect 23488 5280 24530 5290
rect 24544 5280 24722 5290
rect 24736 5280 25874 5290
rect 25888 5280 26738 5290
rect 26752 5280 27194 5290
rect 3712 5256 6674 5266
rect 6736 5256 16082 5266
rect 17704 5256 20978 5266
rect 20992 5256 24938 5266
rect 3688 5232 14666 5242
rect 14872 5232 25586 5242
rect 3640 5208 16298 5218
rect 17200 5208 18578 5218
rect 18976 5208 19010 5218
rect 19384 5208 24530 5218
rect 3568 5184 3914 5194
rect 3928 5184 11978 5194
rect 11992 5184 19562 5194
rect 19576 5184 20426 5194
rect 20440 5184 22658 5194
rect 22672 5184 24950 5194
rect 3544 5160 13730 5170
rect 13744 5160 21410 5170
rect 21424 5160 23306 5170
rect 23416 5160 23546 5170
rect 3496 5136 20522 5146
rect 21232 5136 24338 5146
rect 3472 5112 6434 5122
rect 6448 5112 8282 5122
rect 8296 5112 23354 5122
rect 23368 5112 23402 5122
rect 24496 5112 24626 5122
rect 3448 5088 8642 5098
rect 8656 5088 9194 5098
rect 9208 5088 10106 5098
rect 10120 5088 13514 5098
rect 13528 5088 15002 5098
rect 15016 5088 17018 5098
rect 17032 5088 21554 5098
rect 21568 5088 23906 5098
rect 23920 5088 24482 5098
rect 24496 5088 24890 5098
rect 3400 5064 13670 5074
rect 13684 5064 25706 5074
rect 3136 5040 5618 5050
rect 5632 5040 6458 5050
rect 6472 5040 7226 5050
rect 7240 5040 7850 5050
rect 7864 5040 10418 5050
rect 10432 5040 11810 5050
rect 11824 5040 13490 5050
rect 13504 5040 14930 5050
rect 14944 5040 17258 5050
rect 17272 5040 17378 5050
rect 17392 5040 20186 5050
rect 20200 5040 22034 5050
rect 3064 5016 19034 5026
rect 19264 5016 27242 5026
rect 3040 4992 9962 5002
rect 10048 4992 12086 5002
rect 12100 4992 20954 5002
rect 21040 4992 25082 5002
rect 3016 4968 4082 4978
rect 4168 4968 4250 4978
rect 4264 4968 18962 4978
rect 18976 4968 24290 4978
rect 2968 4944 10898 4954
rect 10912 4944 11906 4954
rect 11920 4944 21986 4954
rect 2944 4920 4514 4930
rect 4528 4920 10178 4930
rect 10192 4920 12314 4930
rect 12448 4920 13874 4930
rect 14656 4920 22970 4930
rect 2920 4896 5906 4906
rect 5920 4896 6818 4906
rect 6832 4896 9290 4906
rect 9304 4896 13058 4906
rect 13072 4896 14234 4906
rect 14248 4896 20450 4906
rect 20464 4896 22682 4906
rect 22696 4896 22922 4906
rect 22936 4896 23258 4906
rect 24064 4896 24410 4906
rect 2848 4872 9050 4882
rect 9064 4872 9170 4882
rect 9400 4872 9482 4882
rect 9640 4872 12218 4882
rect 12232 4872 12650 4882
rect 12664 4872 18386 4882
rect 18400 4872 22490 4882
rect 23152 4872 23330 4882
rect 23608 4872 23642 4882
rect 24040 4872 24062 4882
rect 24616 4872 24734 4882
rect 2800 4848 7010 4858
rect 7024 4848 13898 4858
rect 14104 4848 14306 4858
rect 14320 4848 14342 4858
rect 14608 4848 21758 4858
rect 21832 4848 21950 4858
rect 23128 4848 25034 4858
rect 25120 4848 25154 4858
rect 2752 4824 5786 4834
rect 5992 4824 22106 4834
rect 22120 4824 26690 4834
rect 2728 4800 5690 4810
rect 5704 4800 11570 4810
rect 11584 4800 23930 4810
rect 23944 4800 25106 4810
rect 2704 4776 3170 4786
rect 3184 4776 5642 4786
rect 5656 4776 8810 4786
rect 8824 4776 9506 4786
rect 9520 4776 11354 4786
rect 11368 4776 11642 4786
rect 11656 4776 20570 4786
rect 20584 4776 23882 4786
rect 23896 4776 27602 4786
rect 2656 4752 15314 4762
rect 15760 4752 23618 4762
rect 23680 4752 24146 4762
rect 24304 4752 24362 4762
rect 24688 4752 26378 4762
rect 2608 4728 8474 4738
rect 8584 4728 18938 4738
rect 19096 4728 19106 4738
rect 20056 4728 24434 4738
rect 24904 4728 24950 4738
rect 25480 4728 26234 4738
rect 2536 4704 4130 4714
rect 4144 4704 10130 4714
rect 10144 4704 13610 4714
rect 14128 4704 25730 4714
rect 2512 4680 7034 4690
rect 7048 4680 12122 4690
rect 12136 4680 13298 4690
rect 13312 4680 14210 4690
rect 14224 4680 14522 4690
rect 14536 4680 20474 4690
rect 20488 4680 21338 4690
rect 21352 4680 21386 4690
rect 21400 4680 24026 4690
rect 24040 4680 24122 4690
rect 24136 4680 24458 4690
rect 24472 4680 24602 4690
rect 24616 4680 25634 4690
rect 25648 4680 26762 4690
rect 26776 4680 27794 4690
rect 2488 4656 3650 4666
rect 3664 4656 5882 4666
rect 5896 4656 17162 4666
rect 17176 4656 17234 4666
rect 17248 4656 20906 4666
rect 20920 4656 26954 4666
rect 2440 4632 7562 4642
rect 7576 4632 22010 4642
rect 22360 4632 27122 4642
rect 2392 4608 9362 4618
rect 9376 4608 9530 4618
rect 9544 4608 10274 4618
rect 10288 4608 12002 4618
rect 12016 4608 16058 4618
rect 16072 4608 25418 4618
rect 26776 4608 26786 4618
rect 2368 4584 3098 4594
rect 3112 4584 6242 4594
rect 6256 4584 15026 4594
rect 15040 4584 19058 4594
rect 20416 4584 24098 4594
rect 2320 4560 13850 4570
rect 14176 4560 14738 4570
rect 14752 4560 27818 4570
rect 2272 4536 8234 4546
rect 8248 4536 11618 4546
rect 11632 4536 11954 4546
rect 11968 4536 18722 4546
rect 18856 4536 26930 4546
rect 2248 4512 6098 4522
rect 6112 4512 6170 4522
rect 6184 4512 10538 4522
rect 10552 4512 11330 4522
rect 11344 4512 17834 4522
rect 17848 4512 18074 4522
rect 18088 4512 24866 4522
rect 24880 4512 24914 4522
rect 2200 4488 3482 4498
rect 3496 4488 6698 4498
rect 6712 4488 19634 4498
rect 20896 4488 21050 4498
rect 21352 4488 21602 4498
rect 22480 4488 23834 4498
rect 23848 4488 27362 4498
rect 2176 4464 5834 4474
rect 5848 4464 9386 4474
rect 9400 4464 9818 4474
rect 9832 4464 10226 4474
rect 10240 4464 15866 4474
rect 15880 4464 21674 4474
rect 22528 4464 22850 4474
rect 23224 4464 27722 4474
rect 2056 4440 24818 4450
rect 2032 4416 20594 4426
rect 20608 4416 23162 4426
rect 23320 4416 23426 4426
rect 23944 4416 26090 4426
rect 26104 4416 27890 4426
rect 2008 4392 27554 4402
rect 1936 4368 9578 4378
rect 9592 4368 16034 4378
rect 16048 4368 16994 4378
rect 17008 4368 25346 4378
rect 1912 4344 10562 4354
rect 10576 4344 18794 4354
rect 18808 4344 20546 4354
rect 20920 4344 21158 4354
rect 21568 4344 23546 4354
rect 1888 4320 19442 4330
rect 22864 4320 27770 4330
rect 1840 4296 12458 4306
rect 12520 4296 18458 4306
rect 18472 4296 21794 4306
rect 23368 4296 23498 4306
rect 1816 4272 11450 4282
rect 11464 4272 14378 4282
rect 14560 4272 26258 4282
rect 1768 4248 4754 4258
rect 4768 4248 6242 4258
rect 6304 4248 15530 4258
rect 15952 4248 16010 4258
rect 16144 4248 19658 4258
rect 1768 4224 8450 4234
rect 8704 4224 13994 4234
rect 14224 4224 15914 4234
rect 16408 4224 16826 4234
rect 17416 4224 17474 4234
rect 17536 4224 18266 4234
rect 18352 4224 25778 4234
rect 1696 4200 10082 4210
rect 10144 4200 10154 4210
rect 10480 4200 23954 4210
rect 1672 4176 26354 4186
rect 1648 4152 5642 4162
rect 5656 4152 14450 4162
rect 14464 4152 14498 4162
rect 14512 4152 20018 4162
rect 1624 4128 4898 4138
rect 4912 4128 23234 4138
rect 23248 4128 23570 4138
rect 23584 4128 25394 4138
rect 25408 4128 26810 4138
rect 84 4104 2090 4114
rect 2152 4104 3314 4114
rect 3328 4104 3794 4114
rect 3808 4104 7586 4114
rect 7600 4104 15002 4114
rect 15184 4104 25250 4114
rect 25408 4104 25586 4114
rect 84 4080 10490 4090
rect 10624 4080 12746 4090
rect 12760 4080 15722 4090
rect 15736 4080 26426 4090
rect 84 4056 4538 4066
rect 4600 4056 9242 4066
rect 9256 4056 12386 4066
rect 12688 4056 13154 4066
rect 13312 4056 13670 4066
rect 13864 4056 14234 4066
rect 14392 4056 14618 4066
rect 14680 4056 14690 4066
rect 14872 4056 23522 4066
rect 84 4032 10706 4042
rect 10888 4032 14954 4042
rect 16456 4032 16754 4042
rect 17800 4032 17858 4042
rect 17968 4032 18818 4042
rect 1624 4008 4706 4018
rect 4792 4008 6386 4018
rect 6400 4008 15842 4018
rect 15856 4008 24314 4018
rect 1672 3984 11834 3994
rect 11968 3984 11978 3994
rect 12064 3984 12482 3994
rect 12928 3984 21842 3994
rect 1720 3960 7346 3970
rect 7408 3960 19334 3970
rect 1864 3936 20234 3946
rect 1960 3912 10658 3922
rect 11032 3912 22394 3922
rect 2080 3888 7898 3898
rect 7960 3888 10370 3898
rect 10528 3888 16778 3898
rect 17848 3888 18038 3898
rect 18088 3888 18194 3898
rect 18280 3888 18866 3898
rect 2248 3864 2282 3874
rect 2296 3864 3626 3874
rect 3640 3864 7778 3874
rect 7792 3864 8330 3874
rect 8344 3864 9794 3874
rect 9808 3864 13202 3874
rect 13216 3864 21578 3874
rect 21592 3864 21698 3874
rect 21712 3864 25298 3874
rect 25312 3864 27626 3874
rect 2296 3840 4274 3850
rect 4288 3840 6002 3850
rect 6016 3840 6194 3850
rect 6208 3840 6482 3850
rect 6496 3840 8618 3850
rect 8632 3840 11162 3850
rect 11176 3840 14090 3850
rect 14104 3840 14474 3850
rect 14488 3840 21890 3850
rect 2440 3816 14018 3826
rect 14032 3816 17354 3826
rect 21592 3816 21866 3826
rect 2464 3792 2546 3802
rect 2560 3792 3722 3802
rect 3736 3792 5738 3802
rect 5752 3792 7610 3802
rect 7624 3792 8882 3802
rect 8896 3792 9146 3802
rect 9160 3792 9482 3802
rect 9496 3792 11138 3802
rect 11152 3792 12026 3802
rect 12040 3792 12362 3802
rect 12376 3792 13394 3802
rect 13408 3792 14342 3802
rect 14356 3792 16538 3802
rect 16552 3792 19994 3802
rect 20008 3792 25514 3802
rect 25528 3792 26546 3802
rect 26560 3792 26666 3802
rect 26680 3792 27410 3802
rect 27424 3792 27530 3802
rect 2488 3768 21194 3778
rect 21712 3768 22058 3778
rect 2536 3744 7754 3754
rect 7768 3744 11738 3754
rect 11752 3744 12818 3754
rect 12832 3744 14282 3754
rect 14296 3744 14498 3754
rect 14512 3744 15146 3754
rect 15160 3744 18002 3754
rect 18016 3744 19130 3754
rect 19144 3744 20978 3754
rect 20992 3744 23570 3754
rect 23584 3744 25178 3754
rect 25192 3744 25826 3754
rect 25840 3744 26378 3754
rect 2584 3720 12770 3730
rect 12952 3720 17642 3730
rect 21208 3720 21410 3730
rect 21904 3720 22130 3730
rect 2584 3696 9962 3706
rect 9976 3696 22898 3706
rect 22912 3696 23594 3706
rect 23608 3696 27170 3706
rect 2608 3672 14762 3682
rect 17368 3672 17426 3682
rect 2632 3648 24818 3658
rect 2824 3624 19202 3634
rect 3160 3600 21818 3610
rect 3208 3576 18674 3586
rect 3232 3552 5186 3562
rect 5200 3552 17762 3562
rect 17776 3552 25202 3562
rect 25216 3552 25274 3562
rect 25288 3552 25658 3562
rect 25672 3552 26882 3562
rect 3256 3528 6002 3538
rect 6064 3528 8738 3538
rect 8848 3528 13970 3538
rect 14032 3528 24770 3538
rect 3352 3504 24434 3514
rect 24784 3504 26570 3514
rect 26584 3504 27842 3514
rect 3400 3480 5114 3490
rect 5128 3480 9002 3490
rect 9016 3480 15026 3490
rect 15040 3480 17282 3490
rect 17296 3480 19850 3490
rect 19864 3480 20762 3490
rect 20776 3480 21650 3490
rect 21664 3480 24062 3490
rect 24076 3480 27770 3490
rect 3448 3456 5762 3466
rect 5776 3456 7442 3466
rect 7456 3456 12290 3466
rect 12304 3456 13754 3466
rect 13768 3456 23042 3466
rect 23056 3456 25538 3466
rect 3544 3432 11234 3442
rect 11248 3432 25970 3442
rect 3592 3408 15722 3418
rect 3592 3384 6674 3394
rect 6688 3384 10322 3394
rect 10336 3384 12578 3394
rect 13216 3384 18986 3394
rect 19000 3384 21290 3394
rect 21304 3384 22946 3394
rect 22960 3384 25010 3394
rect 3616 3360 11498 3370
rect 11512 3360 21482 3370
rect 22960 3360 22970 3370
rect 3664 3336 8522 3346
rect 8848 3336 9602 3346
rect 9616 3336 16154 3346
rect 3856 3312 10250 3322
rect 10336 3312 10370 3322
rect 11032 3312 11282 3322
rect 11344 3312 11426 3322
rect 11560 3312 11714 3322
rect 11776 3312 23066 3322
rect 3904 3288 6314 3298
rect 6328 3288 8018 3298
rect 8032 3288 9914 3298
rect 9928 3288 16106 3298
rect 16120 3288 20618 3298
rect 3928 3264 12890 3274
rect 12904 3264 19154 3274
rect 19168 3264 24314 3274
rect 24328 3264 25322 3274
rect 3976 3240 11786 3250
rect 11800 3240 17114 3250
rect 19168 3240 19334 3250
rect 4024 3216 4994 3226
rect 5008 3216 8258 3226
rect 8272 3216 14138 3226
rect 14272 3216 24626 3226
rect 4120 3192 7154 3202
rect 7168 3192 17882 3202
rect 17896 3192 21074 3202
rect 21088 3192 23258 3202
rect 23272 3192 24734 3202
rect 24748 3192 25298 3202
rect 4168 3168 12146 3178
rect 12160 3168 26330 3178
rect 4216 3144 5906 3154
rect 5920 3144 12170 3154
rect 12184 3144 23138 3154
rect 26344 3144 26402 3154
rect 4360 3120 26642 3130
rect 4360 3096 8546 3106
rect 8560 3096 8906 3106
rect 8920 3096 13178 3106
rect 13192 3096 18746 3106
rect 18760 3096 24386 3106
rect 24400 3096 25634 3106
rect 25648 3096 27314 3106
rect 4408 3072 14306 3082
rect 14416 3072 26210 3082
rect 4456 3048 13274 3058
rect 13432 3048 13802 3058
rect 4456 3024 25154 3034
rect 4504 3000 8354 3010
rect 9016 3000 10754 3010
rect 11056 3000 20594 3010
rect 4696 2976 12986 2986
rect 13000 2976 13370 2986
rect 13528 2976 14042 2986
rect 4816 2952 9602 2962
rect 9664 2952 13586 2962
rect 5056 2928 21530 2938
rect 5440 2904 10634 2914
rect 10768 2904 12194 2914
rect 12208 2904 14906 2914
rect 14920 2904 23450 2914
rect 5488 2880 14594 2890
rect 14608 2880 20738 2890
rect 20752 2880 22586 2890
rect 5536 2856 25346 2866
rect 5680 2832 14786 2842
rect 5992 2808 17690 2818
rect 17704 2808 21506 2818
rect 6040 2784 11402 2794
rect 11416 2784 20354 2794
rect 21520 2784 21758 2794
rect 6088 2760 15578 2770
rect 6136 2736 6890 2746
rect 6904 2736 9986 2746
rect 10000 2736 23642 2746
rect 6184 2712 13946 2722
rect 13960 2712 20210 2722
rect 20224 2712 27506 2722
rect 6232 2688 17570 2698
rect 17584 2688 22082 2698
rect 22096 2688 24578 2698
rect 6352 2664 13610 2674
rect 20224 2664 20330 2674
rect 6616 2640 12410 2650
rect 12592 2640 12794 2650
rect 13192 2640 13334 2650
rect 13552 2640 19010 2650
rect 6784 2616 6938 2626
rect 7072 2616 7442 2626
rect 7456 2616 13562 2626
rect 13576 2616 16370 2626
rect 16384 2616 22994 2626
rect 6976 2592 9086 2602
rect 9100 2592 10586 2602
rect 10600 2592 12242 2602
rect 12256 2592 13706 2602
rect 13720 2592 17498 2602
rect 17512 2592 20834 2602
rect 20848 2592 21218 2602
rect 21232 2592 21950 2602
rect 21964 2592 24218 2602
rect 24232 2592 25610 2602
rect 7096 2568 7634 2578
rect 7648 2568 17594 2578
rect 7144 2544 17306 2554
rect 17512 2544 26138 2554
rect 7408 2520 8306 2530
rect 8320 2520 12458 2530
rect 12472 2520 22754 2530
rect 22768 2520 23114 2530
rect 7480 2496 28227 2506
rect 7720 2472 9266 2482
rect 9280 2472 21002 2482
rect 21016 2472 25274 2482
rect 7816 2448 13250 2458
rect 7960 2424 20714 2434
rect 8008 2400 11306 2410
rect 11392 2400 11522 2410
rect 11608 2400 19298 2410
rect 8056 2376 21794 2386
rect 8056 2352 8378 2362
rect 9088 2352 9218 2362
rect 9280 2352 9314 2362
rect 9520 2352 23330 2362
rect 8152 2328 26282 2338
rect 8176 2304 24242 2314
rect 9184 2280 9194 2290
rect 9304 2280 11474 2290
rect 11680 2280 20930 2290
rect 24256 2280 24266 2290
rect 9640 2256 19418 2266
rect 20944 2256 21362 2266
rect 9712 2232 27674 2242
rect 9880 2208 20090 2218
rect 10048 2184 20498 2194
rect 10168 2160 14186 2170
rect 11200 2136 27098 2146
rect 11296 2112 26186 2122
rect 11464 2088 12866 2098
rect 14200 2088 17378 2098
rect 17392 2088 18530 2098
rect 18544 2088 24794 2098
rect 24808 2088 26114 2098
rect 11776 2064 19610 2074
rect 27904 2064 28227 2074
rect 11848 2040 14978 2050
rect 14992 2040 24938 2050
rect 27880 2040 28227 2050
rect 11992 2016 12626 2026
rect 12640 2016 16874 2026
rect 27856 2016 28227 2026
rect 12040 1992 12086 2002
rect 12328 1992 17666 2002
rect 27832 1992 28227 2002
rect 12088 1968 23018 1978
rect 27808 1968 28227 1978
rect 12400 1944 13778 1954
rect 13792 1944 27266 1954
rect 27784 1944 28227 1954
rect 27435 1915 27795 1925
rect 27435 1892 27795 1902
rect 27435 1854 27795 1879
rect 27435 1209 27795 1234
rect 16264 1111 21962 1121
rect 16216 1087 18866 1097
rect 16000 1063 22370 1073
rect 15904 1039 16274 1049
rect 17248 1039 19010 1049
rect 15808 1015 22802 1025
rect 10432 991 11666 1001
rect 11728 991 17858 1001
rect 10384 967 17258 977
rect 17488 967 22298 977
rect 9688 943 25730 953
rect 9352 919 12818 929
rect 12832 919 18050 929
rect 18064 919 21314 929
rect 21328 919 21938 929
rect 21952 919 26570 929
rect 26584 919 26810 929
rect 9136 895 12410 905
rect 12424 895 17570 905
rect 18640 895 24338 905
rect 8440 871 13658 881
rect 13792 871 18602 881
rect 8320 847 20258 857
rect 20320 847 25970 857
rect 8104 823 25802 833
rect 7312 799 9746 809
rect 10072 799 11066 809
rect 11488 799 14354 809
rect 14944 799 21098 809
rect 6880 775 6938 785
rect 7216 775 18650 785
rect 19072 775 22706 785
rect 6832 751 16562 761
rect 16576 751 21170 761
rect 21184 751 24386 761
rect 6760 727 7322 737
rect 7336 727 23618 737
rect 6736 703 13346 713
rect 13456 703 17594 713
rect 17680 703 21242 713
rect 21760 703 23522 713
rect 6520 679 17906 689
rect 18040 679 21914 689
rect 21928 679 24122 689
rect 6352 655 10778 665
rect 10792 655 12842 665
rect 12856 655 22130 665
rect 22144 655 23498 665
rect 23512 655 24002 665
rect 24016 655 26762 665
rect 6280 631 10994 641
rect 11056 631 24722 641
rect 5968 607 22778 617
rect 22792 607 24626 617
rect 5896 583 7658 593
rect 7672 583 8066 593
rect 8080 583 12146 593
rect 12160 583 26834 593
rect 5800 559 22898 569
rect 4960 535 23690 545
rect 4936 511 6554 521
rect 6568 511 19106 521
rect 4816 487 7178 497
rect 7192 487 10826 497
rect 11536 487 20090 497
rect 20104 487 20498 497
rect 4744 463 23162 473
rect 4672 439 11090 449
rect 11872 439 20138 449
rect 4600 415 19346 425
rect 4408 391 25418 401
rect 4336 367 25850 377
rect 4072 343 11426 353
rect 11896 343 13946 353
rect 14080 343 23042 353
rect 4048 319 18482 329
rect 18496 319 21410 329
rect 21424 319 26858 329
rect 3832 295 21890 305
rect 21904 295 26786 305
rect 3760 271 10442 281
rect 10624 271 21770 281
rect 3520 247 21026 257
rect 3376 223 20810 233
rect 20824 223 26714 233
rect 2824 199 18914 209
rect 2704 175 13634 185
rect 15064 175 26618 185
rect 2680 151 17042 161
rect 17296 151 21122 161
rect 1720 127 19898 137
rect 26740 127 28227 137
rect 1648 103 20834 113
rect 26872 103 28227 113
rect 84 79 22274 89
rect 26848 79 28227 89
rect 84 55 1754 65
rect 2656 55 16682 65
rect 16696 55 19754 65
rect 26824 55 28227 65
rect 84 31 12578 41
rect 12640 31 19946 41
rect 26800 31 28227 41
rect 84 7 16442 17
rect 26776 7 28227 17
<< m2contact >>
rect 18818 8775 18832 8789
rect 24734 8775 24748 8789
rect 16922 8751 16936 8765
rect 23198 8751 23212 8765
rect 13370 8727 13384 8741
rect 20126 8727 20140 8741
rect 13034 8703 13048 8717
rect 17054 8703 17068 8717
rect 18674 8703 18688 8717
rect 27842 8703 27856 8717
rect 12242 8679 12256 8693
rect 12674 8679 12688 8693
rect 21662 8679 21676 8693
rect 7130 8655 7144 8669
rect 10850 8655 10864 8669
rect 18866 8655 18880 8669
rect 20102 8655 20116 8669
rect 23834 8655 23848 8669
rect 70 8631 84 8645
rect 25778 8631 25792 8645
rect 70 8607 84 8621
rect 1706 8607 1720 8621
rect 2858 8607 2872 8621
rect 4694 8607 4708 8621
rect 6938 8607 6952 8621
rect 27866 8607 27880 8621
rect 70 8583 84 8597
rect 1754 8583 1768 8597
rect 3110 8583 3124 8597
rect 9218 8583 9232 8597
rect 10346 8583 10360 8597
rect 27818 8583 27832 8597
rect 27842 8583 27856 8597
rect 28227 8583 28241 8597
rect 4658 8559 4672 8573
rect 7826 8559 7840 8573
rect 8738 8559 8752 8573
rect 11090 8559 11104 8573
rect 26270 8559 26284 8573
rect 27722 8559 27736 8573
rect 28227 8559 28241 8573
rect 7082 8535 7096 8549
rect 27842 8535 27856 8549
rect 27866 8535 27880 8549
rect 28227 8535 28241 8549
rect 13946 8511 13960 8525
rect 23186 8511 23200 8525
rect 27770 8511 27784 8525
rect 27794 8511 27808 8525
rect 27842 8511 27856 8525
rect 28227 8511 28241 8525
rect 15494 8487 15508 8501
rect 25562 8487 25576 8501
rect 27794 8487 27808 8501
rect 28227 8487 28241 8501
rect 16826 8463 16840 8477
rect 27794 8463 27808 8477
rect 27818 8463 27832 8477
rect 28227 8463 28241 8477
rect 17030 8439 17044 8453
rect 22850 8439 22864 8453
rect 27794 8439 27808 8453
rect 28227 8439 28241 8453
rect 13106 7606 13120 7620
rect 13778 7606 13792 7620
rect 12194 7582 12208 7596
rect 12962 7582 12976 7596
rect 13082 7582 13096 7596
rect 13250 7582 13264 7596
rect 13826 7582 13840 7596
rect 21362 7582 21376 7596
rect 12098 7558 12112 7572
rect 12650 7558 12664 7572
rect 12770 7558 12784 7572
rect 15890 7558 15904 7572
rect 11786 7534 11800 7548
rect 24266 7534 24280 7548
rect 11714 7510 11728 7524
rect 24362 7510 24376 7524
rect 11642 7486 11656 7500
rect 23426 7486 23440 7500
rect 25562 7486 25576 7500
rect 25778 7486 25792 7500
rect 11258 7462 11272 7476
rect 11306 7462 11320 7476
rect 11570 7462 11584 7476
rect 11786 7462 11800 7476
rect 11882 7462 11896 7476
rect 25562 7462 25576 7476
rect 11234 7438 11248 7452
rect 23714 7438 23728 7452
rect 11186 7414 11200 7428
rect 24218 7414 24232 7428
rect 11066 7390 11080 7404
rect 17066 7390 17080 7404
rect 10706 7366 10720 7380
rect 21266 7366 21280 7380
rect 10562 7342 10576 7356
rect 22298 7342 22312 7356
rect 10538 7318 10552 7332
rect 17474 7318 17488 7332
rect 10274 7294 10288 7308
rect 17306 7294 17320 7308
rect 17618 7294 17632 7308
rect 17642 7294 17656 7308
rect 10010 7270 10024 7284
rect 10658 7270 10672 7284
rect 12482 7270 12496 7284
rect 12746 7270 12760 7284
rect 12794 7270 12808 7284
rect 12842 7270 12856 7284
rect 21314 7270 21328 7284
rect 9938 7246 9952 7260
rect 9986 7246 10000 7260
rect 10058 7246 10072 7260
rect 16514 7246 16528 7260
rect 20858 7246 20872 7260
rect 22058 7246 22072 7260
rect 9914 7222 9928 7236
rect 17618 7222 17632 7236
rect 9866 7198 9880 7212
rect 24194 7198 24208 7212
rect 9842 7174 9856 7188
rect 21386 7174 21400 7188
rect 9818 7150 9832 7164
rect 13130 7150 13144 7164
rect 13658 7150 13672 7164
rect 17858 7150 17872 7164
rect 9458 7126 9472 7140
rect 12962 7126 12976 7140
rect 13034 7126 13048 7140
rect 13154 7126 13168 7140
rect 13466 7126 13480 7140
rect 25490 7126 25504 7140
rect 26858 7126 26872 7140
rect 9098 7102 9112 7116
rect 11138 7102 11152 7116
rect 13226 7102 13240 7116
rect 13706 7102 13720 7116
rect 17978 7102 17992 7116
rect 9050 7078 9064 7092
rect 19490 7078 19504 7092
rect 24986 7078 25000 7092
rect 27290 7078 27304 7092
rect 8978 7054 8992 7068
rect 9086 7054 9100 7068
rect 9434 7054 9448 7068
rect 13802 7054 13816 7068
rect 25682 7054 25696 7068
rect 8282 7030 8296 7044
rect 8306 7030 8320 7044
rect 8426 7030 8440 7044
rect 9458 7030 9472 7044
rect 12722 7030 12736 7044
rect 16730 7030 16744 7044
rect 19322 7030 19336 7044
rect 22250 7030 22264 7044
rect 8210 7006 8224 7020
rect 10298 7006 10312 7020
rect 10490 7006 10504 7020
rect 21146 7006 21160 7020
rect 8186 6982 8200 6996
rect 10922 6982 10936 6996
rect 12722 6982 12736 6996
rect 21098 6982 21112 6996
rect 22562 6982 22576 6996
rect 8162 6958 8176 6972
rect 11714 6958 11728 6972
rect 13226 6958 13240 6972
rect 19106 6958 19120 6972
rect 19946 6958 19960 6972
rect 8138 6934 8152 6948
rect 14714 6934 14728 6948
rect 8114 6910 8128 6924
rect 8258 6910 8272 6924
rect 9410 6910 9424 6924
rect 12050 6910 12064 6924
rect 12266 6910 12280 6924
rect 18146 6910 18160 6924
rect 24650 6910 24664 6924
rect 8090 6886 8104 6900
rect 27458 6886 27472 6900
rect 7994 6862 8008 6876
rect 19778 6862 19792 6876
rect 24986 6862 25000 6876
rect 7874 6838 7888 6852
rect 11690 6838 11704 6852
rect 12338 6838 12352 6852
rect 19706 6838 19720 6852
rect 23666 6838 23680 6852
rect 7802 6814 7816 6828
rect 18170 6814 18184 6828
rect 22826 6814 22840 6828
rect 23186 6814 23200 6828
rect 25202 6814 25216 6828
rect 7778 6790 7792 6804
rect 9026 6790 9040 6804
rect 17738 6790 17752 6804
rect 7754 6766 7768 6780
rect 19082 6766 19096 6780
rect 7706 6742 7720 6756
rect 20546 6742 20560 6756
rect 7610 6718 7624 6732
rect 20378 6718 20392 6732
rect 7586 6694 7600 6708
rect 7610 6694 7624 6708
rect 7658 6694 7672 6708
rect 7874 6694 7888 6708
rect 9122 6694 9136 6708
rect 9746 6694 9760 6708
rect 13538 6694 13552 6708
rect 18146 6694 18160 6708
rect 7490 6670 7504 6684
rect 13274 6670 13288 6684
rect 13322 6670 13336 6684
rect 13826 6670 13840 6684
rect 7370 6646 7384 6660
rect 15074 6646 15088 6660
rect 7346 6622 7360 6636
rect 25922 6622 25936 6636
rect 7322 6598 7336 6612
rect 25442 6598 25456 6612
rect 7298 6574 7312 6588
rect 17402 6574 17416 6588
rect 7274 6550 7288 6564
rect 26018 6550 26032 6564
rect 7178 6526 7192 6540
rect 8930 6526 8944 6540
rect 27074 6526 27088 6540
rect 7034 6502 7048 6516
rect 23738 6502 23752 6516
rect 6986 6478 7000 6492
rect 13130 6478 13144 6492
rect 21434 6478 21448 6492
rect 23786 6478 23800 6492
rect 23834 6478 23848 6492
rect 6842 6454 6856 6468
rect 7538 6454 7552 6468
rect 13334 6454 13348 6468
rect 14426 6454 14440 6468
rect 14618 6454 14632 6468
rect 19826 6454 19840 6468
rect 23282 6454 23296 6468
rect 27002 6454 27016 6468
rect 27218 6454 27232 6468
rect 6770 6430 6784 6444
rect 10394 6430 10408 6444
rect 10442 6430 10456 6444
rect 10682 6430 10696 6444
rect 10946 6430 10960 6444
rect 18674 6430 18688 6444
rect 23786 6430 23800 6444
rect 6650 6406 6664 6420
rect 9554 6406 9568 6420
rect 15962 6406 15976 6420
rect 18026 6406 18040 6420
rect 20330 6406 20344 6420
rect 20786 6406 20800 6420
rect 20954 6406 20968 6420
rect 6602 6382 6616 6396
rect 21938 6382 21952 6396
rect 6530 6358 6544 6372
rect 17426 6358 17440 6372
rect 27866 6358 27880 6372
rect 6458 6334 6472 6348
rect 10946 6334 10960 6348
rect 14690 6334 14704 6348
rect 23858 6334 23872 6348
rect 26498 6334 26512 6348
rect 6386 6310 6400 6324
rect 20786 6310 20800 6324
rect 21122 6310 21136 6324
rect 22706 6310 22720 6324
rect 6314 6286 6328 6300
rect 17090 6286 17104 6300
rect 17930 6286 17944 6300
rect 19226 6286 19240 6300
rect 6122 6262 6136 6276
rect 25178 6262 25192 6276
rect 6098 6238 6112 6252
rect 21842 6238 21856 6252
rect 22442 6238 22456 6252
rect 6026 6214 6040 6228
rect 19394 6214 19408 6228
rect 5858 6190 5872 6204
rect 21602 6190 21616 6204
rect 27434 6190 27448 6204
rect 5810 6166 5824 6180
rect 20666 6166 20680 6180
rect 5762 6142 5776 6156
rect 6626 6142 6640 6156
rect 6746 6142 6760 6156
rect 11522 6142 11536 6156
rect 12530 6142 12544 6156
rect 16010 6142 16024 6156
rect 23498 6142 23512 6156
rect 5714 6118 5728 6132
rect 13922 6118 13936 6132
rect 14834 6118 14848 6132
rect 19178 6118 19192 6132
rect 5666 6094 5680 6108
rect 11354 6094 11368 6108
rect 15122 6094 15136 6108
rect 18122 6094 18136 6108
rect 20642 6094 20656 6108
rect 21626 6094 21640 6108
rect 5474 6070 5488 6084
rect 8978 6070 8992 6084
rect 18218 6070 18232 6084
rect 5450 6046 5464 6060
rect 6986 6046 7000 6060
rect 19730 6046 19744 6060
rect 5426 6022 5440 6036
rect 5570 6022 5584 6036
rect 11930 6022 11944 6036
rect 19922 6022 19936 6036
rect 27314 6022 27328 6036
rect 5378 5998 5392 6012
rect 14810 5998 14824 6012
rect 15866 5998 15880 6012
rect 22610 5998 22624 6012
rect 5330 5974 5344 5988
rect 10826 5974 10840 5988
rect 11162 5974 11176 5988
rect 13442 5974 13456 5988
rect 14570 5974 14584 5988
rect 16586 5974 16600 5988
rect 17810 5974 17824 5988
rect 24674 5974 24688 5988
rect 5306 5950 5320 5964
rect 10850 5950 10864 5964
rect 19898 5950 19912 5964
rect 5234 5926 5248 5940
rect 9698 5926 9712 5940
rect 25514 5926 25528 5940
rect 5138 5902 5152 5916
rect 20642 5902 20656 5916
rect 24194 5902 24208 5916
rect 5090 5878 5104 5892
rect 21626 5878 21640 5892
rect 26786 5878 26800 5892
rect 27338 5878 27352 5892
rect 5066 5854 5080 5868
rect 15938 5854 15952 5868
rect 16034 5854 16048 5868
rect 16106 5854 16120 5868
rect 16178 5854 16192 5868
rect 21866 5854 21880 5868
rect 5018 5830 5032 5844
rect 5210 5830 5224 5844
rect 7514 5830 7528 5844
rect 8666 5830 8680 5844
rect 11426 5830 11440 5844
rect 14042 5830 14056 5844
rect 14330 5830 14344 5844
rect 17786 5830 17800 5844
rect 21914 5830 21928 5844
rect 26402 5830 26416 5844
rect 4922 5806 4936 5820
rect 5714 5806 5728 5820
rect 12074 5806 12088 5820
rect 13106 5806 13120 5820
rect 20234 5806 20248 5820
rect 4874 5782 4888 5796
rect 13970 5782 13984 5796
rect 21434 5782 21448 5796
rect 4850 5758 4864 5772
rect 20306 5758 20320 5772
rect 20690 5758 20704 5772
rect 25754 5758 25768 5772
rect 4682 5734 4696 5748
rect 5354 5734 5368 5748
rect 17450 5734 17464 5748
rect 18482 5734 18496 5748
rect 21722 5734 21736 5748
rect 24002 5734 24016 5748
rect 25898 5734 25912 5748
rect 4658 5710 4672 5724
rect 22658 5710 22672 5724
rect 4634 5686 4648 5700
rect 13034 5686 13048 5700
rect 16490 5686 16504 5700
rect 20690 5686 20704 5700
rect 25826 5686 25840 5700
rect 4562 5662 4576 5676
rect 13634 5662 13648 5676
rect 15986 5662 16000 5676
rect 22130 5662 22144 5676
rect 24554 5662 24568 5676
rect 4490 5638 4504 5652
rect 7898 5638 7912 5652
rect 9338 5638 9352 5652
rect 14450 5638 14464 5652
rect 23474 5638 23488 5652
rect 4418 5614 4432 5628
rect 10874 5614 10888 5628
rect 10970 5614 10984 5628
rect 17450 5614 17464 5628
rect 17906 5614 17920 5628
rect 18194 5614 18208 5628
rect 20474 5614 20488 5628
rect 20714 5614 20728 5628
rect 4370 5590 4384 5604
rect 20138 5590 20152 5604
rect 20450 5590 20464 5604
rect 20618 5590 20632 5604
rect 26906 5590 26920 5604
rect 26930 5590 26944 5604
rect 4298 5566 4312 5580
rect 18914 5566 18928 5580
rect 18986 5566 19000 5580
rect 26906 5566 26920 5580
rect 4250 5542 4264 5556
rect 7250 5542 7264 5556
rect 22154 5542 22168 5556
rect 4202 5518 4216 5532
rect 19274 5518 19288 5532
rect 19514 5518 19528 5532
rect 20810 5518 20824 5532
rect 25010 5518 25024 5532
rect 4178 5494 4192 5508
rect 4466 5494 4480 5508
rect 4538 5494 4552 5508
rect 5282 5494 5296 5508
rect 7970 5494 7984 5508
rect 9938 5494 9952 5508
rect 10346 5494 10360 5508
rect 11258 5494 11272 5508
rect 14834 5494 14848 5508
rect 18038 5494 18052 5508
rect 22178 5494 22192 5508
rect 24698 5494 24712 5508
rect 4034 5470 4048 5484
rect 8786 5470 8800 5484
rect 14258 5470 14272 5484
rect 15674 5470 15688 5484
rect 20762 5470 20776 5484
rect 3986 5446 4000 5460
rect 7418 5446 7432 5460
rect 16346 5446 16360 5460
rect 17714 5446 17728 5460
rect 21050 5446 21064 5460
rect 3962 5422 3976 5436
rect 17042 5422 17056 5436
rect 21158 5422 21172 5436
rect 22034 5422 22048 5436
rect 25850 5422 25864 5436
rect 3866 5398 3880 5412
rect 14546 5398 14560 5412
rect 14906 5398 14920 5412
rect 14978 5398 14992 5412
rect 15194 5398 15208 5412
rect 20066 5398 20080 5412
rect 20354 5398 20368 5412
rect 20498 5398 20512 5412
rect 21242 5398 21256 5412
rect 25130 5398 25144 5412
rect 3842 5374 3856 5388
rect 7682 5374 7696 5388
rect 13418 5374 13432 5388
rect 13754 5374 13768 5388
rect 14066 5374 14080 5388
rect 16178 5374 16192 5388
rect 18098 5374 18112 5388
rect 23378 5374 23392 5388
rect 25226 5374 25240 5388
rect 25250 5374 25264 5388
rect 3818 5350 3832 5364
rect 12506 5350 12520 5364
rect 18890 5350 18904 5364
rect 20282 5350 20296 5364
rect 24506 5350 24520 5364
rect 25226 5350 25240 5364
rect 26642 5350 26656 5364
rect 3770 5326 3784 5340
rect 21458 5326 21472 5340
rect 21746 5326 21760 5340
rect 24410 5326 24424 5340
rect 3746 5302 3760 5316
rect 10154 5302 10168 5316
rect 10202 5302 10216 5316
rect 11378 5302 11392 5316
rect 15050 5302 15064 5316
rect 19994 5302 20008 5316
rect 20258 5302 20272 5316
rect 23810 5302 23824 5316
rect 3722 5278 3736 5292
rect 3938 5278 3952 5292
rect 5858 5278 5872 5292
rect 10010 5278 10024 5292
rect 11546 5278 11560 5292
rect 12290 5278 12304 5292
rect 13082 5278 13096 5292
rect 17138 5278 17152 5292
rect 20882 5278 20896 5292
rect 23474 5278 23488 5292
rect 24530 5278 24544 5292
rect 24722 5278 24736 5292
rect 25874 5278 25888 5292
rect 26738 5278 26752 5292
rect 27194 5278 27208 5292
rect 3698 5254 3712 5268
rect 6674 5254 6688 5268
rect 6722 5254 6736 5268
rect 16082 5254 16096 5268
rect 17690 5254 17704 5268
rect 20978 5254 20992 5268
rect 24938 5254 24952 5268
rect 3674 5230 3688 5244
rect 14666 5230 14680 5244
rect 14858 5230 14872 5244
rect 25586 5230 25600 5244
rect 3626 5206 3640 5220
rect 16298 5206 16312 5220
rect 17186 5206 17200 5220
rect 18578 5206 18592 5220
rect 18962 5206 18976 5220
rect 19010 5206 19024 5220
rect 19370 5206 19384 5220
rect 24530 5206 24544 5220
rect 3554 5182 3568 5196
rect 3914 5182 3928 5196
rect 11978 5182 11992 5196
rect 19562 5182 19576 5196
rect 20426 5182 20440 5196
rect 22658 5182 22672 5196
rect 24950 5182 24964 5196
rect 3530 5158 3544 5172
rect 13730 5158 13744 5172
rect 21410 5158 21424 5172
rect 23306 5158 23320 5172
rect 23402 5158 23416 5172
rect 23546 5158 23560 5172
rect 3482 5134 3496 5148
rect 20522 5134 20536 5148
rect 21218 5134 21232 5148
rect 24338 5134 24352 5148
rect 3458 5110 3472 5124
rect 6434 5110 6448 5124
rect 8282 5110 8296 5124
rect 23354 5110 23368 5124
rect 23402 5110 23416 5124
rect 24482 5110 24496 5124
rect 24626 5110 24640 5124
rect 3434 5086 3448 5100
rect 8642 5086 8656 5100
rect 9194 5086 9208 5100
rect 10106 5086 10120 5100
rect 13514 5086 13528 5100
rect 15002 5086 15016 5100
rect 17018 5086 17032 5100
rect 21554 5086 21568 5100
rect 23906 5086 23920 5100
rect 24482 5086 24496 5100
rect 24890 5086 24904 5100
rect 3386 5062 3400 5076
rect 13670 5062 13684 5076
rect 25706 5062 25720 5076
rect 3122 5038 3136 5052
rect 5618 5038 5632 5052
rect 6458 5038 6472 5052
rect 7226 5038 7240 5052
rect 7850 5038 7864 5052
rect 10418 5038 10432 5052
rect 11810 5038 11824 5052
rect 13490 5038 13504 5052
rect 14930 5038 14944 5052
rect 17258 5038 17272 5052
rect 17378 5038 17392 5052
rect 20186 5038 20200 5052
rect 22034 5038 22048 5052
rect 3050 5014 3064 5028
rect 19034 5014 19048 5028
rect 19250 5014 19264 5028
rect 27242 5014 27256 5028
rect 3026 4990 3040 5004
rect 9962 4990 9976 5004
rect 10034 4990 10048 5004
rect 12086 4990 12100 5004
rect 20954 4990 20968 5004
rect 21026 4990 21040 5004
rect 25082 4990 25096 5004
rect 3002 4966 3016 4980
rect 4082 4966 4096 4980
rect 4154 4966 4168 4980
rect 4250 4966 4264 4980
rect 18962 4966 18976 4980
rect 24290 4966 24304 4980
rect 2954 4942 2968 4956
rect 10898 4942 10912 4956
rect 11906 4942 11920 4956
rect 21986 4942 22000 4956
rect 2930 4918 2944 4932
rect 4514 4918 4528 4932
rect 10178 4918 10192 4932
rect 12314 4918 12328 4932
rect 12434 4918 12448 4932
rect 13874 4918 13888 4932
rect 14642 4918 14656 4932
rect 22970 4918 22984 4932
rect 2906 4894 2920 4908
rect 5906 4894 5920 4908
rect 6818 4894 6832 4908
rect 9290 4894 9304 4908
rect 13058 4894 13072 4908
rect 14234 4894 14248 4908
rect 20450 4894 20464 4908
rect 22682 4894 22696 4908
rect 22922 4894 22936 4908
rect 23258 4894 23272 4908
rect 24050 4894 24064 4908
rect 24410 4894 24424 4908
rect 2834 4870 2848 4884
rect 9050 4870 9064 4884
rect 9170 4870 9184 4884
rect 9386 4870 9400 4884
rect 9482 4870 9496 4884
rect 9626 4870 9640 4884
rect 12218 4870 12232 4884
rect 12650 4870 12664 4884
rect 18386 4870 18400 4884
rect 22490 4870 22504 4884
rect 23138 4870 23152 4884
rect 23330 4870 23344 4884
rect 23594 4870 23608 4884
rect 23642 4870 23656 4884
rect 24026 4870 24040 4884
rect 24062 4870 24076 4884
rect 24602 4870 24616 4884
rect 24734 4870 24748 4884
rect 2786 4846 2800 4860
rect 7010 4846 7024 4860
rect 13898 4846 13912 4860
rect 14090 4846 14104 4860
rect 14306 4846 14320 4860
rect 14342 4846 14356 4860
rect 14594 4846 14608 4860
rect 21758 4846 21772 4860
rect 21818 4846 21832 4860
rect 21950 4846 21964 4860
rect 23114 4846 23128 4860
rect 25034 4846 25048 4860
rect 25106 4846 25120 4860
rect 25154 4846 25168 4860
rect 2738 4822 2752 4836
rect 5786 4822 5800 4836
rect 5978 4822 5992 4836
rect 22106 4822 22120 4836
rect 26690 4822 26704 4836
rect 2714 4798 2728 4812
rect 5690 4798 5704 4812
rect 11570 4798 11584 4812
rect 23930 4798 23944 4812
rect 25106 4798 25120 4812
rect 2690 4774 2704 4788
rect 3170 4774 3184 4788
rect 5642 4774 5656 4788
rect 8810 4774 8824 4788
rect 9506 4774 9520 4788
rect 11354 4774 11368 4788
rect 11642 4774 11656 4788
rect 20570 4774 20584 4788
rect 23882 4774 23896 4788
rect 27602 4774 27616 4788
rect 2642 4750 2656 4764
rect 15314 4750 15328 4764
rect 15746 4750 15760 4764
rect 23618 4750 23632 4764
rect 23666 4750 23680 4764
rect 24146 4750 24160 4764
rect 24290 4750 24304 4764
rect 24362 4750 24376 4764
rect 24674 4750 24688 4764
rect 26378 4750 26392 4764
rect 2594 4726 2608 4740
rect 8474 4726 8488 4740
rect 8570 4726 8584 4740
rect 18938 4726 18952 4740
rect 19082 4726 19096 4740
rect 19106 4726 19120 4740
rect 20042 4726 20056 4740
rect 24434 4726 24448 4740
rect 24890 4726 24904 4740
rect 24950 4726 24964 4740
rect 25466 4726 25480 4740
rect 26234 4726 26248 4740
rect 2522 4702 2536 4716
rect 4130 4702 4144 4716
rect 10130 4702 10144 4716
rect 13610 4702 13624 4716
rect 14114 4702 14128 4716
rect 25730 4702 25744 4716
rect 2498 4678 2512 4692
rect 7034 4678 7048 4692
rect 12122 4678 12136 4692
rect 13298 4678 13312 4692
rect 14210 4678 14224 4692
rect 14522 4678 14536 4692
rect 20474 4678 20488 4692
rect 21338 4678 21352 4692
rect 21386 4678 21400 4692
rect 24026 4678 24040 4692
rect 24122 4678 24136 4692
rect 24458 4678 24472 4692
rect 24602 4678 24616 4692
rect 25634 4678 25648 4692
rect 26762 4678 26776 4692
rect 27794 4678 27808 4692
rect 2474 4654 2488 4668
rect 3650 4654 3664 4668
rect 5882 4654 5896 4668
rect 17162 4654 17176 4668
rect 17234 4654 17248 4668
rect 20906 4654 20920 4668
rect 26954 4654 26968 4668
rect 2426 4630 2440 4644
rect 7562 4630 7576 4644
rect 22010 4630 22024 4644
rect 22346 4630 22360 4644
rect 27122 4630 27136 4644
rect 2378 4606 2392 4620
rect 9362 4606 9376 4620
rect 9530 4606 9544 4620
rect 10274 4606 10288 4620
rect 12002 4606 12016 4620
rect 16058 4606 16072 4620
rect 25418 4606 25432 4620
rect 26762 4606 26776 4620
rect 26786 4606 26800 4620
rect 2354 4582 2368 4596
rect 3098 4582 3112 4596
rect 6242 4582 6256 4596
rect 15026 4582 15040 4596
rect 19058 4582 19072 4596
rect 20402 4582 20416 4596
rect 24098 4582 24112 4596
rect 2306 4558 2320 4572
rect 13850 4558 13864 4572
rect 14162 4558 14176 4572
rect 14738 4558 14752 4572
rect 27818 4558 27832 4572
rect 2258 4534 2272 4548
rect 8234 4534 8248 4548
rect 11618 4534 11632 4548
rect 11954 4534 11968 4548
rect 18722 4534 18736 4548
rect 18842 4534 18856 4548
rect 26930 4534 26944 4548
rect 2234 4510 2248 4524
rect 6098 4510 6112 4524
rect 6170 4510 6184 4524
rect 10538 4510 10552 4524
rect 11330 4510 11344 4524
rect 17834 4510 17848 4524
rect 18074 4510 18088 4524
rect 24866 4510 24880 4524
rect 24914 4510 24928 4524
rect 2186 4486 2200 4500
rect 3482 4486 3496 4500
rect 6698 4486 6712 4500
rect 19634 4486 19648 4500
rect 20882 4486 20896 4500
rect 21050 4486 21064 4500
rect 21338 4486 21352 4500
rect 21602 4486 21616 4500
rect 22466 4486 22480 4500
rect 23834 4486 23848 4500
rect 27362 4486 27376 4500
rect 2162 4462 2176 4476
rect 5834 4462 5848 4476
rect 9386 4462 9400 4476
rect 9818 4462 9832 4476
rect 10226 4462 10240 4476
rect 15866 4462 15880 4476
rect 21674 4462 21688 4476
rect 22514 4462 22528 4476
rect 22850 4462 22864 4476
rect 23210 4462 23224 4476
rect 27722 4462 27736 4476
rect 2042 4438 2056 4452
rect 24818 4438 24832 4452
rect 2018 4414 2032 4428
rect 20594 4414 20608 4428
rect 23162 4414 23176 4428
rect 23306 4414 23320 4428
rect 23426 4414 23440 4428
rect 23930 4414 23944 4428
rect 26090 4414 26104 4428
rect 27890 4414 27904 4428
rect 1994 4390 2008 4404
rect 27554 4390 27568 4404
rect 1922 4366 1936 4380
rect 9578 4366 9592 4380
rect 16034 4366 16048 4380
rect 16994 4366 17008 4380
rect 25346 4366 25360 4380
rect 1898 4342 1912 4356
rect 10562 4342 10576 4356
rect 18794 4342 18808 4356
rect 20546 4342 20560 4356
rect 20906 4342 20920 4356
rect 21158 4342 21172 4356
rect 21554 4342 21568 4356
rect 23546 4342 23560 4356
rect 1874 4318 1888 4332
rect 19442 4318 19456 4332
rect 22850 4318 22864 4332
rect 27770 4318 27784 4332
rect 1826 4294 1840 4308
rect 12458 4294 12472 4308
rect 12506 4294 12520 4308
rect 18458 4294 18472 4308
rect 21794 4294 21808 4308
rect 23354 4294 23368 4308
rect 23498 4294 23512 4308
rect 1802 4270 1816 4284
rect 11450 4270 11464 4284
rect 14378 4270 14392 4284
rect 14546 4270 14560 4284
rect 26258 4270 26272 4284
rect 1754 4246 1768 4260
rect 4754 4246 4768 4260
rect 6242 4246 6256 4260
rect 6290 4246 6304 4260
rect 15530 4246 15544 4260
rect 15938 4246 15952 4260
rect 16010 4246 16024 4260
rect 16130 4246 16144 4260
rect 19658 4246 19672 4260
rect 1754 4222 1768 4236
rect 8450 4222 8464 4236
rect 8690 4222 8704 4236
rect 13994 4222 14008 4236
rect 14210 4222 14224 4236
rect 15914 4222 15928 4236
rect 16394 4222 16408 4236
rect 16826 4222 16840 4236
rect 17402 4222 17416 4236
rect 17474 4222 17488 4236
rect 17522 4222 17536 4236
rect 18266 4222 18280 4236
rect 18338 4222 18352 4236
rect 25778 4222 25792 4236
rect 1682 4198 1696 4212
rect 10082 4198 10096 4212
rect 10130 4198 10144 4212
rect 10154 4198 10168 4212
rect 10466 4198 10480 4212
rect 23954 4198 23968 4212
rect 1658 4174 1672 4188
rect 26354 4174 26368 4188
rect 1634 4150 1648 4164
rect 5642 4150 5656 4164
rect 14450 4150 14464 4164
rect 14498 4150 14512 4164
rect 20018 4150 20032 4164
rect 1610 4126 1624 4140
rect 4898 4126 4912 4140
rect 23234 4126 23248 4140
rect 23570 4126 23584 4140
rect 25394 4126 25408 4140
rect 26810 4126 26824 4140
rect 70 4102 84 4116
rect 2090 4102 2104 4116
rect 2138 4102 2152 4116
rect 3314 4102 3328 4116
rect 3794 4102 3808 4116
rect 7586 4102 7600 4116
rect 15002 4102 15016 4116
rect 15170 4102 15184 4116
rect 25250 4102 25264 4116
rect 25394 4102 25408 4116
rect 25586 4102 25600 4116
rect 70 4078 84 4092
rect 10490 4078 10504 4092
rect 10610 4078 10624 4092
rect 12746 4078 12760 4092
rect 15722 4078 15736 4092
rect 26426 4078 26440 4092
rect 70 4054 84 4068
rect 4538 4054 4552 4068
rect 4586 4054 4600 4068
rect 9242 4054 9256 4068
rect 12386 4054 12400 4068
rect 12674 4054 12688 4068
rect 13154 4054 13168 4068
rect 13298 4054 13312 4068
rect 13670 4054 13684 4068
rect 13850 4054 13864 4068
rect 14234 4054 14248 4068
rect 14378 4054 14392 4068
rect 14618 4054 14632 4068
rect 14666 4054 14680 4068
rect 14690 4054 14704 4068
rect 14858 4054 14872 4068
rect 23522 4054 23536 4068
rect 70 4030 84 4044
rect 10706 4030 10720 4044
rect 10874 4030 10888 4044
rect 14954 4030 14968 4044
rect 16442 4030 16456 4044
rect 16754 4030 16768 4044
rect 17786 4030 17800 4044
rect 17858 4030 17872 4044
rect 17954 4030 17968 4044
rect 18818 4030 18832 4044
rect 1610 4006 1624 4020
rect 4706 4006 4720 4020
rect 4778 4006 4792 4020
rect 6386 4006 6400 4020
rect 15842 4006 15856 4020
rect 24314 4006 24328 4020
rect 1658 3982 1672 3996
rect 11834 3982 11848 3996
rect 11954 3982 11968 3996
rect 11978 3982 11992 3996
rect 12050 3982 12064 3996
rect 12482 3982 12496 3996
rect 12914 3982 12928 3996
rect 21842 3982 21856 3996
rect 1706 3958 1720 3972
rect 7346 3958 7360 3972
rect 7394 3958 7408 3972
rect 19334 3958 19348 3972
rect 1850 3934 1864 3948
rect 20234 3934 20248 3948
rect 1946 3910 1960 3924
rect 10658 3910 10672 3924
rect 11018 3910 11032 3924
rect 22394 3910 22408 3924
rect 2066 3886 2080 3900
rect 7898 3886 7912 3900
rect 7946 3886 7960 3900
rect 10370 3886 10384 3900
rect 10514 3886 10528 3900
rect 16778 3886 16792 3900
rect 17834 3886 17848 3900
rect 18038 3886 18052 3900
rect 18074 3886 18088 3900
rect 18194 3886 18208 3900
rect 18266 3886 18280 3900
rect 18866 3886 18880 3900
rect 2234 3862 2248 3876
rect 2282 3862 2296 3876
rect 3626 3862 3640 3876
rect 7778 3862 7792 3876
rect 8330 3862 8344 3876
rect 9794 3862 9808 3876
rect 13202 3862 13216 3876
rect 21578 3862 21592 3876
rect 21698 3862 21712 3876
rect 25298 3862 25312 3876
rect 27626 3862 27640 3876
rect 2282 3838 2296 3852
rect 4274 3838 4288 3852
rect 6002 3838 6016 3852
rect 6194 3838 6208 3852
rect 6482 3838 6496 3852
rect 8618 3838 8632 3852
rect 11162 3838 11176 3852
rect 14090 3838 14104 3852
rect 14474 3838 14488 3852
rect 21890 3838 21904 3852
rect 2426 3814 2440 3828
rect 14018 3814 14032 3828
rect 17354 3814 17368 3828
rect 21578 3814 21592 3828
rect 21866 3814 21880 3828
rect 2450 3790 2464 3804
rect 2546 3790 2560 3804
rect 3722 3790 3736 3804
rect 5738 3790 5752 3804
rect 7610 3790 7624 3804
rect 8882 3790 8896 3804
rect 9146 3790 9160 3804
rect 9482 3790 9496 3804
rect 11138 3790 11152 3804
rect 12026 3790 12040 3804
rect 12362 3790 12376 3804
rect 13394 3790 13408 3804
rect 14342 3790 14356 3804
rect 16538 3790 16552 3804
rect 19994 3790 20008 3804
rect 25514 3790 25528 3804
rect 26546 3790 26560 3804
rect 26666 3790 26680 3804
rect 27410 3790 27424 3804
rect 27530 3790 27544 3804
rect 2474 3766 2488 3780
rect 21194 3766 21208 3780
rect 21698 3766 21712 3780
rect 22058 3766 22072 3780
rect 2522 3742 2536 3756
rect 7754 3742 7768 3756
rect 11738 3742 11752 3756
rect 12818 3742 12832 3756
rect 14282 3742 14296 3756
rect 14498 3742 14512 3756
rect 15146 3742 15160 3756
rect 18002 3742 18016 3756
rect 19130 3742 19144 3756
rect 20978 3742 20992 3756
rect 23570 3742 23584 3756
rect 25178 3742 25192 3756
rect 25826 3742 25840 3756
rect 26378 3742 26392 3756
rect 2570 3718 2584 3732
rect 12770 3718 12784 3732
rect 12938 3718 12952 3732
rect 17642 3718 17656 3732
rect 21194 3718 21208 3732
rect 21410 3718 21424 3732
rect 21890 3718 21904 3732
rect 22130 3718 22144 3732
rect 2570 3694 2584 3708
rect 9962 3694 9976 3708
rect 22898 3694 22912 3708
rect 23594 3694 23608 3708
rect 27170 3694 27184 3708
rect 2594 3670 2608 3684
rect 14762 3670 14776 3684
rect 17354 3670 17368 3684
rect 17426 3670 17440 3684
rect 2618 3646 2632 3660
rect 24818 3646 24832 3660
rect 2810 3622 2824 3636
rect 19202 3622 19216 3636
rect 3146 3598 3160 3612
rect 21818 3598 21832 3612
rect 3194 3574 3208 3588
rect 18674 3574 18688 3588
rect 3218 3550 3232 3564
rect 5186 3550 5200 3564
rect 17762 3550 17776 3564
rect 25202 3550 25216 3564
rect 25274 3550 25288 3564
rect 25658 3550 25672 3564
rect 26882 3550 26896 3564
rect 3242 3526 3256 3540
rect 6002 3526 6016 3540
rect 6050 3526 6064 3540
rect 8738 3526 8752 3540
rect 8834 3526 8848 3540
rect 13970 3526 13984 3540
rect 14018 3526 14032 3540
rect 24770 3526 24784 3540
rect 3338 3502 3352 3516
rect 24434 3502 24448 3516
rect 24770 3502 24784 3516
rect 26570 3502 26584 3516
rect 27842 3502 27856 3516
rect 3386 3478 3400 3492
rect 5114 3478 5128 3492
rect 9002 3478 9016 3492
rect 15026 3478 15040 3492
rect 17282 3478 17296 3492
rect 19850 3478 19864 3492
rect 20762 3478 20776 3492
rect 21650 3478 21664 3492
rect 24062 3478 24076 3492
rect 27770 3478 27784 3492
rect 3434 3454 3448 3468
rect 5762 3454 5776 3468
rect 7442 3454 7456 3468
rect 12290 3454 12304 3468
rect 13754 3454 13768 3468
rect 23042 3454 23056 3468
rect 25538 3454 25552 3468
rect 3530 3430 3544 3444
rect 11234 3430 11248 3444
rect 25970 3430 25984 3444
rect 3578 3406 3592 3420
rect 15722 3406 15736 3420
rect 3578 3382 3592 3396
rect 6674 3382 6688 3396
rect 10322 3382 10336 3396
rect 12578 3382 12592 3396
rect 13202 3382 13216 3396
rect 18986 3382 19000 3396
rect 21290 3382 21304 3396
rect 22946 3382 22960 3396
rect 25010 3382 25024 3396
rect 3602 3358 3616 3372
rect 11498 3358 11512 3372
rect 21482 3358 21496 3372
rect 22946 3358 22960 3372
rect 22970 3358 22984 3372
rect 3650 3334 3664 3348
rect 8522 3334 8536 3348
rect 8834 3334 8848 3348
rect 9602 3334 9616 3348
rect 16154 3334 16168 3348
rect 3842 3310 3856 3324
rect 10250 3310 10264 3324
rect 10322 3310 10336 3324
rect 10370 3310 10384 3324
rect 11018 3310 11032 3324
rect 11282 3310 11296 3324
rect 11330 3310 11344 3324
rect 11426 3310 11440 3324
rect 11546 3310 11560 3324
rect 11714 3310 11728 3324
rect 11762 3310 11776 3324
rect 23066 3310 23080 3324
rect 3890 3286 3904 3300
rect 6314 3286 6328 3300
rect 8018 3286 8032 3300
rect 9914 3286 9928 3300
rect 16106 3286 16120 3300
rect 20618 3286 20632 3300
rect 3914 3262 3928 3276
rect 12890 3262 12904 3276
rect 19154 3262 19168 3276
rect 24314 3262 24328 3276
rect 25322 3262 25336 3276
rect 3962 3238 3976 3252
rect 11786 3238 11800 3252
rect 17114 3238 17128 3252
rect 19154 3238 19168 3252
rect 19334 3238 19348 3252
rect 4010 3214 4024 3228
rect 4994 3214 5008 3228
rect 8258 3214 8272 3228
rect 14138 3214 14152 3228
rect 14258 3214 14272 3228
rect 24626 3214 24640 3228
rect 4106 3190 4120 3204
rect 7154 3190 7168 3204
rect 17882 3190 17896 3204
rect 21074 3190 21088 3204
rect 23258 3190 23272 3204
rect 24734 3190 24748 3204
rect 25298 3190 25312 3204
rect 4154 3166 4168 3180
rect 12146 3166 12160 3180
rect 26330 3166 26344 3180
rect 4202 3142 4216 3156
rect 5906 3142 5920 3156
rect 12170 3142 12184 3156
rect 23138 3142 23152 3156
rect 26330 3142 26344 3156
rect 26402 3142 26416 3156
rect 4346 3118 4360 3132
rect 26642 3118 26656 3132
rect 4346 3094 4360 3108
rect 8546 3094 8560 3108
rect 8906 3094 8920 3108
rect 13178 3094 13192 3108
rect 18746 3094 18760 3108
rect 24386 3094 24400 3108
rect 25634 3094 25648 3108
rect 27314 3094 27328 3108
rect 4394 3070 4408 3084
rect 14306 3070 14320 3084
rect 14402 3070 14416 3084
rect 26210 3070 26224 3084
rect 4442 3046 4456 3060
rect 13274 3046 13288 3060
rect 13418 3046 13432 3060
rect 13802 3046 13816 3060
rect 4442 3022 4456 3036
rect 25154 3022 25168 3036
rect 4490 2998 4504 3012
rect 8354 2998 8368 3012
rect 9002 2998 9016 3012
rect 10754 2998 10768 3012
rect 11042 2998 11056 3012
rect 20594 2998 20608 3012
rect 4682 2974 4696 2988
rect 12986 2974 13000 2988
rect 13370 2974 13384 2988
rect 13514 2974 13528 2988
rect 14042 2974 14056 2988
rect 4802 2950 4816 2964
rect 9602 2950 9616 2964
rect 9650 2950 9664 2964
rect 13586 2950 13600 2964
rect 5042 2926 5056 2940
rect 21530 2926 21544 2940
rect 5426 2902 5440 2916
rect 10634 2902 10648 2916
rect 10754 2902 10768 2916
rect 12194 2902 12208 2916
rect 14906 2902 14920 2916
rect 23450 2902 23464 2916
rect 5474 2878 5488 2892
rect 14594 2878 14608 2892
rect 20738 2878 20752 2892
rect 22586 2878 22600 2892
rect 5522 2854 5536 2868
rect 25346 2854 25360 2868
rect 5666 2830 5680 2844
rect 14786 2830 14800 2844
rect 5978 2806 5992 2820
rect 17690 2806 17704 2820
rect 21506 2806 21520 2820
rect 6026 2782 6040 2796
rect 11402 2782 11416 2796
rect 20354 2782 20368 2796
rect 21506 2782 21520 2796
rect 21758 2782 21772 2796
rect 6074 2758 6088 2772
rect 15578 2758 15592 2772
rect 6122 2734 6136 2748
rect 6890 2734 6904 2748
rect 9986 2734 10000 2748
rect 23642 2734 23656 2748
rect 6170 2710 6184 2724
rect 13946 2710 13960 2724
rect 20210 2710 20224 2724
rect 27506 2710 27520 2724
rect 6218 2686 6232 2700
rect 17570 2686 17584 2700
rect 22082 2686 22096 2700
rect 24578 2686 24592 2700
rect 6338 2662 6352 2676
rect 13610 2662 13624 2676
rect 20210 2662 20224 2676
rect 20330 2662 20344 2676
rect 6602 2638 6616 2652
rect 12410 2638 12424 2652
rect 12578 2638 12592 2652
rect 12794 2638 12808 2652
rect 13178 2638 13192 2652
rect 13334 2638 13348 2652
rect 13538 2638 13552 2652
rect 19010 2638 19024 2652
rect 6770 2614 6784 2628
rect 6938 2614 6952 2628
rect 7058 2614 7072 2628
rect 7442 2614 7456 2628
rect 13562 2614 13576 2628
rect 16370 2614 16384 2628
rect 22994 2614 23008 2628
rect 6962 2590 6976 2604
rect 9086 2590 9100 2604
rect 10586 2590 10600 2604
rect 12242 2590 12256 2604
rect 13706 2590 13720 2604
rect 17498 2590 17512 2604
rect 20834 2590 20848 2604
rect 21218 2590 21232 2604
rect 21950 2590 21964 2604
rect 24218 2590 24232 2604
rect 25610 2590 25624 2604
rect 7082 2566 7096 2580
rect 7634 2566 7648 2580
rect 17594 2566 17608 2580
rect 7130 2542 7144 2556
rect 17306 2542 17320 2556
rect 17498 2542 17512 2556
rect 26138 2542 26152 2556
rect 7394 2518 7408 2532
rect 8306 2518 8320 2532
rect 12458 2518 12472 2532
rect 22754 2518 22768 2532
rect 23114 2518 23128 2532
rect 7466 2494 7480 2508
rect 28227 2494 28241 2508
rect 7706 2470 7720 2484
rect 9266 2470 9280 2484
rect 21002 2470 21016 2484
rect 25274 2470 25288 2484
rect 7802 2446 7816 2460
rect 13250 2446 13264 2460
rect 7946 2422 7960 2436
rect 20714 2422 20728 2436
rect 7994 2398 8008 2412
rect 11306 2398 11320 2412
rect 11378 2398 11392 2412
rect 11522 2398 11536 2412
rect 11594 2398 11608 2412
rect 19298 2398 19312 2412
rect 8042 2374 8056 2388
rect 21794 2374 21808 2388
rect 8042 2350 8056 2364
rect 8378 2350 8392 2364
rect 9074 2350 9088 2364
rect 9218 2350 9232 2364
rect 9266 2350 9280 2364
rect 9314 2350 9328 2364
rect 9506 2350 9520 2364
rect 23330 2350 23344 2364
rect 8138 2326 8152 2340
rect 26282 2326 26296 2340
rect 8162 2302 8176 2316
rect 24242 2302 24256 2316
rect 9170 2278 9184 2292
rect 9194 2278 9208 2292
rect 9290 2278 9304 2292
rect 11474 2278 11488 2292
rect 11666 2278 11680 2292
rect 20930 2278 20944 2292
rect 24242 2278 24256 2292
rect 24266 2278 24280 2292
rect 9626 2254 9640 2268
rect 19418 2254 19432 2268
rect 20930 2254 20944 2268
rect 21362 2254 21376 2268
rect 9698 2230 9712 2244
rect 27674 2230 27688 2244
rect 9866 2206 9880 2220
rect 20090 2206 20104 2220
rect 10034 2182 10048 2196
rect 20498 2182 20512 2196
rect 10154 2158 10168 2172
rect 14186 2158 14200 2172
rect 11186 2134 11200 2148
rect 27098 2134 27112 2148
rect 11282 2110 11296 2124
rect 26186 2110 26200 2124
rect 11450 2086 11464 2100
rect 12866 2086 12880 2100
rect 14186 2086 14200 2100
rect 17378 2086 17392 2100
rect 18530 2086 18544 2100
rect 24794 2086 24808 2100
rect 26114 2086 26128 2100
rect 11762 2062 11776 2076
rect 19610 2062 19624 2076
rect 27890 2062 27904 2076
rect 28227 2062 28241 2076
rect 11834 2038 11848 2052
rect 14978 2038 14992 2052
rect 24938 2038 24952 2052
rect 27866 2038 27880 2052
rect 28227 2038 28241 2052
rect 11978 2014 11992 2028
rect 12626 2014 12640 2028
rect 16874 2014 16888 2028
rect 27842 2014 27856 2028
rect 28227 2014 28241 2028
rect 12026 1990 12040 2004
rect 12086 1990 12100 2004
rect 12314 1990 12328 2004
rect 17666 1990 17680 2004
rect 27818 1990 27832 2004
rect 28227 1990 28241 2004
rect 12074 1966 12088 1980
rect 23018 1966 23032 1980
rect 27794 1966 27808 1980
rect 28227 1966 28241 1980
rect 12386 1942 12400 1956
rect 13778 1942 13792 1956
rect 27266 1942 27280 1956
rect 27770 1942 27784 1956
rect 28227 1942 28241 1956
rect 16250 1109 16264 1123
rect 21962 1109 21976 1123
rect 16202 1085 16216 1099
rect 18866 1085 18880 1099
rect 15986 1061 16000 1075
rect 22370 1061 22384 1075
rect 15890 1037 15904 1051
rect 16274 1037 16288 1051
rect 17234 1037 17248 1051
rect 19010 1037 19024 1051
rect 15794 1013 15808 1027
rect 22802 1013 22816 1027
rect 10418 989 10432 1003
rect 11666 989 11680 1003
rect 11714 989 11728 1003
rect 17858 989 17872 1003
rect 10370 965 10384 979
rect 17258 965 17272 979
rect 17474 965 17488 979
rect 22298 965 22312 979
rect 9674 941 9688 955
rect 25730 941 25744 955
rect 9338 917 9352 931
rect 12818 917 12832 931
rect 18050 917 18064 931
rect 21314 917 21328 931
rect 21938 917 21952 931
rect 26570 917 26584 931
rect 26810 917 26824 931
rect 9122 893 9136 907
rect 12410 893 12424 907
rect 17570 893 17584 907
rect 18626 893 18640 907
rect 24338 893 24352 907
rect 8426 869 8440 883
rect 13658 869 13672 883
rect 13778 869 13792 883
rect 18602 869 18616 883
rect 8306 845 8320 859
rect 20258 845 20272 859
rect 20306 845 20320 859
rect 25970 845 25984 859
rect 8090 821 8104 835
rect 25802 821 25816 835
rect 7298 797 7312 811
rect 9746 797 9760 811
rect 10058 797 10072 811
rect 11066 797 11080 811
rect 11474 797 11488 811
rect 14354 797 14368 811
rect 14930 797 14944 811
rect 21098 797 21112 811
rect 6866 773 6880 787
rect 6938 773 6952 787
rect 7202 773 7216 787
rect 18650 773 18664 787
rect 19058 773 19072 787
rect 22706 773 22720 787
rect 6818 749 6832 763
rect 16562 749 16576 763
rect 21170 749 21184 763
rect 24386 749 24400 763
rect 6746 725 6760 739
rect 7322 725 7336 739
rect 23618 725 23632 739
rect 6722 701 6736 715
rect 13346 701 13360 715
rect 13442 701 13456 715
rect 17594 701 17608 715
rect 17666 701 17680 715
rect 21242 701 21256 715
rect 21746 701 21760 715
rect 23522 701 23536 715
rect 6506 677 6520 691
rect 17906 677 17920 691
rect 18026 677 18040 691
rect 21914 677 21928 691
rect 24122 677 24136 691
rect 6338 653 6352 667
rect 10778 653 10792 667
rect 12842 653 12856 667
rect 22130 653 22144 667
rect 23498 653 23512 667
rect 24002 653 24016 667
rect 26762 653 26776 667
rect 6266 629 6280 643
rect 10994 629 11008 643
rect 11042 629 11056 643
rect 24722 629 24736 643
rect 5954 605 5968 619
rect 22778 605 22792 619
rect 24626 605 24640 619
rect 5882 581 5896 595
rect 7658 581 7672 595
rect 8066 581 8080 595
rect 12146 581 12160 595
rect 26834 581 26848 595
rect 5786 557 5800 571
rect 22898 557 22912 571
rect 4946 533 4960 547
rect 23690 533 23704 547
rect 4922 509 4936 523
rect 6554 509 6568 523
rect 19106 509 19120 523
rect 4802 485 4816 499
rect 7178 485 7192 499
rect 10826 485 10840 499
rect 11522 485 11536 499
rect 20090 485 20104 499
rect 20498 485 20512 499
rect 4730 461 4744 475
rect 23162 461 23176 475
rect 4658 437 4672 451
rect 11090 437 11104 451
rect 11858 437 11872 451
rect 20138 437 20152 451
rect 4586 413 4600 427
rect 19346 413 19360 427
rect 4394 389 4408 403
rect 25418 389 25432 403
rect 4322 365 4336 379
rect 25850 365 25864 379
rect 4058 341 4072 355
rect 11426 341 11440 355
rect 11882 341 11896 355
rect 13946 341 13960 355
rect 14066 341 14080 355
rect 23042 341 23056 355
rect 4034 317 4048 331
rect 18482 317 18496 331
rect 21410 317 21424 331
rect 26858 317 26872 331
rect 3818 293 3832 307
rect 21890 293 21904 307
rect 26786 293 26800 307
rect 3746 269 3760 283
rect 10442 269 10456 283
rect 10610 269 10624 283
rect 21770 269 21784 283
rect 3506 245 3520 259
rect 21026 245 21040 259
rect 3362 221 3376 235
rect 20810 221 20824 235
rect 26714 221 26746 235
rect 2810 197 2824 211
rect 18914 197 18928 211
rect 2690 173 2704 187
rect 13634 173 13648 187
rect 15050 173 15064 187
rect 26618 173 26632 187
rect 2666 149 2680 163
rect 17042 149 17056 163
rect 17282 149 17296 163
rect 21122 149 21136 163
rect 1706 125 1720 139
rect 19898 125 19912 139
rect 26726 125 26740 139
rect 28227 125 28241 139
rect 1634 101 1648 115
rect 20834 101 20848 115
rect 26858 101 26872 115
rect 28227 101 28241 115
rect 70 77 84 91
rect 22274 77 22288 91
rect 26834 77 26848 91
rect 28227 77 28241 91
rect 70 53 84 67
rect 1754 53 1768 67
rect 2642 53 2656 67
rect 16682 53 16696 67
rect 19754 53 19768 67
rect 26810 53 26824 67
rect 28227 53 28241 67
rect 70 29 84 43
rect 12578 29 12592 43
rect 12626 29 12640 43
rect 19946 29 19960 43
rect 26786 29 26800 43
rect 28227 29 28241 43
rect 70 5 84 19
rect 16442 5 16456 19
rect 26762 5 26776 19
rect 28227 5 28241 19
<< metal2 >>
rect 0 8632 70 8644
rect 0 8608 70 8620
rect 0 8584 70 8596
rect 123 8429 323 8799
rect 339 8429 351 8799
rect 363 8429 375 8799
rect 387 8429 399 8799
rect 411 8429 423 8799
rect 1707 8429 1719 8607
rect 1755 8429 1767 8583
rect 2859 8429 2871 8607
rect 3111 8597 3123 8799
rect 4659 8573 4671 8799
rect 4695 8621 4707 8799
rect 7143 8669 7155 8799
rect 7144 8655 7162 8669
rect 6939 8429 6951 8607
rect 7083 8429 7095 8535
rect 7131 8429 7143 8655
rect 8751 8573 8763 8799
rect 10851 8669 10863 8799
rect 12255 8693 12267 8799
rect 12256 8679 12274 8693
rect 8752 8559 8770 8573
rect 7827 8429 7839 8559
rect 8739 8429 8751 8559
rect 9219 8429 9231 8583
rect 10347 8429 10359 8583
rect 11091 8429 11103 8559
rect 12243 8429 12255 8679
rect 12675 8429 12687 8679
rect 13035 8429 13047 8703
rect 13371 8429 13383 8727
rect 13947 8525 13959 8799
rect 15495 8501 15507 8799
rect 16827 8429 16839 8463
rect 16923 8429 16935 8751
rect 17031 8453 17043 8799
rect 17055 8717 17067 8799
rect 18675 8429 18687 8703
rect 18819 8429 18831 8775
rect 20103 8669 20115 8799
rect 20127 8741 20139 8799
rect 21663 8693 21675 8799
rect 23199 8765 23211 8799
rect 24735 8789 24747 8799
rect 18867 8429 18879 8655
rect 22851 8429 22863 8439
rect 23187 8429 23199 8511
rect 23835 8429 23847 8655
rect 25563 8429 25575 8487
rect 25779 8429 25791 8631
rect 26271 8573 26283 8799
rect 27843 8597 27855 8703
rect 27723 8429 27735 8559
rect 27771 8429 27783 8511
rect 27795 8501 27807 8511
rect 27819 8477 27831 8583
rect 27867 8549 27879 8607
rect 27843 8525 27855 8535
rect 27795 8453 27807 8463
rect 27915 8429 28115 8799
rect 28241 8584 28311 8596
rect 28241 8560 28311 8572
rect 28241 8536 28311 8548
rect 28241 8512 28311 8524
rect 28241 8488 28311 8500
rect 28241 8464 28311 8476
rect 28241 8440 28311 8452
rect 0 4103 70 4115
rect 0 4079 70 4091
rect 0 4055 70 4067
rect 0 4031 70 4043
rect 123 1932 323 7630
rect 339 1932 351 7630
rect 363 1932 375 7630
rect 387 1932 399 7630
rect 411 1932 423 7630
rect 1611 4140 1623 7630
rect 1635 4164 1647 7630
rect 1659 4188 1671 7630
rect 1611 1932 1623 4006
rect 1659 1932 1671 3982
rect 1683 1932 1695 4198
rect 1707 3972 1719 7630
rect 1755 4260 1767 7630
rect 1803 4284 1815 7630
rect 1827 4308 1839 7630
rect 1755 1932 1767 4222
rect 1851 3948 1863 7630
rect 1899 4356 1911 7630
rect 1923 4380 1935 7630
rect 1875 1932 1887 4318
rect 1947 3924 1959 7630
rect 1995 4404 2007 7630
rect 2019 4428 2031 7630
rect 2043 4452 2055 7630
rect 2067 3900 2079 7630
rect 2091 4116 2103 7630
rect 2139 4116 2151 7630
rect 2163 4476 2175 7630
rect 2187 4500 2199 7630
rect 2235 4524 2247 7630
rect 2259 4548 2271 7630
rect 2283 3876 2295 7630
rect 2307 4572 2319 7630
rect 2355 4596 2367 7630
rect 2379 4620 2391 7630
rect 2427 4644 2439 7630
rect 2475 4668 2487 7630
rect 2499 4692 2511 7630
rect 2523 4716 2535 7630
rect 2235 1932 2247 3862
rect 2283 1932 2295 3838
rect 2427 1932 2439 3814
rect 2451 1932 2463 3790
rect 2475 1932 2487 3766
rect 2523 1932 2535 3742
rect 2547 1932 2559 3790
rect 2571 3732 2583 7630
rect 2595 4740 2607 7630
rect 2571 1932 2583 3694
rect 2595 1932 2607 3670
rect 2619 3660 2631 7630
rect 2643 4764 2655 7630
rect 2691 4788 2703 7630
rect 2715 4812 2727 7630
rect 2739 4836 2751 7630
rect 2787 4860 2799 7630
rect 2811 3636 2823 7630
rect 2835 4884 2847 7630
rect 2907 4908 2919 7630
rect 2931 4932 2943 7630
rect 2955 4956 2967 7630
rect 3003 4980 3015 7630
rect 3027 5004 3039 7630
rect 3051 5028 3063 7630
rect 3099 4596 3111 7630
rect 3123 5052 3135 7630
rect 3147 3612 3159 7630
rect 3171 1932 3183 4774
rect 3195 3588 3207 7630
rect 3219 1932 3231 3550
rect 3243 3540 3255 7630
rect 3315 4116 3327 7630
rect 3339 3516 3351 7630
rect 3387 5076 3399 7630
rect 3435 5100 3447 7630
rect 3459 5124 3471 7630
rect 3483 5148 3495 7630
rect 3531 5172 3543 7630
rect 3555 5196 3567 7630
rect 3387 1932 3399 3478
rect 3435 1932 3447 3454
rect 3483 1932 3495 4486
rect 3531 1932 3543 3430
rect 3579 3420 3591 7630
rect 3627 5220 3639 7630
rect 3651 4668 3663 7630
rect 3675 5244 3687 7630
rect 3723 5292 3735 7630
rect 3747 5316 3759 7630
rect 3771 5340 3783 7630
rect 3819 5364 3831 7630
rect 3843 5388 3855 7630
rect 3867 5412 3879 7630
rect 3579 1932 3591 3382
rect 3603 1932 3615 3358
rect 3627 1932 3639 3862
rect 3651 1932 3663 3334
rect 3699 1932 3711 5254
rect 3915 5196 3927 7630
rect 3939 5292 3951 7630
rect 3963 5436 3975 7630
rect 3987 5460 3999 7630
rect 4035 5484 4047 7630
rect 4083 4980 4095 7630
rect 4155 4980 4167 7630
rect 4179 5508 4191 7630
rect 4203 5532 4215 7630
rect 4251 5556 4263 7630
rect 3723 1932 3735 3790
rect 3795 1932 3807 4102
rect 3843 1932 3855 3310
rect 3891 1932 3903 3286
rect 3915 1932 3927 3262
rect 3963 1932 3975 3238
rect 4011 1932 4023 3214
rect 4107 1932 4119 3190
rect 4131 1932 4143 4702
rect 4155 1932 4167 3166
rect 4203 1932 4215 3142
rect 4251 1932 4263 4966
rect 4275 3852 4287 7630
rect 4299 5580 4311 7630
rect 4347 3132 4359 7630
rect 4371 5604 4383 7630
rect 4347 1932 4359 3094
rect 4395 3084 4407 7630
rect 4419 5628 4431 7630
rect 4443 3060 4455 7630
rect 4491 5652 4503 7630
rect 4443 1932 4455 3022
rect 4467 1932 4479 5494
rect 4515 4932 4527 7630
rect 4539 5508 4551 7630
rect 4563 5676 4575 7630
rect 4587 4068 4599 7630
rect 4635 5700 4647 7630
rect 4659 5724 4671 7630
rect 4683 5748 4695 7630
rect 4491 1932 4503 2998
rect 4539 1932 4551 4054
rect 4707 4020 4719 7630
rect 4755 4260 4767 7630
rect 4683 1932 4695 2974
rect 4779 1932 4791 4006
rect 4803 2964 4815 7630
rect 4875 5796 4887 7630
rect 4923 5820 4935 7630
rect 4851 1932 4863 5758
rect 4899 1932 4911 4126
rect 4995 3228 5007 7630
rect 5019 5844 5031 7630
rect 5043 2940 5055 7630
rect 5091 5892 5103 7630
rect 5067 1932 5079 5854
rect 5115 3492 5127 7630
rect 5139 5916 5151 7630
rect 5187 3564 5199 7630
rect 5211 5844 5223 7630
rect 5235 5940 5247 7630
rect 5283 5508 5295 7630
rect 5307 5964 5319 7630
rect 5331 5988 5343 7630
rect 5355 5748 5367 7630
rect 5379 6012 5391 7630
rect 5427 6036 5439 7630
rect 5451 6060 5463 7630
rect 5475 6084 5487 7630
rect 5427 1932 5439 2902
rect 5475 1932 5487 2878
rect 5523 2868 5535 7630
rect 5571 6036 5583 7630
rect 5619 1932 5631 5038
rect 5643 4788 5655 7630
rect 5667 6108 5679 7630
rect 5691 4812 5703 7630
rect 5715 6132 5727 7630
rect 5763 6156 5775 7630
rect 5643 1932 5655 4150
rect 5667 1932 5679 2830
rect 5715 1932 5727 5806
rect 5787 4836 5799 7630
rect 5811 6180 5823 7630
rect 5859 6204 5871 7630
rect 5739 1932 5751 3790
rect 5763 1932 5775 3454
rect 5835 1932 5847 4462
rect 5859 1932 5871 5278
rect 5907 4908 5919 7630
rect 5979 4836 5991 7630
rect 5883 1932 5895 4654
rect 6003 3852 6015 7630
rect 6027 6228 6039 7630
rect 5907 1932 5919 3142
rect 5979 1932 5991 2806
rect 6003 1932 6015 3526
rect 6027 1932 6039 2782
rect 6051 1932 6063 3526
rect 6075 2772 6087 7630
rect 6099 6252 6111 7630
rect 6123 6276 6135 7630
rect 6171 4524 6183 7630
rect 6099 1932 6111 4510
rect 6195 3852 6207 7630
rect 6243 4596 6255 7630
rect 6291 4260 6303 7630
rect 6315 6300 6327 7630
rect 6123 1932 6135 2734
rect 6171 1932 6183 2710
rect 6219 1932 6231 2686
rect 6243 1932 6255 4246
rect 6315 1932 6327 3286
rect 6339 2676 6351 7630
rect 6387 6324 6399 7630
rect 6459 6348 6471 7630
rect 6531 6372 6543 7630
rect 6603 6396 6615 7630
rect 6627 6156 6639 7630
rect 6651 6420 6663 7630
rect 6675 5268 6687 7630
rect 6723 5268 6735 7630
rect 6747 6156 6759 7630
rect 6771 6444 6783 7630
rect 6387 1932 6399 4006
rect 6435 1932 6447 5110
rect 6459 1932 6471 5038
rect 6819 4908 6831 7630
rect 6843 6468 6855 7630
rect 6483 1932 6495 3838
rect 6603 1932 6615 2638
rect 6675 1932 6687 3382
rect 6699 1932 6711 4486
rect 6891 2748 6903 7630
rect 6939 2628 6951 7630
rect 6987 6492 6999 7630
rect 6771 1932 6783 2614
rect 6963 1932 6975 2590
rect 6987 1932 6999 6046
rect 7011 4860 7023 7630
rect 7035 6516 7047 7630
rect 7035 1932 7047 4678
rect 7059 2628 7071 7630
rect 7083 1932 7095 2566
rect 7131 2556 7143 7630
rect 7179 6540 7191 7630
rect 7227 5052 7239 7630
rect 7299 6588 7311 7630
rect 7323 6612 7335 7630
rect 7347 6636 7359 7630
rect 7371 6660 7383 7630
rect 7155 1932 7167 3190
rect 7251 1932 7263 5542
rect 7275 1932 7287 6550
rect 7395 3972 7407 7630
rect 7347 1932 7359 3958
rect 7395 1932 7407 2518
rect 7419 1932 7431 5446
rect 7443 3468 7455 7630
rect 7491 6684 7503 7630
rect 7443 1932 7455 2614
rect 7467 1932 7479 2494
rect 7515 1932 7527 5830
rect 7539 1932 7551 6454
rect 7563 4644 7575 7630
rect 7587 6708 7599 7630
rect 7611 6732 7623 7630
rect 7659 6708 7671 7630
rect 7587 1932 7599 4102
rect 7611 3804 7623 6694
rect 7683 5388 7695 7630
rect 7707 6756 7719 7630
rect 7755 6780 7767 7630
rect 7779 6804 7791 7630
rect 7803 6828 7815 7630
rect 7875 6852 7887 7630
rect 7635 1932 7647 2566
rect 7707 1932 7719 2470
rect 7755 1932 7767 3742
rect 7779 1932 7791 3862
rect 7803 1932 7815 2446
rect 7851 1932 7863 5038
rect 7875 1932 7887 6694
rect 7899 5652 7911 7630
rect 7947 3900 7959 7630
rect 7995 6876 8007 7630
rect 7899 1932 7911 3886
rect 7947 1932 7959 2422
rect 7971 1932 7983 5494
rect 8019 3300 8031 7630
rect 7995 1932 8007 2398
rect 8043 2388 8055 7630
rect 8091 6900 8103 7630
rect 8115 6924 8127 7630
rect 8139 6948 8151 7630
rect 8163 6972 8175 7630
rect 8187 6996 8199 7630
rect 8043 1932 8055 2350
rect 8139 1932 8151 2326
rect 8163 1932 8175 2302
rect 8211 1932 8223 7006
rect 8235 4548 8247 7630
rect 8259 6924 8271 7630
rect 8283 7044 8295 7630
rect 8259 1932 8271 3214
rect 8283 1932 8295 5110
rect 8307 2532 8319 7030
rect 8331 3876 8343 7630
rect 8355 3012 8367 7630
rect 8379 2364 8391 7630
rect 8427 7044 8439 7630
rect 8451 4236 8463 7630
rect 8475 4740 8487 7630
rect 8523 3348 8535 7630
rect 8547 3108 8559 7630
rect 8571 4740 8583 7630
rect 8619 3852 8631 7630
rect 8643 5100 8655 7630
rect 8667 5844 8679 7630
rect 8691 4236 8703 7630
rect 8739 3540 8751 7630
rect 8787 5484 8799 7630
rect 8811 4788 8823 7630
rect 8835 3540 8847 7630
rect 8883 3804 8895 7630
rect 8835 1932 8847 3334
rect 8907 3108 8919 7630
rect 8931 6540 8943 7630
rect 8979 7068 8991 7630
rect 8979 1932 8991 6070
rect 9003 3492 9015 7630
rect 9051 7092 9063 7630
rect 9099 7116 9111 7630
rect 9003 1932 9015 2998
rect 9027 1932 9039 6790
rect 9051 1932 9063 4870
rect 9087 2604 9099 7054
rect 9123 6708 9135 7630
rect 9147 3804 9159 7630
rect 9171 4884 9183 7630
rect 9075 1932 9087 2350
rect 9195 2292 9207 5086
rect 9219 2364 9231 7630
rect 9171 1932 9183 2278
rect 9243 1932 9255 4054
rect 9267 2484 9279 7630
rect 9291 4908 9303 7630
rect 9315 2364 9327 7630
rect 9267 1932 9279 2350
rect 9291 1932 9303 2278
rect 9339 1932 9351 5638
rect 9363 4620 9375 7630
rect 9387 4884 9399 7630
rect 9411 6924 9423 7630
rect 9435 7068 9447 7630
rect 9459 7140 9471 7630
rect 9387 1932 9399 4462
rect 9459 1932 9471 7030
rect 9483 3804 9495 4870
rect 9507 4788 9519 7630
rect 9531 4620 9543 7630
rect 9555 6420 9567 7630
rect 9507 1932 9519 2350
rect 9579 1932 9591 4366
rect 9603 3348 9615 7630
rect 9627 4884 9639 7630
rect 9651 2964 9663 7630
rect 9699 5940 9711 7630
rect 9747 6708 9759 7630
rect 9819 7164 9831 7630
rect 9843 7188 9855 7630
rect 9867 7212 9879 7630
rect 9915 7236 9927 7630
rect 9939 7260 9951 7630
rect 9603 1932 9615 2950
rect 9627 1932 9639 2254
rect 9699 1932 9711 2230
rect 9795 1932 9807 3862
rect 9819 1932 9831 4462
rect 9867 1932 9879 2206
rect 9915 1932 9927 3286
rect 9939 1932 9951 5494
rect 9963 5004 9975 7630
rect 10011 7284 10023 7630
rect 9963 1932 9975 3694
rect 9987 2748 9999 7246
rect 10011 1932 10023 5278
rect 10035 5004 10047 7630
rect 10059 7260 10071 7630
rect 10083 4212 10095 7630
rect 10035 1932 10047 2182
rect 10107 1932 10119 5086
rect 10131 4716 10143 7630
rect 10155 4212 10167 5302
rect 10179 4932 10191 7630
rect 10131 1932 10143 4198
rect 10155 1932 10167 2158
rect 10203 1932 10215 5302
rect 10227 1932 10239 4462
rect 10251 3324 10263 7630
rect 10275 7308 10287 7630
rect 10299 7020 10311 7630
rect 10275 1932 10287 4606
rect 10323 3396 10335 7630
rect 10395 6444 10407 7630
rect 10323 1932 10335 3310
rect 10347 1932 10359 5494
rect 10419 5052 10431 7630
rect 10443 6444 10455 7630
rect 10491 7020 10503 7630
rect 10371 3324 10383 3886
rect 10467 1932 10479 4198
rect 10491 1932 10503 4078
rect 10515 3900 10527 7630
rect 10539 7332 10551 7630
rect 10563 7356 10575 7630
rect 10539 1932 10551 4510
rect 10563 1932 10575 4342
rect 10611 4092 10623 7630
rect 10635 2916 10647 7630
rect 10659 7284 10671 7630
rect 10707 7380 10719 7630
rect 10587 1932 10599 2590
rect 10659 1932 10671 3910
rect 10683 1932 10695 6430
rect 10707 1932 10719 4030
rect 10755 3012 10767 7630
rect 10827 5988 10839 7630
rect 10851 5964 10863 7630
rect 10875 5628 10887 7630
rect 10923 6996 10935 7630
rect 10947 6444 10959 7630
rect 10755 1932 10767 2902
rect 10875 1932 10887 4030
rect 10899 1932 10911 4942
rect 10947 1932 10959 6334
rect 10971 5628 10983 7630
rect 11019 3924 11031 7630
rect 11019 1932 11031 3310
rect 11043 3012 11055 7630
rect 11067 7404 11079 7630
rect 11139 7116 11151 7630
rect 11163 5988 11175 7630
rect 11187 7428 11199 7630
rect 11235 7452 11247 7630
rect 11259 7476 11271 7630
rect 11139 1932 11151 3790
rect 11163 1932 11175 3838
rect 11187 1932 11199 2134
rect 11235 1932 11247 3430
rect 11259 1932 11271 5494
rect 11283 3324 11295 7630
rect 11307 2412 11319 7462
rect 11331 4524 11343 7630
rect 11355 6108 11367 7630
rect 11379 5316 11391 7630
rect 11283 1932 11295 2110
rect 11331 1932 11343 3310
rect 11355 1932 11367 4774
rect 11403 2796 11415 7630
rect 11427 3324 11439 5830
rect 11451 4284 11463 7630
rect 11379 1932 11391 2398
rect 11475 2292 11487 7630
rect 11499 3372 11511 7630
rect 11523 2412 11535 6142
rect 11547 5292 11559 7630
rect 11571 7476 11583 7630
rect 11451 1932 11463 2086
rect 11547 1932 11559 3310
rect 11571 1932 11583 4798
rect 11595 2412 11607 7630
rect 11643 7500 11655 7630
rect 11619 1932 11631 4534
rect 11643 1932 11655 4774
rect 11667 2292 11679 7630
rect 11691 6852 11703 7630
rect 11715 7524 11727 7630
rect 11715 3324 11727 6958
rect 11739 1932 11751 3742
rect 11763 3324 11775 7630
rect 11787 7548 11799 7630
rect 11787 3252 11799 7462
rect 11763 1932 11775 2062
rect 11811 1932 11823 5038
rect 11835 3996 11847 7630
rect 11883 7476 11895 7630
rect 11907 4956 11919 7630
rect 11835 1932 11847 2038
rect 11931 1932 11943 6022
rect 11955 4548 11967 7630
rect 11979 3996 11991 5182
rect 12003 4620 12015 7630
rect 11955 1932 11967 3982
rect 12027 3804 12039 7630
rect 12051 6924 12063 7630
rect 12075 5820 12087 7630
rect 12099 7572 12111 7630
rect 11979 1932 11991 2014
rect 12027 1932 12039 1990
rect 12051 1932 12063 3982
rect 12087 2004 12099 4990
rect 12075 1932 12087 1966
rect 12123 1932 12135 4678
rect 12147 3180 12159 7630
rect 12171 3156 12183 7630
rect 12195 7596 12207 7630
rect 12219 4884 12231 7630
rect 12195 1932 12207 2902
rect 12243 1932 12255 2590
rect 12267 1932 12279 6910
rect 12291 5292 12303 7630
rect 12315 4932 12327 7630
rect 12339 6852 12351 7630
rect 12387 4068 12399 7630
rect 12291 1932 12303 3454
rect 12315 1932 12327 1990
rect 12363 1932 12375 3790
rect 12411 2652 12423 7630
rect 12435 4932 12447 7630
rect 12459 4308 12471 7630
rect 12483 3996 12495 7270
rect 12507 5364 12519 7630
rect 12531 6156 12543 7630
rect 12387 1932 12399 1942
rect 12459 1932 12471 2518
rect 12507 1932 12519 4294
rect 12579 3396 12591 7630
rect 12579 1932 12591 2638
rect 12627 2028 12639 7630
rect 12651 7572 12663 7630
rect 12723 7044 12735 7630
rect 12747 7284 12759 7630
rect 12771 7572 12783 7630
rect 12651 1932 12663 4870
rect 12675 1932 12687 4054
rect 12723 1932 12735 6982
rect 12747 1932 12759 4078
rect 12771 1932 12783 3718
rect 12795 2652 12807 7270
rect 12819 3756 12831 7630
rect 12843 7284 12855 7630
rect 12843 1932 12855 7270
rect 12867 2100 12879 7630
rect 12915 3996 12927 7630
rect 12963 7596 12975 7630
rect 13035 7140 13047 7630
rect 13083 7596 13095 7630
rect 13107 7620 13119 7630
rect 13131 7164 13143 7630
rect 12891 1932 12903 3262
rect 12939 1932 12951 3718
rect 12963 1932 12975 7126
rect 12987 1932 12999 2974
rect 13035 1932 13047 5686
rect 13059 1932 13071 4894
rect 13083 1932 13095 5278
rect 13107 1932 13119 5806
rect 13131 1932 13143 6478
rect 13155 4068 13167 7126
rect 13179 3108 13191 7630
rect 13203 3876 13215 7630
rect 13227 7116 13239 7630
rect 13179 1932 13191 2638
rect 13203 1932 13215 3382
rect 13227 1932 13239 6958
rect 13251 2460 13263 7582
rect 13275 6684 13287 7630
rect 13299 4692 13311 7630
rect 13323 6684 13335 7630
rect 13275 1932 13287 3046
rect 13299 1932 13311 4054
rect 13335 2652 13347 6454
rect 13371 2988 13383 7630
rect 13419 5388 13431 7630
rect 13443 5988 13455 7630
rect 13467 7140 13479 7630
rect 13515 5100 13527 7630
rect 13539 6708 13551 7630
rect 13395 1932 13407 3790
rect 13419 1932 13431 3046
rect 13491 1932 13503 5038
rect 13515 1932 13527 2974
rect 13539 1932 13551 2638
rect 13563 2628 13575 7630
rect 13611 4716 13623 7630
rect 13635 5676 13647 7630
rect 13659 7164 13671 7630
rect 13707 7116 13719 7630
rect 13755 5388 13767 7630
rect 13671 4068 13683 5062
rect 13587 1932 13599 2950
rect 13611 1932 13623 2662
rect 13707 1932 13719 2590
rect 13731 1932 13743 5158
rect 13755 1932 13767 3454
rect 13779 1956 13791 7606
rect 13827 7596 13839 7630
rect 13803 3060 13815 7054
rect 13827 1932 13839 6670
rect 13851 4572 13863 7630
rect 13851 1932 13863 4054
rect 13875 1932 13887 4918
rect 13899 4860 13911 7630
rect 13923 1932 13935 6118
rect 13947 2724 13959 7630
rect 13971 5796 13983 7630
rect 13971 1932 13983 3526
rect 13995 1932 14007 4222
rect 14019 3828 14031 7630
rect 14019 1932 14031 3526
rect 14043 2988 14055 5830
rect 14067 5388 14079 7630
rect 14091 4860 14103 7630
rect 14091 1932 14103 3838
rect 14115 1932 14127 4702
rect 14139 3228 14151 7630
rect 14163 1932 14175 4558
rect 14187 2172 14199 7630
rect 14211 4692 14223 7630
rect 14259 5484 14271 7630
rect 14187 1932 14199 2086
rect 14211 1932 14223 4222
rect 14235 4068 14247 4894
rect 14307 4860 14319 7630
rect 14331 5844 14343 7630
rect 14343 3804 14355 4846
rect 14379 4284 14391 7630
rect 14427 6468 14439 7630
rect 14451 5652 14463 7630
rect 14499 4164 14511 7630
rect 14547 5412 14559 7630
rect 14571 5988 14583 7630
rect 14595 4860 14607 7630
rect 14259 1932 14271 3214
rect 14283 1932 14295 3742
rect 14307 1932 14319 3070
rect 14379 1932 14391 4054
rect 14403 1932 14415 3070
rect 14451 1932 14463 4150
rect 14475 1932 14487 3838
rect 14499 1932 14511 3742
rect 14523 1932 14535 4678
rect 14547 1932 14559 4270
rect 14619 4068 14631 6454
rect 14643 4932 14655 7630
rect 14667 5244 14679 7630
rect 14715 6948 14727 7630
rect 14691 4068 14703 6334
rect 14595 1932 14607 2878
rect 14667 1932 14679 4054
rect 14739 1932 14751 4558
rect 14763 3684 14775 7630
rect 14787 2844 14799 7630
rect 14811 6012 14823 7630
rect 14835 6132 14847 7630
rect 14835 1932 14847 5494
rect 14859 5244 14871 7630
rect 14907 5412 14919 7630
rect 14931 5052 14943 7630
rect 14859 1932 14871 4054
rect 14955 4044 14967 7630
rect 14907 1932 14919 2902
rect 14979 2052 14991 5398
rect 15003 5100 15015 7630
rect 15027 4596 15039 7630
rect 15051 5316 15063 7630
rect 15075 6660 15087 7630
rect 15123 6108 15135 7630
rect 15003 1932 15015 4102
rect 15147 3756 15159 7630
rect 15195 5412 15207 7630
rect 15315 4764 15327 7630
rect 15675 5484 15687 7630
rect 15027 1932 15039 3478
rect 15171 1932 15183 4102
rect 15531 1932 15543 4246
rect 15723 4092 15735 7630
rect 15867 6012 15879 7630
rect 15891 7572 15903 7630
rect 15579 1932 15591 2758
rect 15723 1932 15735 3406
rect 15747 1932 15759 4750
rect 15843 1932 15855 4006
rect 15867 1932 15879 4462
rect 15915 4236 15927 7630
rect 15939 5868 15951 7630
rect 15939 1932 15951 4246
rect 15963 1932 15975 6406
rect 15987 5676 15999 7630
rect 16011 4260 16023 6142
rect 16035 5868 16047 7630
rect 16179 5868 16191 7630
rect 16035 1932 16047 4366
rect 16059 1932 16071 4606
rect 16083 1932 16095 5254
rect 16107 3300 16119 5854
rect 16131 1932 16143 4246
rect 16155 1932 16167 3334
rect 16179 1932 16191 5374
rect 16299 1932 16311 5206
rect 16347 1932 16359 5446
rect 16371 1932 16383 2614
rect 16395 1932 16407 4222
rect 16443 1932 16455 4030
rect 16491 1932 16503 5686
rect 16515 1932 16527 7246
rect 16539 3804 16551 7630
rect 16587 5988 16599 7630
rect 16731 7044 16743 7630
rect 16755 4044 16767 7630
rect 16779 3900 16791 7630
rect 16827 4236 16839 7630
rect 16875 2028 16887 7630
rect 16995 4380 17007 7630
rect 17019 5100 17031 7630
rect 17043 5436 17055 7630
rect 17067 7404 17079 7630
rect 17091 1932 17103 6286
rect 17115 3252 17127 7630
rect 17139 5292 17151 7630
rect 17163 4668 17175 7630
rect 17187 5220 17199 7630
rect 17235 4668 17247 7630
rect 17259 5052 17271 7630
rect 17283 3492 17295 7630
rect 17307 7308 17319 7630
rect 17355 3828 17367 7630
rect 17379 5052 17391 7630
rect 17403 6588 17415 7630
rect 17307 1932 17319 2542
rect 17355 1932 17367 3670
rect 17379 1932 17391 2086
rect 17403 1932 17415 4222
rect 17427 3684 17439 6358
rect 17451 5748 17463 7630
rect 17451 1932 17463 5614
rect 17475 4236 17487 7318
rect 17499 2604 17511 7630
rect 17499 1932 17511 2542
rect 17523 1932 17535 4222
rect 17571 2700 17583 7630
rect 17595 2580 17607 7630
rect 17619 7308 17631 7630
rect 17619 1932 17631 7222
rect 17643 3732 17655 7294
rect 17667 2004 17679 7630
rect 17691 5268 17703 7630
rect 17715 5460 17727 7630
rect 17691 1932 17703 2806
rect 17739 1932 17751 6790
rect 17763 3564 17775 7630
rect 17787 5844 17799 7630
rect 17787 1932 17799 4030
rect 17811 1932 17823 5974
rect 17835 4524 17847 7630
rect 17859 4044 17871 7150
rect 17835 1932 17847 3886
rect 17883 3204 17895 7630
rect 17907 5628 17919 7630
rect 17931 6300 17943 7630
rect 17979 7116 17991 7630
rect 17955 1932 17967 4030
rect 18003 3756 18015 7630
rect 18027 6420 18039 7630
rect 18039 3900 18051 5494
rect 18075 4524 18087 7630
rect 18099 5388 18111 7630
rect 18147 6924 18159 7630
rect 18075 1932 18087 3886
rect 18123 1932 18135 6094
rect 18147 1932 18159 6694
rect 18171 1932 18183 6814
rect 18195 3900 18207 5614
rect 18219 1932 18231 6070
rect 18267 4236 18279 7630
rect 18675 6444 18687 7630
rect 18267 1932 18279 3886
rect 18339 1932 18351 4222
rect 18387 1932 18399 4870
rect 18459 1932 18471 4294
rect 18483 1932 18495 5734
rect 18531 1932 18543 2086
rect 18579 1932 18591 5206
rect 18675 1932 18687 3574
rect 18723 1932 18735 4534
rect 18747 1932 18759 3094
rect 18795 1932 18807 4342
rect 18819 4044 18831 7630
rect 18843 1932 18855 4534
rect 18867 3900 18879 7630
rect 18915 5580 18927 7630
rect 18891 1932 18903 5350
rect 18939 4740 18951 7630
rect 18963 5220 18975 7630
rect 18987 5580 18999 7630
rect 18963 1932 18975 4966
rect 18987 1932 18999 3382
rect 19011 2652 19023 5206
rect 19035 5028 19047 7630
rect 19059 4596 19071 7630
rect 19083 6780 19095 7630
rect 19107 4740 19119 6958
rect 19083 1932 19095 4726
rect 19131 3756 19143 7630
rect 19155 3276 19167 7630
rect 19179 6132 19191 7630
rect 19227 6300 19239 7630
rect 19251 5028 19263 7630
rect 19275 5532 19287 7630
rect 19155 1932 19167 3238
rect 19203 1932 19215 3622
rect 19299 2412 19311 7630
rect 19323 7044 19335 7630
rect 19371 5220 19383 7630
rect 19395 6228 19407 7630
rect 19335 3252 19347 3958
rect 19419 2268 19431 7630
rect 19443 4332 19455 7630
rect 19491 7092 19503 7630
rect 19515 5532 19527 7630
rect 19563 5196 19575 7630
rect 19611 2076 19623 7630
rect 19635 4500 19647 7630
rect 19659 4260 19671 7630
rect 19707 6852 19719 7630
rect 19731 6060 19743 7630
rect 19779 6876 19791 7630
rect 19827 6468 19839 7630
rect 19851 3492 19863 7630
rect 19899 5964 19911 7630
rect 19947 6972 19959 7630
rect 19923 1932 19935 6022
rect 19995 5316 20007 7630
rect 20067 5412 20079 7630
rect 19995 1932 20007 3790
rect 20019 1932 20031 4150
rect 20043 1932 20055 4726
rect 20091 2220 20103 7630
rect 20139 5604 20151 7630
rect 20187 5052 20199 7630
rect 20211 2724 20223 7630
rect 20235 5820 20247 7630
rect 20259 5316 20271 7630
rect 20307 5772 20319 7630
rect 20211 1932 20223 2662
rect 20235 1932 20247 3934
rect 20283 1932 20295 5350
rect 20331 2676 20343 6406
rect 20355 5412 20367 7630
rect 20355 1932 20367 2782
rect 20379 1932 20391 6718
rect 20427 5196 20439 7630
rect 20451 5604 20463 7630
rect 20475 5628 20487 7630
rect 20403 1932 20415 4582
rect 20451 1932 20463 4894
rect 20475 1932 20487 4678
rect 20499 2196 20511 5398
rect 20523 5148 20535 7630
rect 20547 6756 20559 7630
rect 20547 1932 20559 4342
rect 20571 1932 20583 4774
rect 20595 4428 20607 7630
rect 20643 6108 20655 7630
rect 20667 6180 20679 7630
rect 20619 3300 20631 5590
rect 20595 1932 20607 2998
rect 20643 1932 20655 5902
rect 20691 5772 20703 7630
rect 20691 1932 20703 5686
rect 20715 2436 20727 5614
rect 20739 2892 20751 7630
rect 20763 5484 20775 7630
rect 20787 6420 20799 7630
rect 20763 1932 20775 3478
rect 20787 1932 20799 6310
rect 20811 1932 20823 5518
rect 20835 2604 20847 7630
rect 20859 7260 20871 7630
rect 20883 5292 20895 7630
rect 20907 4668 20919 7630
rect 20883 1932 20895 4486
rect 20907 1932 20919 4342
rect 20931 2292 20943 7630
rect 20955 5004 20967 6406
rect 20979 5268 20991 7630
rect 21027 5004 21039 7630
rect 21099 6996 21111 7630
rect 21123 6324 21135 7630
rect 21147 7020 21159 7630
rect 21051 4500 21063 5446
rect 21159 4356 21171 5422
rect 21195 3780 21207 7630
rect 21219 5148 21231 7630
rect 21243 5412 21255 7630
rect 21267 7380 21279 7630
rect 21315 7284 21327 7630
rect 21339 4692 21351 7630
rect 20931 1932 20943 2254
rect 20979 1932 20991 3742
rect 21003 1932 21015 2470
rect 21075 1932 21087 3190
rect 21195 1932 21207 3718
rect 21219 1932 21231 2590
rect 21291 1932 21303 3382
rect 21339 1932 21351 4486
rect 21363 2268 21375 7582
rect 21387 7188 21399 7630
rect 21435 6492 21447 7630
rect 21387 1932 21399 4678
rect 21411 3732 21423 5158
rect 21435 1932 21447 5782
rect 21459 5340 21471 7630
rect 21483 1932 21495 3358
rect 21507 2820 21519 7630
rect 21555 5100 21567 7630
rect 21507 1932 21519 2782
rect 21531 1932 21543 2926
rect 21555 1932 21567 4342
rect 21579 3876 21591 7630
rect 21603 4500 21615 6190
rect 21627 6108 21639 7630
rect 21579 1932 21591 3814
rect 21627 1932 21639 5878
rect 21675 4476 21687 7630
rect 21699 3876 21711 7630
rect 21723 5748 21735 7630
rect 21747 5340 21759 7630
rect 21651 1932 21663 3478
rect 21699 1932 21711 3766
rect 21759 2796 21771 4846
rect 21795 4308 21807 7630
rect 21819 4860 21831 7630
rect 21843 6252 21855 7630
rect 21795 1932 21807 2374
rect 21819 1932 21831 3598
rect 21843 1932 21855 3982
rect 21867 3828 21879 5854
rect 21891 3852 21903 7630
rect 21915 5844 21927 7630
rect 21939 6396 21951 7630
rect 21987 4956 21999 7630
rect 22035 5436 22047 7630
rect 21891 1932 21903 3718
rect 21951 2604 21963 4846
rect 22011 1932 22023 4630
rect 22035 1932 22047 5038
rect 22059 3780 22071 7246
rect 22107 4836 22119 7630
rect 22131 3732 22143 5662
rect 22155 5556 22167 7630
rect 22299 7356 22311 7630
rect 22083 1932 22095 2686
rect 22179 1932 22191 5494
rect 22251 1932 22263 7030
rect 22347 1932 22359 4630
rect 22395 1932 22407 3910
rect 22443 1932 22455 6238
rect 22467 1932 22479 4486
rect 22491 1932 22503 4870
rect 22515 1932 22527 4462
rect 22563 1932 22575 6982
rect 22587 1932 22599 2878
rect 22611 1932 22623 5998
rect 22659 5724 22671 7630
rect 22707 6324 22719 7630
rect 22659 1932 22671 5182
rect 22683 1932 22695 4894
rect 22755 1932 22767 2518
rect 22827 1932 22839 6814
rect 22851 4476 22863 7630
rect 22851 1932 22863 4318
rect 22899 3708 22911 7630
rect 22923 1932 22935 4894
rect 22947 3396 22959 7630
rect 22971 3372 22983 4918
rect 22947 1932 22959 3358
rect 22995 1932 23007 2614
rect 23019 1980 23031 7630
rect 23043 3468 23055 7630
rect 23067 3324 23079 7630
rect 23115 4860 23127 7630
rect 23139 4884 23151 7630
rect 23163 4428 23175 7630
rect 23115 1932 23127 2518
rect 23139 1932 23151 3142
rect 23187 1932 23199 6814
rect 23211 1932 23223 4462
rect 23235 4140 23247 7630
rect 23259 4908 23271 7630
rect 23259 1932 23271 3190
rect 23283 1932 23295 6454
rect 23307 5172 23319 7630
rect 23355 5124 23367 7630
rect 23379 5388 23391 7630
rect 23403 5172 23415 7630
rect 23307 1932 23319 4414
rect 23331 2364 23343 4870
rect 23355 1932 23367 4294
rect 23403 1932 23415 5110
rect 23427 4428 23439 7486
rect 23451 2916 23463 7630
rect 23475 5652 23487 7630
rect 23475 1932 23487 5278
rect 23499 4308 23511 6142
rect 23523 4068 23535 7630
rect 23547 4356 23559 5158
rect 23571 4140 23583 7630
rect 23595 4884 23607 7630
rect 23619 4764 23631 7630
rect 23667 6852 23679 7630
rect 23715 7452 23727 7630
rect 23571 1932 23583 3742
rect 23595 1932 23607 3694
rect 23643 2748 23655 4870
rect 23667 1932 23679 4750
rect 23739 1932 23751 6502
rect 23787 6492 23799 7630
rect 23787 1932 23799 6430
rect 23811 5316 23823 7630
rect 23835 4500 23847 6478
rect 23859 1932 23871 6334
rect 23883 4788 23895 7630
rect 23907 5100 23919 7630
rect 23931 4812 23943 7630
rect 23931 1932 23943 4414
rect 23955 4212 23967 7630
rect 24003 5748 24015 7630
rect 24027 4884 24039 7630
rect 24051 4908 24063 7630
rect 24027 1932 24039 4678
rect 24063 3492 24075 4870
rect 24099 4596 24111 7630
rect 24123 4692 24135 7630
rect 24147 4764 24159 7630
rect 24195 7212 24207 7630
rect 24219 7428 24231 7630
rect 24195 1932 24207 5902
rect 24219 1932 24231 2590
rect 24243 2316 24255 7630
rect 24267 2292 24279 7534
rect 24291 4980 24303 7630
rect 24243 1932 24255 2278
rect 24291 1932 24303 4750
rect 24315 4020 24327 7630
rect 24339 5148 24351 7630
rect 24363 4764 24375 7510
rect 24315 1932 24327 3262
rect 24387 3108 24399 7630
rect 24411 5340 24423 7630
rect 24411 1932 24423 4894
rect 24435 4740 24447 7630
rect 24459 4692 24471 7630
rect 24483 5124 24495 7630
rect 24435 1932 24447 3502
rect 24483 1932 24495 5086
rect 24507 1932 24519 5350
rect 24531 5292 24543 7630
rect 24555 5676 24567 7630
rect 24531 1932 24543 5206
rect 24603 4884 24615 7630
rect 24651 6924 24663 7630
rect 24675 5988 24687 7630
rect 24579 1932 24591 2686
rect 24603 1932 24615 4678
rect 24627 3228 24639 5110
rect 24675 1932 24687 4750
rect 24699 1932 24711 5494
rect 24723 5292 24735 7630
rect 24735 3204 24747 4870
rect 24771 3540 24783 7630
rect 24819 4452 24831 7630
rect 24891 5100 24903 7630
rect 24771 1932 24783 3502
rect 24795 1932 24807 2086
rect 24819 1932 24831 3646
rect 24867 1932 24879 4510
rect 24891 1932 24903 4726
rect 24915 4524 24927 7630
rect 24939 5268 24951 7630
rect 24987 7092 24999 7630
rect 24951 4740 24963 5182
rect 24939 1932 24951 2038
rect 24987 1932 24999 6862
rect 25011 5532 25023 7630
rect 25011 1932 25023 3382
rect 25035 1932 25047 4846
rect 25083 1932 25095 4990
rect 25107 4860 25119 7630
rect 25179 6276 25191 7630
rect 25203 6828 25215 7630
rect 25107 1932 25119 4798
rect 25131 1932 25143 5398
rect 25227 5388 25239 7630
rect 25155 3036 25167 4846
rect 25179 1932 25191 3742
rect 25203 1932 25215 3550
rect 25227 1932 25239 5350
rect 25251 4116 25263 5374
rect 25275 3564 25287 7630
rect 25299 3876 25311 7630
rect 25347 4380 25359 7630
rect 25395 4140 25407 7630
rect 25419 4620 25431 7630
rect 25443 6612 25455 7630
rect 25491 7140 25503 7630
rect 25515 5940 25527 7630
rect 25563 7500 25575 7630
rect 25275 1932 25287 2470
rect 25299 1932 25311 3190
rect 25323 1932 25335 3262
rect 25347 1932 25359 2854
rect 25395 1932 25407 4102
rect 25467 1932 25479 4726
rect 25515 1932 25527 3790
rect 25539 1932 25551 3454
rect 25563 1932 25575 7462
rect 25587 4116 25599 5230
rect 25611 2604 25623 7630
rect 25635 4692 25647 7630
rect 25683 7068 25695 7630
rect 25635 1932 25647 3094
rect 25659 1932 25671 3550
rect 25707 1932 25719 5062
rect 25731 4716 25743 7630
rect 25755 5772 25767 7630
rect 25779 4236 25791 7486
rect 25827 5700 25839 7630
rect 25851 5436 25863 7630
rect 25875 5292 25887 7630
rect 25899 5748 25911 7630
rect 25923 6636 25935 7630
rect 25827 1932 25839 3742
rect 25971 3444 25983 7630
rect 26019 6564 26031 7630
rect 26091 4428 26103 7630
rect 26115 2100 26127 7630
rect 26139 2556 26151 7630
rect 26187 2124 26199 7630
rect 26211 3084 26223 7630
rect 26235 4740 26247 7630
rect 26259 4284 26271 7630
rect 26283 2340 26295 7630
rect 26331 3180 26343 7630
rect 26355 4188 26367 7630
rect 26379 4764 26391 7630
rect 26331 1932 26343 3142
rect 26379 1932 26391 3742
rect 26403 3156 26415 5830
rect 26427 4092 26439 7630
rect 26499 6348 26511 7630
rect 26547 1932 26559 3790
rect 26571 3516 26583 7630
rect 26643 5364 26655 7630
rect 26667 3804 26679 7630
rect 26691 4836 26703 7630
rect 26739 5292 26751 7630
rect 26763 4692 26775 7630
rect 26787 4620 26799 5878
rect 26643 1932 26655 3118
rect 26763 1932 26775 4606
rect 26811 4140 26823 7630
rect 26859 7140 26871 7630
rect 26883 3564 26895 7630
rect 26907 5604 26919 7630
rect 26907 1932 26919 5566
rect 26931 4548 26943 5590
rect 26955 4668 26967 7630
rect 27003 6468 27015 7630
rect 27075 6540 27087 7630
rect 27099 2148 27111 7630
rect 27123 4644 27135 7630
rect 27171 3708 27183 7630
rect 27195 5292 27207 7630
rect 27219 6468 27231 7630
rect 27243 5028 27255 7630
rect 27291 7092 27303 7630
rect 27315 6036 27327 7630
rect 27339 5892 27351 7630
rect 27363 4500 27375 7630
rect 27411 3804 27423 7630
rect 27435 6204 27447 7630
rect 27459 6900 27471 7630
rect 27267 1932 27279 1942
rect 27315 1932 27327 3094
rect 27507 2724 27519 7630
rect 27531 3804 27543 7630
rect 27555 4404 27567 7630
rect 27603 4788 27615 7630
rect 27627 3876 27639 7630
rect 27675 2244 27687 7630
rect 27723 4476 27735 7630
rect 27771 4332 27783 7630
rect 27771 1956 27783 3478
rect 27795 1980 27807 4678
rect 27819 2004 27831 4558
rect 27843 2028 27855 3502
rect 27867 2052 27879 6358
rect 27891 2076 27903 4414
rect 27915 1932 28115 7630
rect 28241 2495 28311 2507
rect 28241 2063 28311 2075
rect 28241 2039 28311 2051
rect 28241 2015 28311 2027
rect 28241 1991 28311 2003
rect 28241 1967 28311 1979
rect 28241 1943 28311 1955
rect 0 78 70 90
rect 0 54 70 66
rect 0 30 70 42
rect 0 6 70 18
rect 123 0 323 1133
rect 339 0 351 1133
rect 363 0 375 1133
rect 387 0 399 1133
rect 411 0 423 1133
rect 1635 115 1647 1133
rect 1707 139 1719 1133
rect 1755 67 1767 1133
rect 2643 67 2655 1133
rect 2667 163 2679 1133
rect 2691 187 2703 1133
rect 2811 211 2823 1133
rect 3363 235 3375 1133
rect 3507 259 3519 1133
rect 3747 283 3759 1133
rect 3819 307 3831 1133
rect 4035 331 4047 1133
rect 4059 355 4071 1133
rect 4323 379 4335 1133
rect 4395 403 4407 1133
rect 4587 427 4599 1133
rect 4659 451 4671 1133
rect 4731 475 4743 1133
rect 4803 499 4815 1133
rect 4923 523 4935 1133
rect 4947 547 4959 1133
rect 5787 571 5799 1133
rect 5883 595 5895 1133
rect 5955 619 5967 1133
rect 6267 643 6279 1133
rect 6339 667 6351 1133
rect 6507 691 6519 1133
rect 6555 523 6567 1133
rect 6723 715 6735 1133
rect 6747 739 6759 1133
rect 6819 763 6831 1133
rect 6867 787 6879 1133
rect 6939 787 6951 1133
rect 7179 499 7191 1133
rect 7203 787 7215 1133
rect 7299 811 7311 1133
rect 7323 739 7335 1133
rect 7659 595 7671 1133
rect 8067 595 8079 1133
rect 8091 835 8103 1133
rect 8307 859 8319 1133
rect 8427 883 8439 1133
rect 9123 907 9135 1133
rect 9339 931 9351 1133
rect 9675 955 9687 1133
rect 9747 811 9759 1133
rect 10059 811 10071 1133
rect 10371 979 10383 1133
rect 10419 1003 10431 1133
rect 10443 283 10455 1133
rect 10611 283 10623 1133
rect 10779 667 10791 1133
rect 10827 499 10839 1133
rect 10995 643 11007 1133
rect 11043 643 11055 1133
rect 11067 811 11079 1133
rect 11091 451 11103 1133
rect 11427 355 11439 1133
rect 11475 811 11487 1133
rect 11523 499 11535 1133
rect 11667 1003 11679 1133
rect 11715 1003 11727 1133
rect 11859 451 11871 1133
rect 11883 355 11895 1133
rect 12147 595 12159 1133
rect 12411 907 12423 1133
rect 12579 43 12591 1133
rect 12627 43 12639 1133
rect 12819 931 12831 1133
rect 12843 667 12855 1133
rect 13347 715 13359 1133
rect 13443 715 13455 1133
rect 13635 187 13647 1133
rect 13659 883 13671 1133
rect 13779 883 13791 1133
rect 13947 355 13959 1133
rect 14067 355 14079 1133
rect 14355 811 14367 1133
rect 14931 811 14943 1133
rect 15051 187 15063 1133
rect 15795 1027 15807 1133
rect 15891 1051 15903 1133
rect 15987 1075 15999 1133
rect 16203 1099 16215 1133
rect 16251 1123 16263 1133
rect 16275 1051 16287 1133
rect 16443 19 16455 1133
rect 16563 763 16575 1133
rect 16683 67 16695 1133
rect 17043 163 17055 1133
rect 17235 1051 17247 1133
rect 17259 979 17271 1133
rect 17283 163 17295 1133
rect 17475 979 17487 1133
rect 17571 907 17583 1133
rect 17595 715 17607 1133
rect 17667 715 17679 1133
rect 17859 1003 17871 1133
rect 17907 691 17919 1133
rect 18027 691 18039 1133
rect 18051 931 18063 1133
rect 18483 331 18495 1133
rect 18603 883 18615 1133
rect 18627 907 18639 1133
rect 18651 787 18663 1133
rect 18867 1099 18879 1133
rect 18915 211 18927 1133
rect 19011 1051 19023 1133
rect 19059 787 19071 1133
rect 19107 523 19119 1133
rect 19347 427 19359 1133
rect 19755 67 19767 1133
rect 19899 139 19911 1133
rect 19947 43 19959 1133
rect 20091 499 20103 1133
rect 20139 451 20151 1133
rect 20259 859 20271 1133
rect 20307 859 20319 1133
rect 20499 499 20511 1133
rect 20811 235 20823 1133
rect 20835 115 20847 1133
rect 21027 259 21039 1133
rect 21099 811 21111 1133
rect 21123 163 21135 1133
rect 21171 763 21183 1133
rect 21243 715 21255 1133
rect 21315 931 21327 1133
rect 21411 331 21423 1133
rect 21747 715 21759 1133
rect 21771 283 21783 1133
rect 21891 307 21903 1133
rect 21915 691 21927 1133
rect 21939 931 21951 1133
rect 21963 1123 21975 1133
rect 22131 667 22143 1133
rect 22275 91 22287 1133
rect 22299 979 22311 1133
rect 22371 1075 22383 1133
rect 22707 787 22719 1133
rect 22779 619 22791 1133
rect 22803 1027 22815 1133
rect 22899 571 22911 1133
rect 23043 355 23055 1133
rect 23163 475 23175 1133
rect 23499 667 23511 1133
rect 23523 715 23535 1133
rect 23619 739 23631 1133
rect 23691 547 23703 1133
rect 24003 667 24015 1133
rect 24123 691 24135 1133
rect 24339 907 24351 1133
rect 24387 763 24399 1133
rect 24627 619 24639 1133
rect 24723 643 24735 1133
rect 25419 403 25431 1133
rect 25731 955 25743 1133
rect 25803 835 25815 1133
rect 25851 379 25863 1133
rect 25971 859 25983 1133
rect 26571 931 26583 1133
rect 26619 187 26631 1133
rect 26715 235 26727 1133
rect 26727 139 26739 221
rect 26763 19 26775 653
rect 26787 43 26799 293
rect 26811 67 26823 917
rect 26835 91 26847 581
rect 26859 115 26871 317
rect 27915 0 28115 1133
rect 28241 126 28311 138
rect 28241 102 28311 114
rect 28241 78 28311 90
rect 28241 54 28311 66
rect 28241 30 28311 42
rect 28241 6 28311 18
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 7630
box 0 0 1464 799
use nand2 g7994
timestamp 1386234792
transform 1 0 1587 0 1 7630
box 0 0 96 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 1683 0 1 7630
box 0 0 48 799
use rowcrosser AluEn
timestamp 1386086759
transform 1 0 1731 0 1 7630
box 0 0 48 799
use nand2 g8032
timestamp 1386234792
transform 1 0 1779 0 1 7630
box 0 0 96 799
use nand2 g7941
timestamp 1386234792
transform 1 0 1875 0 1 7630
box 0 0 96 799
use nand4 g8197
timestamp 1386234936
transform 1 0 1971 0 1 7630
box 0 0 144 799
use nand2 g8043
timestamp 1386234792
transform 1 0 2115 0 1 7630
box 0 0 96 799
use nand3 g8112
timestamp 1386234893
transform 1 0 2211 0 1 7630
box 0 0 120 799
use and2 g8291
timestamp 1386234845
transform 1 0 2331 0 1 7630
box 0 0 120 799
use nand2 g7923
timestamp 1386234792
transform 1 0 2451 0 1 7630
box 0 0 96 799
use nand3 g8060
timestamp 1386234893
transform 1 0 2547 0 1 7630
box 0 0 120 799
use nand2 g7942
timestamp 1386234792
transform 1 0 2667 0 1 7630
box 0 0 96 799
use nand3 g8182
timestamp 1386234893
transform 1 0 2763 0 1 7630
box 0 0 120 799
use nand2 g8066
timestamp 1386234792
transform 1 0 2883 0 1 7630
box 0 0 96 799
use nand2 g8169
timestamp 1386234792
transform 1 0 2979 0 1 7630
box 0 0 96 799
use nand2 g7934
timestamp 1386234792
transform 1 0 3075 0 1 7630
box 0 0 96 799
use inv g8107
timestamp 1386238110
transform 1 0 3171 0 1 7630
box 0 0 120 799
use and2 g8229
timestamp 1386234845
transform 1 0 3291 0 1 7630
box 0 0 120 799
use nand2 g8039
timestamp 1386234792
transform 1 0 3411 0 1 7630
box 0 0 96 799
use nand2 g8046
timestamp 1386234792
transform 1 0 3507 0 1 7630
box 0 0 96 799
use nand2 g8123
timestamp 1386234792
transform 1 0 3603 0 1 7630
box 0 0 96 799
use nand2 g8222
timestamp 1386234792
transform 1 0 3699 0 1 7630
box 0 0 96 799
use nand2 g8098
timestamp 1386234792
transform 1 0 3795 0 1 7630
box 0 0 96 799
use nand3 g8102
timestamp 1386234893
transform 1 0 3891 0 1 7630
box 0 0 120 799
use inv g8012
timestamp 1386238110
transform 1 0 4011 0 1 7630
box 0 0 120 799
use nand2 g8187
timestamp 1386234792
transform 1 0 4131 0 1 7630
box 0 0 96 799
use nand2 g7951
timestamp 1386234792
transform 1 0 4227 0 1 7630
box 0 0 96 799
use nand4 g8135
timestamp 1386234936
transform 1 0 4323 0 1 7630
box 0 0 144 799
use nand4 g8171
timestamp 1386234936
transform 1 0 4467 0 1 7630
box 0 0 144 799
use nand3 g8295
timestamp 1386234893
transform 1 0 4611 0 1 7630
box 0 0 120 799
use inv g8287
timestamp 1386238110
transform 1 0 4731 0 1 7630
box 0 0 120 799
use inv g8154
timestamp 1386238110
transform 1 0 4851 0 1 7630
box 0 0 120 799
use nand2 g8261
timestamp 1386234792
transform 1 0 4971 0 1 7630
box 0 0 96 799
use nand2 g8276
timestamp 1386234792
transform 1 0 5067 0 1 7630
box 0 0 96 799
use nand2 g8130
timestamp 1386234792
transform 1 0 5163 0 1 7630
box 0 0 96 799
use nand4 g8027
timestamp 1386234936
transform 1 0 5259 0 1 7630
box 0 0 144 799
use nand2 g8082
timestamp 1386234792
transform 1 0 5403 0 1 7630
box 0 0 96 799
use inv g8035
timestamp 1386238110
transform 1 0 5499 0 1 7630
box 0 0 120 799
use nand3 g8019
timestamp 1386234893
transform 1 0 5619 0 1 7630
box 0 0 120 799
use nand2 g8238
timestamp 1386234792
transform 1 0 5739 0 1 7630
box 0 0 96 799
use inv g8168
timestamp 1386238110
transform 1 0 5835 0 1 7630
box 0 0 120 799
use nand2 g7989
timestamp 1386234792
transform 1 0 5955 0 1 7630
box 0 0 96 799
use nand2 g8225
timestamp 1386234792
transform 1 0 6051 0 1 7630
box 0 0 96 799
use and2 g8143
timestamp 1386234845
transform 1 0 6147 0 1 7630
box 0 0 120 799
use nand2 g454
timestamp 1386234792
transform 1 0 6267 0 1 7630
box 0 0 96 799
use trisbuf g8042
timestamp 1386237216
transform 1 0 6363 0 1 7630
box 0 0 216 799
use nand3 g8069
timestamp 1386234893
transform 1 0 6579 0 1 7630
box 0 0 120 799
use nand2 g8149
timestamp 1386234792
transform 1 0 6699 0 1 7630
box 0 0 96 799
use and2 g7926
timestamp 1386234845
transform 1 0 6795 0 1 7630
box 0 0 120 799
use rowcrosser PcSel_91_1_93_
timestamp 1386086759
transform 1 0 6915 0 1 7630
box 0 0 48 799
use nand4 g8280
timestamp 1386234936
transform 1 0 6963 0 1 7630
box 0 0 144 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 7107 0 1 7630
box 0 0 48 799
use inv g7985
timestamp 1386238110
transform 1 0 7155 0 1 7630
box 0 0 120 799
use nand4 g8249
timestamp 1386234936
transform 1 0 7275 0 1 7630
box 0 0 144 799
use inv g8064
timestamp 1386238110
transform 1 0 7419 0 1 7630
box 0 0 120 799
use nand2 g8235
timestamp 1386234792
transform 1 0 7539 0 1 7630
box 0 0 96 799
use nand2 g7948
timestamp 1386234792
transform 1 0 7635 0 1 7630
box 0 0 96 799
use nand3 g8058
timestamp 1386234893
transform 1 0 7731 0 1 7630
box 0 0 120 799
use nor2 g8009
timestamp 1386235306
transform 1 0 7851 0 1 7630
box 0 0 120 799
use nand2 g7939
timestamp 1386234792
transform 1 0 7971 0 1 7630
box 0 0 96 799
use nand4 g8088
timestamp 1386234936
transform 1 0 8067 0 1 7630
box 0 0 144 799
use nand2 g8055
timestamp 1386234792
transform 1 0 8211 0 1 7630
box 0 0 96 799
use nand2 g7947
timestamp 1386234792
transform 1 0 8307 0 1 7630
box 0 0 96 799
use nand2 g7960
timestamp 1386234792
transform 1 0 8403 0 1 7630
box 0 0 96 799
use nand2 g8214
timestamp 1386234792
transform 1 0 8499 0 1 7630
box 0 0 96 799
use nand3 g8056
timestamp 1386234893
transform 1 0 8595 0 1 7630
box 0 0 120 799
use rowcrosser AluOR_91_0_93_
timestamp 1386086759
transform 1 0 8715 0 1 7630
box 0 0 48 799
use nand2 g8281
timestamp 1386234792
transform 1 0 8763 0 1 7630
box 0 0 96 799
use nand2 g8269
timestamp 1386234792
transform 1 0 8859 0 1 7630
box 0 0 96 799
use and2 g8183
timestamp 1386234845
transform 1 0 8955 0 1 7630
box 0 0 120 799
use nand3 g8170
timestamp 1386234893
transform 1 0 9075 0 1 7630
box 0 0 120 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 9195 0 1 7630
box 0 0 48 799
use nand2 g8124
timestamp 1386234792
transform 1 0 9243 0 1 7630
box 0 0 96 799
use nand4 g8106
timestamp 1386234936
transform 1 0 9339 0 1 7630
box 0 0 144 799
use nand2 g8119
timestamp 1386234792
transform 1 0 9483 0 1 7630
box 0 0 96 799
use nand2 g8275
timestamp 1386234792
transform 1 0 9579 0 1 7630
box 0 0 96 799
use inv g8146
timestamp 1386238110
transform 1 0 9675 0 1 7630
box 0 0 120 799
use nand2 g8127
timestamp 1386234792
transform 1 0 9795 0 1 7630
box 0 0 96 799
use nand2 g8155
timestamp 1386234792
transform 1 0 9891 0 1 7630
box 0 0 96 799
use nand3 g8290
timestamp 1386234893
transform 1 0 9987 0 1 7630
box 0 0 120 799
use inv g7909
timestamp 1386238110
transform 1 0 10107 0 1 7630
box 0 0 120 799
use nand4 g8033
timestamp 1386234936
transform 1 0 10227 0 1 7630
box 0 0 144 799
use nand2 g7921
timestamp 1386234792
transform 1 0 10371 0 1 7630
box 0 0 96 799
use nand3 g8252
timestamp 1386234893
transform 1 0 10467 0 1 7630
box 0 0 120 799
use nand2 g7978
timestamp 1386234792
transform 1 0 10587 0 1 7630
box 0 0 96 799
use inv g8244
timestamp 1386238110
transform 1 0 10683 0 1 7630
box 0 0 120 799
use nand2 g7930
timestamp 1386234792
transform 1 0 10803 0 1 7630
box 0 0 96 799
use nand2 g7972
timestamp 1386234792
transform 1 0 10899 0 1 7630
box 0 0 96 799
use nand3 g8240
timestamp 1386234893
transform 1 0 10995 0 1 7630
box 0 0 120 799
use nand2 g8054
timestamp 1386234792
transform 1 0 11115 0 1 7630
box 0 0 96 799
use nand2 g8139
timestamp 1386234792
transform 1 0 11211 0 1 7630
box 0 0 96 799
use nand3 g8023
timestamp 1386234893
transform 1 0 11307 0 1 7630
box 0 0 120 799
use nand2 g8118
timestamp 1386234792
transform 1 0 11427 0 1 7630
box 0 0 96 799
use nand2 g7981
timestamp 1386234792
transform 1 0 11523 0 1 7630
box 0 0 96 799
use nand3 g8111
timestamp 1386234893
transform 1 0 11619 0 1 7630
box 0 0 120 799
use and2 g8120
timestamp 1386234845
transform 1 0 11739 0 1 7630
box 0 0 120 799
use nor2 g8091
timestamp 1386235306
transform 1 0 11859 0 1 7630
box 0 0 120 799
use nand4 g7918
timestamp 1386234936
transform 1 0 11979 0 1 7630
box 0 0 144 799
use nand4 g8134
timestamp 1386234936
transform 1 0 12123 0 1 7630
box 0 0 144 799
use nand2 g8050
timestamp 1386234792
transform 1 0 12267 0 1 7630
box 0 0 96 799
use nand3 g8218
timestamp 1386234893
transform 1 0 12363 0 1 7630
box 0 0 120 799
use and2 g7995
timestamp 1386234845
transform 1 0 12483 0 1 7630
box 0 0 120 799
use nand2 g7945
timestamp 1386234792
transform 1 0 12603 0 1 7630
box 0 0 96 799
use nand2 g8284
timestamp 1386234792
transform 1 0 12699 0 1 7630
box 0 0 96 799
use nand2 g7964
timestamp 1386234792
transform 1 0 12795 0 1 7630
box 0 0 96 799
use inv g8198
timestamp 1386238110
transform 1 0 12891 0 1 7630
box 0 0 120 799
use rowcrosser g8048
timestamp 1386086759
transform 1 0 13011 0 1 7630
box 0 0 48 799
use nand2 g8272
timestamp 1386234792
transform 1 0 13059 0 1 7630
box 0 0 96 799
use nand2 g8199
timestamp 1386234792
transform 1 0 13155 0 1 7630
box 0 0 96 799
use nand2 g8221
timestamp 1386234792
transform 1 0 13251 0 1 7630
box 0 0 96 799
use rowcrosser Op1Sel
timestamp 1386086759
transform 1 0 13347 0 1 7630
box 0 0 48 799
use nand2 g8220
timestamp 1386234792
transform 1 0 13395 0 1 7630
box 0 0 96 799
use nand2 g8230
timestamp 1386234792
transform 1 0 13491 0 1 7630
box 0 0 96 799
use nand2 g8271
timestamp 1386234792
transform 1 0 13587 0 1 7630
box 0 0 96 799
use inv g8004
timestamp 1386238110
transform 1 0 13683 0 1 7630
box 0 0 120 799
use and2 g8074
timestamp 1386234845
transform 1 0 13803 0 1 7630
box 0 0 120 799
use and2 g8209
timestamp 1386234845
transform 1 0 13923 0 1 7630
box 0 0 120 799
use and2 g8103
timestamp 1386234845
transform 1 0 14043 0 1 7630
box 0 0 120 799
use nor2 g8283
timestamp 1386235306
transform 1 0 14163 0 1 7630
box 0 0 120 799
use nor2 g8268
timestamp 1386235306
transform 1 0 14283 0 1 7630
box 0 0 120 799
use and2 g8180
timestamp 1386234845
transform 1 0 14403 0 1 7630
box 0 0 120 799
use nand2 g8005
timestamp 1386234792
transform 1 0 14523 0 1 7630
box 0 0 96 799
use and2 g8052
timestamp 1386234845
transform 1 0 14619 0 1 7630
box 0 0 120 799
use nand4 g8136
timestamp 1386234936
transform 1 0 14739 0 1 7630
box 0 0 144 799
use nand2 g8110
timestamp 1386234792
transform 1 0 14883 0 1 7630
box 0 0 96 799
use nand3 g8153
timestamp 1386234893
transform 1 0 14979 0 1 7630
box 0 0 120 799
use nor2 StatusReg_reg_91_3_93_
timestamp 1386235306
transform 1 0 15099 0 1 7630
box 0 0 120 799
use scandtype g7922
timestamp 1386241841
transform 1 0 15219 0 1 7630
box 0 0 624 799
use nand3 g8308
timestamp 1386234893
transform 1 0 15843 0 1 7630
box 0 0 120 799
use inv stateSub_reg_91_2_93_
timestamp 1386238110
transform 1 0 15963 0 1 7630
box 0 0 120 799
use scandtype g7943
timestamp 1386241841
transform 1 0 16083 0 1 7630
box 0 0 624 799
use nand2 g8024
timestamp 1386234792
transform 1 0 16707 0 1 7630
box 0 0 96 799
use rowcrosser RwSel_91_1_93_
timestamp 1386086759
transform 1 0 16803 0 1 7630
box 0 0 48 799
use inv g8099
timestamp 1386238110
transform 1 0 16851 0 1 7630
box 0 0 120 799
use nand3 g8057
timestamp 1386234893
transform 1 0 16971 0 1 7630
box 0 0 120 799
use nand3 g8190
timestamp 1386234893
transform 1 0 17091 0 1 7630
box 0 0 120 799
use nand3 g8045
timestamp 1386234893
transform 1 0 17211 0 1 7630
box 0 0 120 799
use nand2 g8304
timestamp 1386234792
transform 1 0 17331 0 1 7630
box 0 0 96 799
use inv g8018
timestamp 1386238110
transform 1 0 17427 0 1 7630
box 0 0 120 799
use nand2 g8092
timestamp 1386234792
transform 1 0 17547 0 1 7630
box 0 0 96 799
use nand2 g8277
timestamp 1386234792
transform 1 0 17643 0 1 7630
box 0 0 96 799
use nor2 g8081
timestamp 1386235306
transform 1 0 17739 0 1 7630
box 0 0 120 799
use nand2 g8243
timestamp 1386234792
transform 1 0 17859 0 1 7630
box 0 0 96 799
use nand2 g8234
timestamp 1386234792
transform 1 0 17955 0 1 7630
box 0 0 96 799
use and2 StatusReg_reg_91_1_93_
timestamp 1386234845
transform 1 0 18051 0 1 7630
box 0 0 120 799
use scandtype g7933
timestamp 1386241841
transform 1 0 18171 0 1 7630
box 0 0 624 799
use rowcrosser RegWe
timestamp 1386086759
transform 1 0 18795 0 1 7630
box 0 0 48 799
use rowcrosser nWait
timestamp 1386086759
transform 1 0 18843 0 1 7630
box 0 0 48 799
use nand3 g8028
timestamp 1386234893
transform 1 0 18891 0 1 7630
box 0 0 120 799
use nand2 g8213
timestamp 1386234792
transform 1 0 19011 0 1 7630
box 0 0 96 799
use nand2 g7963
timestamp 1386234792
transform 1 0 19107 0 1 7630
box 0 0 96 799
use nand4 g8096
timestamp 1386234936
transform 1 0 19203 0 1 7630
box 0 0 144 799
use nand3 g8212
timestamp 1386234893
transform 1 0 19347 0 1 7630
box 0 0 120 799
use and2 g8015
timestamp 1386234845
transform 1 0 19467 0 1 7630
box 0 0 120 799
use nand2 g8084
timestamp 1386234792
transform 1 0 19587 0 1 7630
box 0 0 96 799
use nor2 g8265
timestamp 1386235306
transform 1 0 19683 0 1 7630
box 0 0 120 799
use nor2 g8200
timestamp 1386235306
transform 1 0 19803 0 1 7630
box 0 0 120 799
use inv g8108
timestamp 1386238110
transform 1 0 19923 0 1 7630
box 0 0 120 799
use nor2 g8049
timestamp 1386235306
transform 1 0 20043 0 1 7630
box 0 0 120 799
use nand3 g8159
timestamp 1386234893
transform 1 0 20163 0 1 7630
box 0 0 120 799
use inv g8144
timestamp 1386238110
transform 1 0 20283 0 1 7630
box 0 0 120 799
use nand2 g8177
timestamp 1386234792
transform 1 0 20403 0 1 7630
box 0 0 96 799
use and2 g7996
timestamp 1386234845
transform 1 0 20499 0 1 7630
box 0 0 120 799
use nand2 g8251
timestamp 1386234792
transform 1 0 20619 0 1 7630
box 0 0 96 799
use nand2 g8036
timestamp 1386234792
transform 1 0 20715 0 1 7630
box 0 0 96 799
use nand4 g8226
timestamp 1386234936
transform 1 0 20811 0 1 7630
box 0 0 144 799
use inv g7929
timestamp 1386238110
transform 1 0 20955 0 1 7630
box 0 0 120 799
use nand2 g7979
timestamp 1386234792
transform 1 0 21075 0 1 7630
box 0 0 96 799
use nand3 g8264
timestamp 1386234893
transform 1 0 21171 0 1 7630
box 0 0 120 799
use nor2 g8089
timestamp 1386235306
transform 1 0 21291 0 1 7630
box 0 0 120 799
use and2 g8206
timestamp 1386234845
transform 1 0 21411 0 1 7630
box 0 0 120 799
use and2 g8237
timestamp 1386234845
transform 1 0 21531 0 1 7630
box 0 0 120 799
use nand3 g8016
timestamp 1386234893
transform 1 0 21651 0 1 7630
box 0 0 120 799
use nand2 g8278
timestamp 1386234792
transform 1 0 21771 0 1 7630
box 0 0 96 799
use nand2 g8181
timestamp 1386234792
transform 1 0 21867 0 1 7630
box 0 0 96 799
use inv g8216
timestamp 1386238110
transform 1 0 21963 0 1 7630
box 0 0 120 799
use inv StatusReg_reg_91_0_93_
timestamp 1386238110
transform 1 0 22083 0 1 7630
box 0 0 120 799
use scandtype g8253
timestamp 1386241841
transform 1 0 22203 0 1 7630
box 0 0 624 799
use rowcrosser Op2Sel_91_0_93_
timestamp 1386086759
transform 1 0 22827 0 1 7630
box 0 0 48 799
use inv g8186
timestamp 1386238110
transform 1 0 22875 0 1 7630
box 0 0 120 799
use nand2 g7946
timestamp 1386234792
transform 1 0 22995 0 1 7630
box 0 0 96 799
use nand3 g8090
timestamp 1386234893
transform 1 0 23091 0 1 7630
box 0 0 120 799
use and2 g8223
timestamp 1386234845
transform 1 0 23211 0 1 7630
box 0 0 120 799
use nand2 g8195
timestamp 1386234792
transform 1 0 23331 0 1 7630
box 0 0 96 799
use nor2 g8077
timestamp 1386235306
transform 1 0 23427 0 1 7630
box 0 0 120 799
use nand2 g8133
timestamp 1386234792
transform 1 0 23547 0 1 7630
box 0 0 96 799
use inv g7971
timestamp 1386238110
transform 1 0 23643 0 1 7630
box 0 0 120 799
use nand2 g8041
timestamp 1386234792
transform 1 0 23763 0 1 7630
box 0 0 96 799
use nand3 g8289
timestamp 1386234893
transform 1 0 23859 0 1 7630
box 0 0 120 799
use nand2 g8002
timestamp 1386234792
transform 1 0 23979 0 1 7630
box 0 0 96 799
use nand2 g8128
timestamp 1386234792
transform 1 0 24075 0 1 7630
box 0 0 96 799
use nand2 g8029
timestamp 1386234792
transform 1 0 24171 0 1 7630
box 0 0 96 799
use nand2 g8100
timestamp 1386234792
transform 1 0 24267 0 1 7630
box 0 0 96 799
use nand4 g8117
timestamp 1386234936
transform 1 0 24363 0 1 7630
box 0 0 144 799
use and2 g8167
timestamp 1386234845
transform 1 0 24507 0 1 7630
box 0 0 120 799
use and2 g7982
timestamp 1386234845
transform 1 0 24627 0 1 7630
box 0 0 120 799
use inv g8227
timestamp 1386238110
transform 1 0 24747 0 1 7630
box 0 0 120 799
use nand2 g8191
timestamp 1386234792
transform 1 0 24867 0 1 7630
box 0 0 96 799
use xor2 g7975
timestamp 1386237344
transform 1 0 24963 0 1 7630
box 0 0 192 799
use nand2 g8270
timestamp 1386234792
transform 1 0 25155 0 1 7630
box 0 0 96 799
use nor2 g8073
timestamp 1386235306
transform 1 0 25251 0 1 7630
box 0 0 120 799
use nand2 g8163
timestamp 1386234792
transform 1 0 25371 0 1 7630
box 0 0 96 799
use nor2 g8273
timestamp 1386235306
transform 1 0 25467 0 1 7630
box 0 0 120 799
use and2 g7969
timestamp 1386234845
transform 1 0 25587 0 1 7630
box 0 0 120 799
use nand2 g8051
timestamp 1386234792
transform 1 0 25707 0 1 7630
box 0 0 96 799
use nand4 g8147
timestamp 1386234936
transform 1 0 25803 0 1 7630
box 0 0 144 799
use inv g7955
timestamp 1386238110
transform 1 0 25947 0 1 7630
box 0 0 120 799
use nand2 g7928
timestamp 1386234792
transform 1 0 26067 0 1 7630
box 0 0 96 799
use nand4 g8030
timestamp 1386234936
transform 1 0 26163 0 1 7630
box 0 0 144 799
use nand2 g1
timestamp 1386234792
transform 1 0 26307 0 1 7630
box 0 0 96 799
use trisbuf g8217
timestamp 1386237216
transform 1 0 26403 0 1 7630
box 0 0 216 799
use nand2 g8114
timestamp 1386234792
transform 1 0 26619 0 1 7630
box 0 0 96 799
use and2 g8174
timestamp 1386234845
transform 1 0 26715 0 1 7630
box 0 0 120 799
use nand2 g8305
timestamp 1386234792
transform 1 0 26835 0 1 7630
box 0 0 96 799
use inv g8241
timestamp 1386238110
transform 1 0 26931 0 1 7630
box 0 0 120 799
use nand2 g8067
timestamp 1386234792
transform 1 0 27051 0 1 7630
box 0 0 96 799
use nand3 g7990
timestamp 1386234893
transform 1 0 27147 0 1 7630
box 0 0 120 799
use nand3 g8158
timestamp 1386234893
transform 1 0 27267 0 1 7630
box 0 0 120 799
use nand2 g8063
timestamp 1386234792
transform 1 0 27387 0 1 7630
box 0 0 96 799
use nand2 g8257
timestamp 1386234792
transform 1 0 27483 0 1 7630
box 0 0 96 799
use and2 RwSel_91_0_93_
timestamp 1386234845
transform 1 0 27579 0 1 7630
box 0 0 120 799
use rowcrosser nME
timestamp 1386086759
transform 1 0 27699 0 1 7630
box 0 0 48 799
use rowcrosser PcSel_91_0_93_
timestamp 1386086759
transform 1 0 27747 0 1 7630
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 27795 0 1 7630
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 1133
box 0 0 1464 799
use nand4 stateSub_reg_91_0_93_
timestamp 1386234936
transform 1 0 1587 0 1 1133
box 0 0 144 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 1731 0 1 1133
box 0 0 48 799
use scandtype g8020
timestamp 1386241841
transform 1 0 1779 0 1 1133
box 0 0 624 799
use nand2 g8150
timestamp 1386234792
transform 1 0 2403 0 1 1133
box 0 0 96 799
use nand3 g8178
timestamp 1386234893
transform 1 0 2499 0 1 1133
box 0 0 120 799
use nand2 state_reg_91_1_93_
timestamp 1386234792
transform 1 0 2619 0 1 1133
box 0 0 96 799
use scandtype g8250
timestamp 1386241841
transform 1 0 2715 0 1 1133
box 0 0 624 799
use nor2 g8148
timestamp 1386235306
transform 1 0 3339 0 1 1133
box 0 0 120 799
use nand2 g7976
timestamp 1386234792
transform 1 0 3459 0 1 1133
box 0 0 96 799
use nand3 g7993
timestamp 1386234893
transform 1 0 3555 0 1 1133
box 0 0 120 799
use nand2 g8211
timestamp 1386234792
transform 1 0 3675 0 1 1133
box 0 0 96 799
use nand2 g8196
timestamp 1386234792
transform 1 0 3771 0 1 1133
box 0 0 96 799
use and2 g8175
timestamp 1386234845
transform 1 0 3867 0 1 1133
box 0 0 120 799
use nand2 g8078
timestamp 1386234792
transform 1 0 3987 0 1 1133
box 0 0 96 799
use nand2 g8093
timestamp 1386234792
transform 1 0 4083 0 1 1133
box 0 0 96 799
use inv g7974
timestamp 1386238110
transform 1 0 4179 0 1 1133
box 0 0 120 799
use and2 g8104
timestamp 1386234845
transform 1 0 4299 0 1 1133
box 0 0 120 799
use nand2 g8307
timestamp 1386234792
transform 1 0 4419 0 1 1133
box 0 0 96 799
use inv g7940
timestamp 1386238110
transform 1 0 4515 0 1 1133
box 0 0 120 799
use nor2 g8160
timestamp 1386235306
transform 1 0 4635 0 1 1133
box 0 0 120 799
use nor2 g8076
timestamp 1386235306
transform 1 0 4755 0 1 1133
box 0 0 120 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 4875 0 1 1133
box 0 0 96 799
use scandtype g8224
timestamp 1386241841
transform 1 0 4971 0 1 1133
box 0 0 624 799
use nand2 g8161
timestamp 1386234792
transform 1 0 5595 0 1 1133
box 0 0 96 799
use nand3 g8094
timestamp 1386234893
transform 1 0 5691 0 1 1133
box 0 0 120 799
use nand3 g7910
timestamp 1386234893
transform 1 0 5811 0 1 1133
box 0 0 120 799
use nand4 g8121
timestamp 1386234936
transform 1 0 5931 0 1 1133
box 0 0 144 799
use and2 g8037
timestamp 1386234845
transform 1 0 6075 0 1 1133
box 0 0 120 799
use nand2 g8266
timestamp 1386234792
transform 1 0 6195 0 1 1133
box 0 0 96 799
use and2 g8189
timestamp 1386234845
transform 1 0 6291 0 1 1133
box 0 0 120 799
use nand3 g8125
timestamp 1386234893
transform 1 0 6411 0 1 1133
box 0 0 120 799
use inv g7915
timestamp 1386238110
transform 1 0 6531 0 1 1133
box 0 0 120 799
use nand4 g8232
timestamp 1386234936
transform 1 0 6651 0 1 1133
box 0 0 144 799
use inv g8152
timestamp 1386238110
transform 1 0 6795 0 1 1133
box 0 0 120 799
use nand2 g8303
timestamp 1386234792
transform 1 0 6915 0 1 1133
box 0 0 96 799
use inv g8080
timestamp 1386238110
transform 1 0 7011 0 1 1133
box 0 0 120 799
use nand2 g7937
timestamp 1386234792
transform 1 0 7131 0 1 1133
box 0 0 96 799
use nand4 g7997
timestamp 1386234936
transform 1 0 7227 0 1 1133
box 0 0 144 799
use nand3 g8282
timestamp 1386234893
transform 1 0 7371 0 1 1133
box 0 0 120 799
use nor2 g8267
timestamp 1386235306
transform 1 0 7491 0 1 1133
box 0 0 120 799
use and2 g8274
timestamp 1386234845
transform 1 0 7611 0 1 1133
box 0 0 120 799
use nand2 g8236
timestamp 1386234792
transform 1 0 7731 0 1 1133
box 0 0 96 799
use nand2 g8101
timestamp 1386234792
transform 1 0 7827 0 1 1133
box 0 0 96 799
use nand2 g8011
timestamp 1386234792
transform 1 0 7923 0 1 1133
box 0 0 96 799
use nand2 g7919
timestamp 1386234792
transform 1 0 8019 0 1 1133
box 0 0 96 799
use nor2 g8185
timestamp 1386235306
transform 1 0 8115 0 1 1133
box 0 0 120 799
use nand2 IntReq_reg
timestamp 1386234792
transform 1 0 8235 0 1 1133
box 0 0 96 799
use scandtype g7927
timestamp 1386241841
transform 1 0 8331 0 1 1133
box 0 0 624 799
use nand4 g8255
timestamp 1386234936
transform 1 0 8955 0 1 1133
box 0 0 144 799
use inv g8086
timestamp 1386238110
transform 1 0 9099 0 1 1133
box 0 0 120 799
use nand2 g8301
timestamp 1386234792
transform 1 0 9219 0 1 1133
box 0 0 96 799
use inv g7962
timestamp 1386238110
transform 1 0 9315 0 1 1133
box 0 0 120 799
use inv g8192
timestamp 1386238110
transform 1 0 9435 0 1 1133
box 0 0 120 799
use nand2 g7988
timestamp 1386234792
transform 1 0 9555 0 1 1133
box 0 0 96 799
use nor2 g8292
timestamp 1386235306
transform 1 0 9651 0 1 1133
box 0 0 120 799
use nor2 g8254
timestamp 1386235306
transform 1 0 9771 0 1 1133
box 0 0 120 799
use nand2 g8116
timestamp 1386234792
transform 1 0 9891 0 1 1133
box 0 0 96 799
use nand2 g8166
timestamp 1386234792
transform 1 0 9987 0 1 1133
box 0 0 96 799
use nand2 g8145
timestamp 1386234792
transform 1 0 10083 0 1 1133
box 0 0 96 799
use and2 g8014
timestamp 1386234845
transform 1 0 10179 0 1 1133
box 0 0 120 799
use nand2 g7959
timestamp 1386234792
transform 1 0 10299 0 1 1133
box 0 0 96 799
use nand3 g8001
timestamp 1386234893
transform 1 0 10395 0 1 1133
box 0 0 120 799
use nand3 g7998
timestamp 1386234893
transform 1 0 10515 0 1 1133
box 0 0 120 799
use nand2 g8228
timestamp 1386234792
transform 1 0 10635 0 1 1133
box 0 0 96 799
use and2 g8072
timestamp 1386234845
transform 1 0 10731 0 1 1133
box 0 0 120 799
use nor2 g7966
timestamp 1386235306
transform 1 0 10851 0 1 1133
box 0 0 120 799
use nand4 g8279
timestamp 1386234936
transform 1 0 10971 0 1 1133
box 0 0 144 799
use nand2 g8105
timestamp 1386234792
transform 1 0 11115 0 1 1133
box 0 0 96 799
use nand2 g8259
timestamp 1386234792
transform 1 0 11211 0 1 1133
box 0 0 96 799
use nand2 g8129
timestamp 1386234792
transform 1 0 11307 0 1 1133
box 0 0 96 799
use nand2 g8122
timestamp 1386234792
transform 1 0 11403 0 1 1133
box 0 0 96 799
use nand2 g8059
timestamp 1386234792
transform 1 0 11499 0 1 1133
box 0 0 96 799
use nand2 g8097
timestamp 1386234792
transform 1 0 11595 0 1 1133
box 0 0 96 799
use nand2 g8062
timestamp 1386234792
transform 1 0 11691 0 1 1133
box 0 0 96 799
use nand3 g8025
timestamp 1386234893
transform 1 0 11787 0 1 1133
box 0 0 120 799
use nand2 g8247
timestamp 1386234792
transform 1 0 11907 0 1 1133
box 0 0 96 799
use nand2 g8263
timestamp 1386234792
transform 1 0 12003 0 1 1133
box 0 0 96 799
use nor2 g8131
timestamp 1386235306
transform 1 0 12099 0 1 1133
box 0 0 120 799
use nand3 g8256
timestamp 1386234893
transform 1 0 12219 0 1 1133
box 0 0 120 799
use nand2 g8087
timestamp 1386234792
transform 1 0 12339 0 1 1133
box 0 0 96 799
use inv g7970
timestamp 1386238110
transform 1 0 12435 0 1 1133
box 0 0 120 799
use rowcrosser Flags_91_3_93_
timestamp 1386086759
transform 1 0 12555 0 1 1133
box 0 0 48 799
use nand2 g7932
timestamp 1386234792
transform 1 0 12603 0 1 1133
box 0 0 96 799
use nand2 g8286
timestamp 1386234792
transform 1 0 12699 0 1 1133
box 0 0 96 799
use and2 g7991
timestamp 1386234845
transform 1 0 12795 0 1 1133
box 0 0 120 799
use nand2 g8137
timestamp 1386234792
transform 1 0 12915 0 1 1133
box 0 0 96 799
use nand4 g8201
timestamp 1386234936
transform 1 0 13011 0 1 1133
box 0 0 144 799
use nand2 g7936
timestamp 1386234792
transform 1 0 13155 0 1 1133
box 0 0 96 799
use nor2 g8242
timestamp 1386235306
transform 1 0 13251 0 1 1133
box 0 0 120 799
use nand2 g8207
timestamp 1386234792
transform 1 0 13371 0 1 1133
box 0 0 96 799
use nand2 g8044
timestamp 1386234792
transform 1 0 13467 0 1 1133
box 0 0 96 799
use nand3 g8006
timestamp 1386234893
transform 1 0 13563 0 1 1133
box 0 0 120 799
use nand3 g8173
timestamp 1386234893
transform 1 0 13683 0 1 1133
box 0 0 120 799
use nand2 g7983
timestamp 1386234792
transform 1 0 13803 0 1 1133
box 0 0 96 799
use nand4 g8157
timestamp 1386234936
transform 1 0 13899 0 1 1133
box 0 0 144 799
use nand2 g7956
timestamp 1386234792
transform 1 0 14043 0 1 1133
box 0 0 96 799
use nand2 g8040
timestamp 1386234792
transform 1 0 14139 0 1 1133
box 0 0 96 799
use nand2 g8068
timestamp 1386234792
transform 1 0 14235 0 1 1133
box 0 0 96 799
use nand2 g8140
timestamp 1386234792
transform 1 0 14331 0 1 1133
box 0 0 96 799
use nand4 g452
timestamp 1386234936
transform 1 0 14427 0 1 1133
box 0 0 144 799
use trisbuf g8141
timestamp 1386237216
transform 1 0 14571 0 1 1133
box 0 0 216 799
use mux2 g8210
timestamp 1386235218
transform 1 0 14787 0 1 1133
box 0 0 192 799
use nand2 InISR_reg
timestamp 1386234792
transform 1 0 14979 0 1 1133
box 0 0 96 799
use scandtype g8003
timestamp 1386241841
transform 1 0 15075 0 1 1133
box 0 0 624 799
use and2 g8203
timestamp 1386234845
transform 1 0 15699 0 1 1133
box 0 0 120 799
use nand2 g8065
timestamp 1386234792
transform 1 0 15819 0 1 1133
box 0 0 96 799
use nand2 g8113
timestamp 1386234792
transform 1 0 15915 0 1 1133
box 0 0 96 799
use nand2 g7977
timestamp 1386234792
transform 1 0 16011 0 1 1133
box 0 0 96 799
use nand3 g8070
timestamp 1386234893
transform 1 0 16107 0 1 1133
box 0 0 120 799
use nand2 g8038
timestamp 1386234792
transform 1 0 16227 0 1 1133
box 0 0 96 799
use nand2 g8233
timestamp 1386234792
transform 1 0 16323 0 1 1133
box 0 0 96 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 16419 0 1 1133
box 0 0 48 799
use nor2 IRQ2_reg
timestamp 1386235306
transform 1 0 16467 0 1 1133
box 0 0 120 799
use scandtype g7980
timestamp 1386241841
transform 1 0 16587 0 1 1133
box 0 0 624 799
use nand3 g7954
timestamp 1386234893
transform 1 0 17211 0 1 1133
box 0 0 120 799
use nand2 g7920
timestamp 1386234792
transform 1 0 17331 0 1 1133
box 0 0 96 799
use nand3 g8151
timestamp 1386234893
transform 1 0 17427 0 1 1133
box 0 0 120 799
use nand2 g7968
timestamp 1386234792
transform 1 0 17547 0 1 1133
box 0 0 96 799
use and2 g8138
timestamp 1386234845
transform 1 0 17643 0 1 1133
box 0 0 120 799
use nand3 g8188
timestamp 1386234893
transform 1 0 17763 0 1 1133
box 0 0 120 799
use inv g8176
timestamp 1386238110
transform 1 0 17883 0 1 1133
box 0 0 120 799
use nand2 g8172
timestamp 1386234792
transform 1 0 18003 0 1 1133
box 0 0 96 799
use nand2 g8026
timestamp 1386234792
transform 1 0 18099 0 1 1133
box 0 0 96 799
use inv g8162
timestamp 1386238110
transform 1 0 18195 0 1 1133
box 0 0 120 799
use inv g8031
timestamp 1386238110
transform 1 0 18315 0 1 1133
box 0 0 120 799
use and2 g7935
timestamp 1386234845
transform 1 0 18435 0 1 1133
box 0 0 120 799
use nand4 g8095
timestamp 1386234936
transform 1 0 18555 0 1 1133
box 0 0 144 799
use and2 g7950
timestamp 1386234845
transform 1 0 18699 0 1 1133
box 0 0 120 799
use nand3 g8013
timestamp 1386234893
transform 1 0 18819 0 1 1133
box 0 0 120 799
use nand2 g8126
timestamp 1386234792
transform 1 0 18939 0 1 1133
box 0 0 96 799
use nand2 g7984
timestamp 1386234792
transform 1 0 19035 0 1 1133
box 0 0 96 799
use inv IRQ1_reg
timestamp 1386238110
transform 1 0 19131 0 1 1133
box 0 0 120 799
use scandtype g7986
timestamp 1386241841
transform 1 0 19251 0 1 1133
box 0 0 624 799
use nand2 g8205
timestamp 1386234792
transform 1 0 19875 0 1 1133
box 0 0 96 799
use nand2 g8164
timestamp 1386234792
transform 1 0 19971 0 1 1133
box 0 0 96 799
use inv g7949
timestamp 1386238110
transform 1 0 20067 0 1 1133
box 0 0 120 799
use nand4 g8017
timestamp 1386234936
transform 1 0 20187 0 1 1133
box 0 0 144 799
use nand2 g8165
timestamp 1386234792
transform 1 0 20331 0 1 1133
box 0 0 96 799
use nand2 g8010
timestamp 1386234792
transform 1 0 20427 0 1 1133
box 0 0 96 799
use nand2 g8260
timestamp 1386234792
transform 1 0 20523 0 1 1133
box 0 0 96 799
use inv g8245
timestamp 1386238110
transform 1 0 20619 0 1 1133
box 0 0 120 799
use nand3 g8034
timestamp 1386234893
transform 1 0 20739 0 1 1133
box 0 0 120 799
use nand2 g8215
timestamp 1386234792
transform 1 0 20859 0 1 1133
box 0 0 96 799
use nand2 g8079
timestamp 1386234792
transform 1 0 20955 0 1 1133
box 0 0 96 799
use nand2 g7999
timestamp 1386234792
transform 1 0 21051 0 1 1133
box 0 0 96 799
use nand3 g8239
timestamp 1386234893
transform 1 0 21147 0 1 1133
box 0 0 120 799
use nand2 g8288
timestamp 1386234792
transform 1 0 21267 0 1 1133
box 0 0 96 799
use nand2 g8007
timestamp 1386234792
transform 1 0 21363 0 1 1133
box 0 0 96 799
use nand4 g8262
timestamp 1386234936
transform 1 0 21459 0 1 1133
box 0 0 144 799
use nor2 g7965
timestamp 1386235306
transform 1 0 21603 0 1 1133
box 0 0 120 799
use nand4 g8109
timestamp 1386234936
transform 1 0 21723 0 1 1133
box 0 0 144 799
use nand3 g8085
timestamp 1386234893
transform 1 0 21867 0 1 1133
box 0 0 120 799
use and2 g8298
timestamp 1386234845
transform 1 0 21987 0 1 1133
box 0 0 120 799
use inv g7944
timestamp 1386238110
transform 1 0 22107 0 1 1133
box 0 0 120 799
use nand2 g8021
timestamp 1386234792
transform 1 0 22227 0 1 1133
box 0 0 96 799
use nand2 g7961
timestamp 1386234792
transform 1 0 22323 0 1 1133
box 0 0 96 799
use nand3 g7931
timestamp 1386234893
transform 1 0 22419 0 1 1133
box 0 0 120 799
use nand2 g8184
timestamp 1386234792
transform 1 0 22539 0 1 1133
box 0 0 96 799
use nand2 g7938
timestamp 1386234792
transform 1 0 22635 0 1 1133
box 0 0 96 799
use nand4 g8132
timestamp 1386234936
transform 1 0 22731 0 1 1133
box 0 0 144 799
use nand2 g8219
timestamp 1386234792
transform 1 0 22875 0 1 1133
box 0 0 96 799
use inv g7916
timestamp 1386238110
transform 1 0 22971 0 1 1133
box 0 0 120 799
use nand4 g8061
timestamp 1386234936
transform 1 0 23091 0 1 1133
box 0 0 144 799
use nand2 g8258
timestamp 1386234792
transform 1 0 23235 0 1 1133
box 0 0 96 799
use inv g8115
timestamp 1386238110
transform 1 0 23331 0 1 1133
box 0 0 120 799
use nand2 g8202
timestamp 1386234792
transform 1 0 23451 0 1 1133
box 0 0 96 799
use nand2 g7973
timestamp 1386234792
transform 1 0 23547 0 1 1133
box 0 0 96 799
use and2 g453
timestamp 1386234845
transform 1 0 23643 0 1 1133
box 0 0 120 799
use trisbuf g8246
timestamp 1386237216
transform 1 0 23763 0 1 1133
box 0 0 216 799
use xor2 g8208
timestamp 1386237344
transform 1 0 23979 0 1 1133
box 0 0 192 799
use nand2 g7958
timestamp 1386234792
transform 1 0 24171 0 1 1133
box 0 0 96 799
use nand2 g8156
timestamp 1386234792
transform 1 0 24267 0 1 1133
box 0 0 96 799
use nand2 g8231
timestamp 1386234792
transform 1 0 24363 0 1 1133
box 0 0 96 799
use nand2 g8047
timestamp 1386234792
transform 1 0 24459 0 1 1133
box 0 0 96 799
use nand2 g7992
timestamp 1386234792
transform 1 0 24555 0 1 1133
box 0 0 96 799
use nand2 g7957
timestamp 1386234792
transform 1 0 24651 0 1 1133
box 0 0 96 799
use nand2 g8179
timestamp 1386234792
transform 1 0 24747 0 1 1133
box 0 0 96 799
use and2 g8022
timestamp 1386234845
transform 1 0 24843 0 1 1133
box 0 0 120 799
use nand2 g8071
timestamp 1386234792
transform 1 0 24963 0 1 1133
box 0 0 96 799
use nand2 g8285
timestamp 1386234792
transform 1 0 25059 0 1 1133
box 0 0 96 799
use nand2 g8083
timestamp 1386234792
transform 1 0 25155 0 1 1133
box 0 0 96 799
use nand3 g7953
timestamp 1386234893
transform 1 0 25251 0 1 1133
box 0 0 120 799
use nor2 g8204
timestamp 1386235306
transform 1 0 25371 0 1 1133
box 0 0 120 799
use nand2 g8053
timestamp 1386234792
transform 1 0 25491 0 1 1133
box 0 0 96 799
use mux2 g8000
timestamp 1386235218
transform 1 0 25587 0 1 1133
box 0 0 192 799
use nand2 state_reg_91_0_93_
timestamp 1386234792
transform 1 0 25779 0 1 1133
box 0 0 96 799
use scandtype g8142
timestamp 1386241841
transform 1 0 25875 0 1 1133
box 0 0 624 799
use mux2 g8302
timestamp 1386235218
transform 1 0 26499 0 1 1133
box 0 0 192 799
use inv stateSub_reg_91_1_93_
timestamp 1386238110
transform 1 0 26691 0 1 1133
box 0 0 120 799
use scandtype Flags_91_0_93_
timestamp 1386241841
transform 1 0 26811 0 1 1133
box 0 0 624 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 27795 0 1 1133
box 0 0 320 799
<< labels >>
rlabel m2contact 27873 8614 27873 8614 6 RwSel[0]
rlabel m2contact 27873 8542 27873 8542 6 RwSel[0]
rlabel m2contact 27849 8710 27849 8710 6 CFlag
rlabel m2contact 27849 8590 27849 8590 6 CFlag
rlabel m2contact 27849 8542 27849 8542 6 Rs1Sel[1]
rlabel m2contact 27849 8518 27849 8518 6 Rs1Sel[1]
rlabel m2contact 27825 8590 27825 8590 6 Rs1Sel[0]
rlabel m2contact 27825 8470 27825 8470 6 Rs1Sel[0]
rlabel m2contact 27801 8518 27801 8518 6 RwSel[1]
rlabel m2contact 27801 8494 27801 8494 6 RwSel[1]
rlabel m2contact 27801 8470 27801 8470 6 AluOR[0]
rlabel m2contact 27801 8446 27801 8446 6 AluOR[0]
rlabel m2contact 27777 8518 27777 8518 6 RwSel[1]
rlabel m2contact 27729 8566 27729 8566 6 RegWe
rlabel m2contact 26277 8566 26277 8566 6 MemEn
rlabel m2contact 25785 8638 25785 8638 6 ALE
rlabel m2contact 25569 8494 25569 8494 6 PcSel[2]
rlabel m2contact 24741 8782 24741 8782 6 IrWe
rlabel m2contact 23841 8662 23841 8662 6 LrEn
rlabel m2contact 23205 8758 23205 8758 6 LrSel
rlabel m2contact 23193 8518 23193 8518 6 PcEn
rlabel m2contact 22857 8446 22857 8446 6 PcSel[1]
rlabel m2contact 21669 8686 21669 8686 6 LrWe
rlabel m2contact 20133 8734 20133 8734 6 WdSel
rlabel m2contact 20109 8662 20109 8662 6 LrEn
rlabel m2contact 18873 8662 18873 8662 6 Op1Sel
rlabel m2contact 18825 8782 18825 8782 6 IrWe
rlabel m2contact 18681 8710 18681 8710 6 CFlag
rlabel m2contact 17061 8710 17061 8710 6 PcSel[0]
rlabel m2contact 17037 8446 17037 8446 6 PcSel[1]
rlabel m2contact 16929 8758 16929 8758 6 LrSel
rlabel m2contact 16833 8470 16833 8470 6 AluOR[0]
rlabel m2contact 15501 8494 15501 8494 6 PcSel[2]
rlabel m2contact 13953 8518 13953 8518 4 PcEn
rlabel m2contact 13377 8734 13377 8734 4 WdSel
rlabel m2contact 13041 8710 13041 8710 4 PcSel[0]
rlabel m2contact 12681 8686 12681 8686 4 LrWe
rlabel metal2 12267 8686 12267 8686 4 PcWe
rlabel m2contact 12249 8686 12249 8686 4 PcWe
rlabel m2contact 11097 8566 11097 8566 4 MemEn
rlabel m2contact 10857 8662 10857 8662 4 Op1Sel
rlabel m2contact 10353 8590 10353 8590 4 Rs1Sel[0]
rlabel m2contact 9225 8590 9225 8590 4 AluEn
rlabel metal2 8763 8566 8763 8566 4 ImmSel
rlabel m2contact 8745 8566 8745 8566 4 ImmSel
rlabel m2contact 7833 8566 7833 8566 4 AluWe
rlabel metal2 7155 8662 7155 8662 4 Op2Sel[0]
rlabel m2contact 7137 8662 7137 8662 4 Op2Sel[0]
rlabel m2contact 7089 8542 7089 8542 4 Rs1Sel[1]
rlabel m2contact 6945 8614 6945 8614 4 RwSel[0]
rlabel m2contact 4701 8614 4701 8614 4 Op2Sel[1]
rlabel m2contact 4665 8566 4665 8566 4 AluWe
rlabel m2contact 3117 8590 3117 8590 4 AluEn
rlabel m2contact 2865 8614 2865 8614 4 Op2Sel[1]
rlabel m2contact 1761 8590 1761 8590 4 nWait
rlabel m2contact 1713 8614 1713 8614 4 nME
rlabel m2contact 26865 324 26865 324 8 OpcodeCondIn[2]
rlabel m2contact 26865 108 26865 108 8 OpcodeCondIn[2]
rlabel m2contact 26841 588 26841 588 8 OpcodeCondIn[7]
rlabel m2contact 26841 84 26841 84 8 OpcodeCondIn[7]
rlabel m2contact 26817 924 26817 924 6 OpcodeCondIn[6]
rlabel m2contact 26817 60 26817 60 8 OpcodeCondIn[6]
rlabel m2contact 26793 300 26793 300 8 OpcodeCondIn[4]
rlabel m2contact 26793 36 26793 36 8 OpcodeCondIn[4]
rlabel m2contact 26769 660 26769 660 8 OpcodeCondIn[5]
rlabel m2contact 26769 12 26769 12 8 OpcodeCondIn[5]
rlabel m2contact 26739 228 26739 228 8 OpcodeCondIn[0]
rlabel m2contact 26733 132 26733 132 8 OpcodeCondIn[0]
rlabel m2contact 26721 228 26721 228 8 OpcodeCondIn[0]
rlabel m2contact 26625 180 26625 180 8 n_43
rlabel m2contact 26577 924 26577 924 6 OpcodeCondIn[6]
rlabel m2contact 25977 852 25977 852 6 n_368
rlabel m2contact 25857 372 25857 372 8 n_262
rlabel m2contact 25809 828 25809 828 6 n_199
rlabel m2contact 25737 948 25737 948 6 n_248
rlabel m2contact 25425 396 25425 396 8 n_295
rlabel m2contact 24729 636 24729 636 8 n_289
rlabel m2contact 24633 612 24633 612 8 n_334
rlabel m2contact 24393 756 24393 756 8 n_116
rlabel m2contact 24345 900 24345 900 6 n_283
rlabel m2contact 24129 684 24129 684 8 n_36
rlabel m2contact 24009 660 24009 660 8 OpcodeCondIn[5]
rlabel m2contact 23697 540 23697 540 8 n_234
rlabel m2contact 23625 732 23625 732 8 n_331
rlabel m2contact 23529 708 23529 708 8 n_146
rlabel m2contact 23505 660 23505 660 8 OpcodeCondIn[5]
rlabel m2contact 23169 468 23169 468 8 n_370
rlabel m2contact 23049 348 23049 348 8 n_109
rlabel m2contact 22905 564 22905 564 8 n_44
rlabel m2contact 22809 1020 22809 1020 6 n_286
rlabel m2contact 22785 612 22785 612 8 n_334
rlabel m2contact 22713 780 22713 780 8 n_130
rlabel m2contact 22377 1068 22377 1068 6 n_238
rlabel m2contact 22305 972 22305 972 6 n_350
rlabel m2contact 22281 84 22281 84 8 Flags[1]
rlabel m2contact 22137 660 22137 660 8 OpcodeCondIn[5]
rlabel m2contact 21969 1116 21969 1116 6 n_69
rlabel m2contact 21945 924 21945 924 6 OpcodeCondIn[6]
rlabel m2contact 21921 684 21921 684 8 n_36
rlabel m2contact 21897 300 21897 300 8 OpcodeCondIn[4]
rlabel m2contact 21777 276 21777 276 8 n_308
rlabel m2contact 21753 708 21753 708 8 n_146
rlabel m2contact 21417 324 21417 324 8 OpcodeCondIn[2]
rlabel m2contact 21321 924 21321 924 6 OpcodeCondIn[6]
rlabel m2contact 21249 708 21249 708 8 n_263
rlabel m2contact 21177 756 21177 756 8 n_116
rlabel m2contact 21129 156 21129 156 8 n_180
rlabel m2contact 21105 804 21105 804 6 n_102
rlabel m2contact 21033 252 21033 252 8 n_52
rlabel m2contact 20841 108 20841 108 8 n_10
rlabel m2contact 20817 228 20817 228 8 OpcodeCondIn[0]
rlabel m2contact 20505 492 20505 492 8 n_152
rlabel m2contact 20313 852 20313 852 6 n_368
rlabel m2contact 20265 852 20265 852 6 n_89
rlabel m2contact 20145 444 20145 444 8 n_153
rlabel m2contact 20097 492 20097 492 8 n_152
rlabel m2contact 19953 36 19953 36 8 n_292
rlabel m2contact 19905 132 19905 132 8 n_191
rlabel m2contact 19761 60 19761 60 8 IRQ1
rlabel m2contact 19353 420 19353 420 8 n_1
rlabel m2contact 19113 516 19113 516 8 n_195
rlabel m2contact 19065 780 19065 780 8 n_130
rlabel m2contact 19017 1044 19017 1044 6 n_220
rlabel m2contact 18921 204 18921 204 8 n_288
rlabel m2contact 18873 1092 18873 1092 6 n_193
rlabel m2contact 18657 780 18657 780 8 n_179
rlabel m2contact 18633 900 18633 900 6 n_283
rlabel m2contact 18609 876 18609 876 6 n_261
rlabel m2contact 18489 324 18489 324 8 OpcodeCondIn[2]
rlabel m2contact 18057 924 18057 924 6 OpcodeCondIn[6]
rlabel m2contact 18033 684 18033 684 8 n_36
rlabel m2contact 17913 684 17913 684 8 n_85
rlabel m2contact 17865 996 17865 996 6 n_67
rlabel m2contact 17673 708 17673 708 8 n_263
rlabel m2contact 17601 708 17601 708 8 n_48
rlabel m2contact 17577 900 17577 900 6 n_25
rlabel m2contact 17481 972 17481 972 6 n_350
rlabel m2contact 17289 156 17289 156 8 n_180
rlabel m2contact 17265 972 17265 972 6 n_218
rlabel m2contact 17241 1044 17241 1044 6 n_220
rlabel m2contact 17049 156 17049 156 8 n_492
rlabel m2contact 16689 60 16689 60 8 IRQ1
rlabel m2contact 16569 756 16569 756 8 n_116
rlabel m2contact 16449 12 16449 12 8 Flags[0]
rlabel m2contact 16281 1044 16281 1044 6 n_38
rlabel m2contact 16257 1116 16257 1116 6 n_69
rlabel m2contact 16209 1092 16209 1092 6 n_193
rlabel m2contact 15993 1068 15993 1068 6 n_238
rlabel m2contact 15897 1044 15897 1044 6 n_38
rlabel m2contact 15801 1020 15801 1020 6 n_286
rlabel m2contact 15057 180 15057 180 8 n_43
rlabel m2contact 14937 804 14937 804 6 n_102
rlabel m2contact 14361 804 14361 804 4 n_141
rlabel m2contact 14073 348 14073 348 2 n_109
rlabel m2contact 13953 348 13953 348 2 n_242
rlabel m2contact 13785 876 13785 876 4 n_261
rlabel m2contact 13665 876 13665 876 4 n_192
rlabel m2contact 13641 180 13641 180 2 n_113
rlabel m2contact 13449 708 13449 708 2 n_48
rlabel m2contact 13353 708 13353 708 2 n_269
rlabel m2contact 12849 660 12849 660 2 OpcodeCondIn[5]
rlabel m2contact 12825 924 12825 924 4 OpcodeCondIn[6]
rlabel m2contact 12633 36 12633 36 2 n_292
rlabel m2contact 12585 36 12585 36 2 Flags[2]
rlabel m2contact 12417 900 12417 900 4 n_25
rlabel m2contact 12153 588 12153 588 2 OpcodeCondIn[7]
rlabel m2contact 11889 348 11889 348 2 n_242
rlabel m2contact 11865 444 11865 444 2 n_153
rlabel m2contact 11721 996 11721 996 4 n_67
rlabel m2contact 11673 996 11673 996 4 n_245
rlabel m2contact 11529 492 11529 492 2 n_152
rlabel m2contact 11481 804 11481 804 4 n_141
rlabel m2contact 11433 348 11433 348 2 n_93
rlabel m2contact 11097 444 11097 444 2 n_327
rlabel m2contact 11073 804 11073 804 4 n_145
rlabel m2contact 11049 636 11049 636 2 n_289
rlabel m2contact 11001 636 11001 636 2 n_271
rlabel m2contact 10833 492 10833 492 2 n_59
rlabel m2contact 10785 660 10785 660 2 OpcodeCondIn[5]
rlabel m2contact 10617 276 10617 276 2 n_308
rlabel m2contact 10449 276 10449 276 2 n_309
rlabel m2contact 10425 996 10425 996 4 n_245
rlabel m2contact 10377 972 10377 972 4 n_218
rlabel m2contact 10065 804 10065 804 4 n_145
rlabel m2contact 9753 804 9753 804 4 n_290
rlabel m2contact 9681 948 9681 948 4 n_248
rlabel m2contact 9345 924 9345 924 4 OpcodeCondIn[6]
rlabel m2contact 9129 900 9129 900 4 n_25
rlabel m2contact 8433 876 8433 876 4 n_192
rlabel m2contact 8313 852 8313 852 4 n_89
rlabel m2contact 8097 828 8097 828 4 n_199
rlabel m2contact 8073 588 8073 588 2 OpcodeCondIn[7]
rlabel m2contact 7665 588 7665 588 2 OpcodeCondIn[7]
rlabel m2contact 7329 732 7329 732 2 n_331
rlabel m2contact 7305 804 7305 804 4 n_290
rlabel m2contact 7209 780 7209 780 2 n_179
rlabel m2contact 7185 492 7185 492 2 n_59
rlabel m2contact 6945 780 6945 780 2 n_106
rlabel m2contact 6873 780 6873 780 2 n_106
rlabel m2contact 6825 756 6825 756 2 n_116
rlabel m2contact 6753 732 6753 732 2 n_331
rlabel m2contact 6729 708 6729 708 2 n_269
rlabel m2contact 6561 516 6561 516 2 n_195
rlabel m2contact 6513 684 6513 684 2 n_85
rlabel m2contact 6345 660 6345 660 2 OpcodeCondIn[5]
rlabel m2contact 6273 636 6273 636 2 n_271
rlabel m2contact 5961 612 5961 612 2 n_334
rlabel m2contact 5889 588 5889 588 2 OpcodeCondIn[7]
rlabel m2contact 5793 564 5793 564 2 n_44
rlabel m2contact 4953 540 4953 540 2 n_234
rlabel m2contact 4929 516 4929 516 2 n_195
rlabel m2contact 4809 492 4809 492 2 n_59
rlabel m2contact 4737 468 4737 468 2 n_370
rlabel m2contact 4665 444 4665 444 2 n_327
rlabel m2contact 4593 420 4593 420 2 n_1
rlabel m2contact 4401 396 4401 396 2 n_295
rlabel m2contact 4329 372 4329 372 2 n_262
rlabel m2contact 4065 348 4065 348 2 n_93
rlabel m2contact 4041 324 4041 324 2 OpcodeCondIn[2]
rlabel m2contact 3825 300 3825 300 2 OpcodeCondIn[4]
rlabel m2contact 3753 276 3753 276 2 n_309
rlabel m2contact 3513 252 3513 252 2 n_52
rlabel m2contact 3369 228 3369 228 2 OpcodeCondIn[0]
rlabel m2contact 2817 204 2817 204 2 n_288
rlabel m2contact 2697 180 2697 180 2 n_113
rlabel m2contact 2673 156 2673 156 2 n_492
rlabel m2contact 2649 60 2649 60 2 IRQ1
rlabel m2contact 1761 60 1761 60 2 Flags[3]
rlabel m2contact 1713 132 1713 132 2 n_191
rlabel m2contact 1641 108 1641 108 2 n_10
rlabel m2contact 27897 4421 27897 4421 6 SysBus[1]
rlabel m2contact 27897 2069 27897 2069 6 SysBus[1]
rlabel m2contact 27873 6365 27873 6365 6 SysBus[0]
rlabel m2contact 27873 2045 27873 2045 6 SysBus[0]
rlabel m2contact 27849 3509 27849 3509 6 SysBus[3]
rlabel m2contact 27849 2021 27849 2021 6 SysBus[3]
rlabel m2contact 27825 4565 27825 4565 6 SysBus[2]
rlabel m2contact 27825 1997 27825 1997 6 SysBus[2]
rlabel m2contact 27801 4685 27801 4685 6 OpcodeCondIn[3]
rlabel m2contact 27801 1973 27801 1973 6 OpcodeCondIn[3]
rlabel m2contact 27777 3485 27777 3485 6 OpcodeCondIn[1]
rlabel m2contact 27777 1949 27777 1949 6 OpcodeCondIn[1]
rlabel m2contact 27777 4325 27777 4325 6 RwSel[1]
rlabel m2contact 27729 4469 27729 4469 6 RegWe
rlabel m2contact 27681 2237 27681 2237 6 n_20
rlabel m2contact 27633 3869 27633 3869 6 stateSub[0]
rlabel m2contact 27609 4781 27609 4781 6 n_258
rlabel m2contact 27561 4397 27561 4397 6 n_241
rlabel m2contact 27537 3797 27537 3797 6 n_275
rlabel m2contact 27513 2717 27513 2717 6 n_240
rlabel m2contact 27465 6893 27465 6893 6 n_115
rlabel m2contact 27441 6197 27441 6197 6 n_105
rlabel m2contact 27417 3797 27417 3797 6 n_275
rlabel m2contact 27369 4493 27369 4493 6 n_342
rlabel m2contact 27345 5885 27345 5885 6 n_19
rlabel m2contact 27321 6029 27321 6029 6 n_291
rlabel m2contact 27321 3101 27321 3101 6 stateSub[1]
rlabel m2contact 27297 7085 27297 7085 6 n_70
rlabel m2contact 27273 1949 27273 1949 6 n_18
rlabel m2contact 27249 5021 27249 5021 6 n_166
rlabel m2contact 27225 6461 27225 6461 6 n_185
rlabel m2contact 27201 5285 27201 5285 6 n_225
rlabel m2contact 27177 3701 27177 3701 6 n_63
rlabel m2contact 27129 4637 27129 4637 6 n_49
rlabel m2contact 27105 2141 27105 2141 6 n_16
rlabel m2contact 27081 6533 27081 6533 6 n_26
rlabel m2contact 27009 6461 27009 6461 6 n_185
rlabel m2contact 26961 4661 26961 4661 6 OpcodeCondIn[7]
rlabel m2contact 26937 5597 26937 5597 6 n_103
rlabel m2contact 26937 4541 26937 4541 6 n_103
rlabel m2contact 26913 5597 26913 5597 6 n_103
rlabel m2contact 26913 5573 26913 5573 6 n_373
rlabel m2contact 26889 3557 26889 3557 6 state[1]
rlabel m2contact 26865 7133 26865 7133 6 n_95
rlabel m2contact 26817 4133 26817 4133 6 n_183
rlabel m2contact 26793 5885 26793 5885 6 n_19
rlabel m2contact 26793 4613 26793 4613 6 n_19
rlabel m2contact 26769 4613 26769 4613 6 n_19
rlabel m2contact 26769 4685 26769 4685 6 OpcodeCondIn[3]
rlabel m2contact 26745 5285 26745 5285 6 n_225
rlabel m2contact 26697 4829 26697 4829 6 n_50
rlabel m2contact 26673 3797 26673 3797 6 n_275
rlabel m2contact 26649 3125 26649 3125 6 n_121
rlabel m2contact 26649 5357 26649 5357 6 n_287
rlabel m2contact 26577 3509 26577 3509 6 SysBus[3]
rlabel m2contact 26553 3797 26553 3797 6 n_275
rlabel m2contact 26505 6341 26505 6341 6 n_224
rlabel m2contact 26433 4085 26433 4085 6 StatusReg[3]
rlabel m2contact 26409 5837 26409 5837 6 n_96
rlabel m2contact 26409 3149 26409 3149 6 n_96
rlabel m2contact 26385 4757 26385 4757 6 n_212
rlabel m2contact 26385 3749 26385 3749 6 state[0]
rlabel m2contact 26361 4181 26361 4181 6 n_182
rlabel m2contact 26337 3149 26337 3149 6 n_96
rlabel m2contact 26337 3173 26337 3173 6 n_211
rlabel m2contact 26289 2333 26289 2333 6 n_379
rlabel m2contact 26265 4277 26265 4277 6 n_66
rlabel m2contact 26241 4733 26241 4733 6 n_344
rlabel m2contact 26217 3077 26217 3077 6 n_186
rlabel m2contact 26193 2117 26193 2117 6 n_148
rlabel m2contact 26145 2549 26145 2549 6 n_338
rlabel m2contact 26121 2093 26121 2093 6 n_337
rlabel m2contact 26097 4421 26097 4421 6 SysBus[1]
rlabel m2contact 26025 6557 26025 6557 6 n_120
rlabel m2contact 25977 3437 25977 3437 6 n_119
rlabel m2contact 25929 6629 25929 6629 6 n_249
rlabel m2contact 25905 5741 25905 5741 6 OpcodeCondIn[2]
rlabel m2contact 25881 5285 25881 5285 6 n_225
rlabel m2contact 25857 5429 25857 5429 6 n_227
rlabel m2contact 25833 5693 25833 5693 6 n_158
rlabel m2contact 25833 3749 25833 3749 6 state[0]
rlabel m2contact 25785 7493 25785 7493 6 PcSel[2]
rlabel m2contact 25785 4229 25785 4229 6 PcSel[2]
rlabel m2contact 25761 5765 25761 5765 6 n_320
rlabel m2contact 25737 4709 25737 4709 6 n_135
rlabel m2contact 25713 5069 25713 5069 6 n_247
rlabel m2contact 25689 7061 25689 7061 6 n_47
rlabel m2contact 25665 3557 25665 3557 6 state[1]
rlabel m2contact 25641 3101 25641 3101 6 stateSub[1]
rlabel m2contact 25641 4685 25641 4685 6 OpcodeCondIn[3]
rlabel m2contact 25617 2597 25617 2597 6 n_303
rlabel m2contact 25593 5237 25593 5237 6 n_150
rlabel m2contact 25593 4109 25593 4109 6 n_150
rlabel m2contact 25569 7493 25569 7493 6 PcSel[2]
rlabel m2contact 25569 7469 25569 7469 6 n_32
rlabel m2contact 25545 3461 25545 3461 6 n_122
rlabel m2contact 25521 5933 25521 5933 6 n_22
rlabel m2contact 25521 3797 25521 3797 6 n_275
rlabel m2contact 25497 7133 25497 7133 6 n_95
rlabel m2contact 25473 4733 25473 4733 6 n_344
rlabel m2contact 25449 6605 25449 6605 6 n_184
rlabel m2contact 25425 4613 25425 4613 6 n_197
rlabel m2contact 25401 4109 25401 4109 6 n_150
rlabel m2contact 25401 4133 25401 4133 6 n_183
rlabel m2contact 25353 2861 25353 2861 6 n_207
rlabel m2contact 25353 4373 25353 4373 6 n_229
rlabel m2contact 25329 3269 25329 3269 6 n_206
rlabel m2contact 25305 3197 25305 3197 6 n_187
rlabel m2contact 25305 3869 25305 3869 6 stateSub[0]
rlabel m2contact 25281 2477 25281 2477 6 n_132
rlabel m2contact 25281 3557 25281 3557 6 state[1]
rlabel m2contact 25257 5381 25257 5381 6 n_364
rlabel m2contact 25257 4109 25257 4109 6 n_364
rlabel m2contact 25233 5381 25233 5381 6 n_364
rlabel m2contact 25233 5357 25233 5357 6 n_287
rlabel m2contact 25209 6821 25209 6821 6 n_363
rlabel m2contact 25209 3557 25209 3557 6 state[1]
rlabel m2contact 25185 6269 25185 6269 6 n_346
rlabel m2contact 25185 3749 25185 3749 6 state[0]
rlabel m2contact 25161 4853 25161 4853 6 n_71
rlabel m2contact 25161 3029 25161 3029 6 n_71
rlabel m2contact 25137 5405 25137 5405 6 n_235
rlabel m2contact 25113 4853 25113 4853 6 n_71
rlabel m2contact 25113 4805 25113 4805 6 n_255
rlabel m2contact 25089 4997 25089 4997 6 n_108
rlabel m2contact 25041 4853 25041 4853 6 n_217
rlabel m2contact 25017 5525 25017 5525 6 OpcodeCondIn[0]
rlabel m2contact 25017 3389 25017 3389 6 n_215
rlabel m2contact 24993 7085 24993 7085 6 n_70
rlabel m2contact 24993 6869 24993 6869 6 n_216
rlabel m2contact 24957 5189 24957 5189 6 n_226
rlabel m2contact 24957 4733 24957 4733 6 n_226
rlabel m2contact 24945 5261 24945 5261 6 n_107
rlabel m2contact 24945 2045 24945 2045 6 n_137
rlabel m2contact 24921 4517 24921 4517 6 n_251
rlabel m2contact 24897 4733 24897 4733 6 n_226
rlabel m2contact 24897 5093 24897 5093 6 n_228
rlabel m2contact 24873 4517 24873 4517 6 n_251
rlabel m2contact 24825 3653 24825 3653 6 n_329
rlabel m2contact 24825 4445 24825 4445 6 n_324
rlabel m2contact 24801 2093 24801 2093 6 n_337
rlabel m2contact 24777 3509 24777 3509 6 SysBus[3]
rlabel m2contact 24777 3533 24777 3533 6 n_323
rlabel m2contact 24741 4877 24741 4877 6 n_187
rlabel m2contact 24741 3197 24741 3197 6 n_187
rlabel m2contact 24729 5285 24729 5285 6 n_225
rlabel m2contact 24705 5501 24705 5501 6 n_221
rlabel m2contact 24681 4757 24681 4757 6 n_212
rlabel m2contact 24681 5981 24681 5981 6 stateSub[2]
rlabel m2contact 24657 6917 24657 6917 6 n_231
rlabel m2contact 24633 5117 24633 5117 6 n_126
rlabel m2contact 24633 3221 24633 3221 6 n_126
rlabel m2contact 24609 4877 24609 4877 6 n_187
rlabel m2contact 24609 4685 24609 4685 6 OpcodeCondIn[3]
rlabel m2contact 24585 2693 24585 2693 6 n_270
rlabel m2contact 24561 5669 24561 5669 6 OpcodeCondIn[4]
rlabel m2contact 24537 5213 24537 5213 6 n_76
rlabel m2contact 24537 5285 24537 5285 6 n_225
rlabel m2contact 24513 5357 24513 5357 6 n_287
rlabel m2contact 24489 5117 24489 5117 6 n_126
rlabel m2contact 24489 5093 24489 5093 6 n_228
rlabel m2contact 24465 4685 24465 4685 6 OpcodeCondIn[3]
rlabel m2contact 24441 4733 24441 4733 6 n_42
rlabel m2contact 24441 3509 24441 3509 6 n_117
rlabel m2contact 24417 4901 24417 4901 6 n_7
rlabel m2contact 24417 5333 24417 5333 6 n_12
rlabel m2contact 24393 3101 24393 3101 6 stateSub[1]
rlabel m2contact 24369 7517 24369 7517 6 n_209
rlabel m2contact 24369 4757 24369 4757 6 n_209
rlabel m2contact 24345 5141 24345 5141 6 n_213
rlabel m2contact 24321 4013 24321 4013 6 n_60
rlabel m2contact 24321 3269 24321 3269 6 n_206
rlabel m2contact 24297 4757 24297 4757 6 n_209
rlabel m2contact 24297 4973 24297 4973 6 n_219
rlabel m2contact 24273 7541 24273 7541 6 n_54
rlabel m2contact 24273 2285 24273 2285 6 n_54
rlabel m2contact 24249 2285 24249 2285 6 n_54
rlabel m2contact 24249 2309 24249 2309 6 n_124
rlabel m2contact 24225 7421 24225 7421 6 n_28
rlabel m2contact 24225 2597 24225 2597 6 n_303
rlabel m2contact 24201 7205 24201 7205 6 n_65
rlabel m2contact 24201 5909 24201 5909 6 n_24
rlabel m2contact 24153 4757 24153 4757 6 n_319
rlabel m2contact 24129 4685 24129 4685 6 OpcodeCondIn[3]
rlabel m2contact 24105 4589 24105 4589 6 n_280
rlabel m2contact 24069 4877 24069 4877 6 OpcodeCondIn[1]
rlabel m2contact 24069 3485 24069 3485 6 OpcodeCondIn[1]
rlabel m2contact 24057 4901 24057 4901 6 n_7
rlabel m2contact 24033 4877 24033 4877 6 OpcodeCondIn[1]
rlabel m2contact 24033 4685 24033 4685 6 OpcodeCondIn[3]
rlabel m2contact 24009 5741 24009 5741 6 OpcodeCondIn[2]
rlabel m2contact 23961 4205 23961 4205 6 n_256
rlabel m2contact 23937 4421 23937 4421 6 SysBus[1]
rlabel m2contact 23937 4805 23937 4805 6 n_255
rlabel m2contact 23913 5093 23913 5093 6 n_228
rlabel m2contact 23889 4781 23889 4781 6 n_258
rlabel m2contact 23865 6341 23865 6341 6 n_224
rlabel m2contact 23841 6485 23841 6485 6 n_342
rlabel m2contact 23841 4493 23841 4493 6 n_342
rlabel m2contact 23817 5309 23817 5309 6 n_250
rlabel m2contact 23793 6485 23793 6485 6 n_342
rlabel m2contact 23793 6437 23793 6437 6 CFlag
rlabel m2contact 23745 6509 23745 6509 6 n_353
rlabel m2contact 23721 7445 23721 7445 6 n_159
rlabel m2contact 23673 4757 23673 4757 6 n_319
rlabel m2contact 23673 6845 23673 6845 6 n_189
rlabel m2contact 23649 4877 23649 4877 6 n_171
rlabel m2contact 23649 2741 23649 2741 6 n_171
rlabel m2contact 23625 4757 23625 4757 6 n_181
rlabel m2contact 23601 4877 23601 4877 6 n_171
rlabel m2contact 23601 3701 23601 3701 6 n_63
rlabel m2contact 23577 3749 23577 3749 6 state[0]
rlabel m2contact 23577 4133 23577 4133 6 n_183
rlabel m2contact 23553 5165 23553 5165 6 n_81
rlabel m2contact 23553 4349 23553 4349 6 n_81
rlabel m2contact 23529 4061 23529 4061 6 n_35
rlabel m2contact 23505 6149 23505 6149 6 n_253
rlabel m2contact 23505 4301 23505 4301 6 n_253
rlabel m2contact 23481 5645 23481 5645 6 OpcodeCondIn[6]
rlabel m2contact 23481 5285 23481 5285 6 n_225
rlabel m2contact 23457 2909 23457 2909 6 n_34
rlabel m2contact 23433 7493 23433 7493 6 n_188
rlabel m2contact 23433 4421 23433 4421 6 n_188
rlabel m2contact 23409 5165 23409 5165 6 n_81
rlabel m2contact 23409 5117 23409 5117 6 n_84
rlabel m2contact 23385 5381 23385 5381 6 n_80
rlabel m2contact 23361 4301 23361 4301 6 n_253
rlabel m2contact 23361 5117 23361 5117 6 n_84
rlabel m2contact 23337 4877 23337 4877 6 n_316
rlabel m2contact 23337 2357 23337 2357 6 n_316
rlabel m2contact 23313 4421 23313 4421 6 n_188
rlabel m2contact 23313 5165 23313 5165 6 n_260
rlabel m2contact 23289 6461 23289 6461 6 n_185
rlabel m2contact 23265 3197 23265 3197 6 n_187
rlabel m2contact 23265 4901 23265 4901 6 n_157
rlabel m2contact 23241 4133 23241 4133 6 n_183
rlabel m2contact 23217 4469 23217 4469 6 RegWe
rlabel m2contact 23193 6821 23193 6821 6 n_363
rlabel m2contact 23169 4421 23169 4421 6 n_366
rlabel m2contact 23145 4877 23145 4877 6 n_316
rlabel m2contact 23145 3149 23145 3149 6 n_384
rlabel m2contact 23121 4853 23121 4853 6 n_217
rlabel m2contact 23121 2525 23121 2525 6 n_335
rlabel m2contact 23073 3317 23073 3317 6 n_88
rlabel m2contact 23049 3461 23049 3461 6 n_122
rlabel m2contact 23025 1973 23025 1973 6 n_41
rlabel m2contact 23001 2621 23001 2621 6 n_306
rlabel m2contact 22977 4925 22977 4925 6 n_140
rlabel m2contact 22977 3365 22977 3365 6 n_140
rlabel m2contact 22953 3365 22953 3365 6 n_140
rlabel m2contact 22953 3389 22953 3389 6 n_215
rlabel m2contact 22929 4901 22929 4901 6 n_157
rlabel m2contact 22905 3701 22905 3701 6 n_63
rlabel m2contact 22857 4325 22857 4325 6 RwSel[1]
rlabel m2contact 22857 4469 22857 4469 6 PcSel[1]
rlabel m2contact 22833 6821 22833 6821 6 n_363
rlabel m2contact 22761 2525 22761 2525 6 n_335
rlabel m2contact 22713 6317 22713 6317 6 StatusReg[0]
rlabel m2contact 22689 4901 22689 4901 6 n_157
rlabel m2contact 22665 5717 22665 5717 6 n_496
rlabel m2contact 22665 5189 22665 5189 6 n_226
rlabel m2contact 22617 6005 22617 6005 6 n_312
rlabel m2contact 22593 2885 22593 2885 6 StatusReg[2]
rlabel m2contact 22569 6989 22569 6989 6 n_313
rlabel m2contact 22521 4469 22521 4469 6 PcSel[1]
rlabel m2contact 22497 4877 22497 4877 6 n_356
rlabel m2contact 22473 4493 22473 4493 6 n_342
rlabel m2contact 22449 6245 22449 6245 6 n_345
rlabel m2contact 22401 3917 22401 3917 6 n_274
rlabel m2contact 22353 4637 22353 4637 6 n_49
rlabel m2contact 22305 7349 22305 7349 6 n_374
rlabel m2contact 22257 7037 22257 7037 6 n_349
rlabel m2contact 22185 5501 22185 5501 6 n_221
rlabel m2contact 22161 5549 22161 5549 6 n_86
rlabel m2contact 22137 5669 22137 5669 6 OpcodeCondIn[4]
rlabel m2contact 22137 3725 22137 3725 6 OpcodeCondIn[4]
rlabel m2contact 22113 4829 22113 4829 6 n_50
rlabel m2contact 22089 2693 22089 2693 6 n_270
rlabel m2contact 22065 7253 22065 7253 6 n_75
rlabel m2contact 22065 3773 22065 3773 6 n_75
rlabel m2contact 22041 5429 22041 5429 6 n_227
rlabel m2contact 22041 5045 22041 5045 6 n_266
rlabel m2contact 22017 4637 22017 4637 6 n_232
rlabel m2contact 21993 4949 21993 4949 6 n_172
rlabel m2contact 21957 4853 21957 4853 6 n_303
rlabel m2contact 21957 2597 21957 2597 6 n_303
rlabel m2contact 21945 6389 21945 6389 6 n_17
rlabel m2contact 21921 5837 21921 5837 6 n_96
rlabel m2contact 21897 3725 21897 3725 6 OpcodeCondIn[4]
rlabel m2contact 21897 3845 21897 3845 6 n_110
rlabel m2contact 21873 5861 21873 5861 6 n_305
rlabel m2contact 21873 3821 21873 3821 6 n_305
rlabel m2contact 21849 3989 21849 3989 6 n_355
rlabel m2contact 21849 6245 21849 6245 6 n_345
rlabel m2contact 21825 4853 21825 4853 6 n_303
rlabel m2contact 21825 3605 21825 3605 6 n_94
rlabel m2contact 21801 4301 21801 4301 6 n_297
rlabel m2contact 21801 2381 21801 2381 6 n_223
rlabel m2contact 21765 4853 21765 4853 6 n_91
rlabel m2contact 21765 2789 21765 2789 6 n_91
rlabel m2contact 21753 5333 21753 5333 6 n_12
rlabel m2contact 21729 5741 21729 5741 6 OpcodeCondIn[2]
rlabel m2contact 21705 3773 21705 3773 6 n_75
rlabel m2contact 21705 3869 21705 3869 6 stateSub[0]
rlabel m2contact 21681 4469 21681 4469 6 n_136
rlabel m2contact 21657 3485 21657 3485 6 OpcodeCondIn[1]
rlabel m2contact 21633 6101 21633 6101 6 n_257
rlabel m2contact 21633 5885 21633 5885 6 n_19
rlabel m2contact 21609 6197 21609 6197 6 n_105
rlabel m2contact 21609 4493 21609 4493 6 n_105
rlabel m2contact 21585 3821 21585 3821 6 n_305
rlabel m2contact 21585 3869 21585 3869 6 stateSub[0]
rlabel m2contact 21561 4349 21561 4349 6 n_81
rlabel m2contact 21561 5093 21561 5093 6 n_228
rlabel m2contact 21537 2933 21537 2933 6 n_97
rlabel m2contact 21513 2789 21513 2789 6 n_91
rlabel m2contact 21513 2813 21513 2813 6 n_296
rlabel m2contact 21489 3365 21489 3365 6 n_293
rlabel m2contact 21465 5333 21465 5333 6 n_142
rlabel m2contact 21441 6485 21441 6485 6 n_205
rlabel m2contact 21441 5789 21441 5789 6 n_15
rlabel m2contact 21417 5165 21417 5165 6 n_260
rlabel m2contact 21417 3725 21417 3725 6 n_260
rlabel m2contact 21393 7181 21393 7181 6 n_6
rlabel m2contact 21393 4685 21393 4685 6 OpcodeCondIn[3]
rlabel m2contact 21369 7589 21369 7589 6 n_194
rlabel m2contact 21369 2261 21369 2261 6 n_194
rlabel m2contact 21345 4493 21345 4493 6 n_105
rlabel m2contact 21345 4685 21345 4685 6 OpcodeCondIn[3]
rlabel m2contact 21321 7277 21321 7277 6 OpcodeCondIn[5]
rlabel m2contact 21297 3389 21297 3389 6 n_215
rlabel m2contact 21273 7373 21273 7373 6 n_310
rlabel m2contact 21249 5405 21249 5405 6 n_235
rlabel m2contact 21225 5141 21225 5141 6 n_213
rlabel m2contact 21225 2597 21225 2597 6 n_303
rlabel m2contact 21201 3725 21201 3725 6 n_260
rlabel m2contact 21201 3773 21201 3773 6 n_276
rlabel m2contact 21165 5429 21165 5429 6 n_227
rlabel m2contact 21165 4349 21165 4349 6 n_227
rlabel m2contact 21153 7013 21153 7013 6 n_315
rlabel m2contact 21129 6317 21129 6317 6 StatusReg[0]
rlabel m2contact 21105 6989 21105 6989 6 n_313
rlabel m2contact 21081 3197 21081 3197 6 n_187
rlabel m2contact 21057 5453 21057 5453 6 n_165
rlabel m2contact 21057 4493 21057 4493 6 n_165
rlabel m2contact 21033 4997 21033 4997 6 n_108
rlabel m2contact 21009 2477 21009 2477 6 n_132
rlabel m2contact 20985 5261 20985 5261 6 n_107
rlabel m2contact 20985 3749 20985 3749 6 state[0]
rlabel m2contact 20961 6413 20961 6413 6 n_40
rlabel m2contact 20961 4997 20961 4997 6 n_40
rlabel m2contact 20937 2261 20937 2261 6 n_194
rlabel m2contact 20937 2285 20937 2285 6 n_155
rlabel m2contact 20913 4349 20913 4349 6 n_227
rlabel m2contact 20913 4661 20913 4661 6 OpcodeCondIn[7]
rlabel m2contact 20889 4493 20889 4493 6 n_165
rlabel m2contact 20889 5285 20889 5285 6 n_225
rlabel m2contact 20865 7253 20865 7253 6 n_75
rlabel m2contact 20841 2597 20841 2597 6 n_303
rlabel m2contact 20817 5525 20817 5525 6 OpcodeCondIn[0]
rlabel m2contact 20793 6413 20793 6413 6 n_40
rlabel m2contact 20793 6317 20793 6317 6 StatusReg[0]
rlabel m2contact 20769 5477 20769 5477 6 n_493
rlabel m2contact 20769 3485 20769 3485 6 OpcodeCondIn[1]
rlabel m2contact 20745 2885 20745 2885 6 StatusReg[2]
rlabel m2contact 20721 5621 20721 5621 6 n_100
rlabel m2contact 20721 2429 20721 2429 6 n_100
rlabel m2contact 20697 5765 20697 5765 6 n_320
rlabel m2contact 20697 5693 20697 5693 6 n_158
rlabel m2contact 20673 6173 20673 6173 6 n_277
rlabel m2contact 20649 6101 20649 6101 6 n_257
rlabel m2contact 20649 5909 20649 5909 6 n_24
rlabel m2contact 20625 5597 20625 5597 6 n_99
rlabel m2contact 20625 3293 20625 3293 6 n_99
rlabel m2contact 20601 3005 20601 3005 6 n_282
rlabel m2contact 20601 4421 20601 4421 6 n_366
rlabel m2contact 20577 4781 20577 4781 6 n_258
rlabel m2contact 20553 6749 20553 6749 6 n_74
rlabel m2contact 20553 4349 20553 4349 6 n_281
rlabel m2contact 20529 5141 20529 5141 6 n_77
rlabel m2contact 20505 5405 20505 5405 6 n_104
rlabel m2contact 20505 2189 20505 2189 6 n_104
rlabel m2contact 20481 5621 20481 5621 6 n_100
rlabel m2contact 20481 4685 20481 4685 6 OpcodeCondIn[3]
rlabel m2contact 20457 5597 20457 5597 6 n_99
rlabel m2contact 20457 4901 20457 4901 6 n_157
rlabel m2contact 20433 5189 20433 5189 6 n_226
rlabel m2contact 20409 4589 20409 4589 6 n_280
rlabel m2contact 20385 6725 20385 6725 6 n_239
rlabel m2contact 20361 5405 20361 5405 6 n_104
rlabel m2contact 20361 2789 20361 2789 6 n_279
rlabel m2contact 20337 6413 20337 6413 6 n_23
rlabel m2contact 20337 2669 20337 2669 6 n_23
rlabel m2contact 20313 5765 20313 5765 6 n_61
rlabel m2contact 20289 5357 20289 5357 6 n_287
rlabel m2contact 20265 5309 20265 5309 6 n_250
rlabel m2contact 20241 5813 20241 5813 6 n_203
rlabel m2contact 20241 3941 20241 3941 6 n_321
rlabel m2contact 20217 2669 20217 2669 6 n_23
rlabel m2contact 20217 2717 20217 2717 6 n_240
rlabel m2contact 20193 5045 20193 5045 6 n_266
rlabel m2contact 20145 5597 20145 5597 6 n_164
rlabel m2contact 20097 2213 20097 2213 6 n_14
rlabel m2contact 20073 5405 20073 5405 6 n_118
rlabel m2contact 20049 4733 20049 4733 6 n_42
rlabel m2contact 20025 4157 20025 4157 6 n_78
rlabel m2contact 20001 5309 20001 5309 6 n_156
rlabel m2contact 20001 3797 20001 3797 6 n_275
rlabel m2contact 19953 6965 19953 6965 6 n_170
rlabel m2contact 19929 6029 19929 6029 6 n_291
rlabel m2contact 19905 5957 19905 5957 6 n_45
rlabel m2contact 19857 3485 19857 3485 6 OpcodeCondIn[1]
rlabel m2contact 19833 6461 19833 6461 6 n_185
rlabel m2contact 19785 6869 19785 6869 6 n_216
rlabel m2contact 19737 6053 19737 6053 6 n_177
rlabel m2contact 19713 6845 19713 6845 6 n_189
rlabel m2contact 19665 4253 19665 4253 6 n_162
rlabel m2contact 19641 4493 19641 4493 6 n_161
rlabel m2contact 19617 2069 19617 2069 6 n_127
rlabel m2contact 19569 5189 19569 5189 6 n_226
rlabel m2contact 19521 5525 19521 5525 6 OpcodeCondIn[0]
rlabel m2contact 19497 7085 19497 7085 6 n_70
rlabel m2contact 19449 4325 19449 4325 6 n_139
rlabel m2contact 19425 2261 19425 2261 6 n_21
rlabel m2contact 19401 6221 19401 6221 6 n_58
rlabel m2contact 19377 5213 19377 5213 6 n_76
rlabel m2contact 19341 3965 19341 3965 6 n_351
rlabel m2contact 19341 3245 19341 3245 6 n_351
rlabel m2contact 19329 7037 19329 7037 6 n_349
rlabel m2contact 19305 2405 19305 2405 6 n_144
rlabel m2contact 19281 5525 19281 5525 6 n_222
rlabel m2contact 19257 5021 19257 5021 6 n_166
rlabel m2contact 19233 6293 19233 6293 6 n_178
rlabel m2contact 19209 3629 19209 3629 6 n_362
rlabel m2contact 19185 6125 19185 6125 6 n_31
rlabel m2contact 19161 3245 19161 3245 6 n_351
rlabel m2contact 19161 3269 19161 3269 6 n_206
rlabel m2contact 19137 3749 19137 3749 6 state[0]
rlabel m2contact 19113 6965 19113 6965 6 n_170
rlabel m2contact 19113 4733 19113 4733 6 n_170
rlabel m2contact 19089 4733 19089 4733 6 n_170
rlabel m2contact 19089 6773 19089 6773 6 n_298
rlabel m2contact 19065 4589 19065 4589 6 n_174
rlabel m2contact 19041 5021 19041 5021 6 n_264
rlabel m2contact 19017 5213 19017 5213 6 n_82
rlabel m2contact 19017 2645 19017 2645 6 n_82
rlabel m2contact 18993 5573 18993 5573 6 n_373
rlabel m2contact 18993 3389 18993 3389 6 n_215
rlabel m2contact 18969 5213 18969 5213 6 n_82
rlabel m2contact 18969 4973 18969 4973 6 n_219
rlabel m2contact 18945 4733 18945 4733 6 n_328
rlabel m2contact 18921 5573 18921 5573 6 n_87
rlabel m2contact 18897 5357 18897 5357 6 n_287
rlabel m2contact 18873 3893 18873 3893 6 Op1Sel
rlabel m2contact 18849 4541 18849 4541 6 n_103
rlabel m2contact 18825 4037 18825 4037 6 IrWe
rlabel m2contact 18801 4349 18801 4349 6 n_281
rlabel m2contact 18753 3101 18753 3101 6 stateSub[1]
rlabel m2contact 18729 4541 18729 4541 6 n_244
rlabel m2contact 18681 6437 18681 6437 6 CFlag
rlabel m2contact 18681 3581 18681 3581 6 n_326
rlabel m2contact 18585 5213 18585 5213 6 n_167
rlabel m2contact 18537 2093 18537 2093 6 n_337
rlabel m2contact 18489 5741 18489 5741 6 OpcodeCondIn[2]
rlabel m2contact 18465 4301 18465 4301 6 n_297
rlabel m2contact 18393 4877 18393 4877 6 n_356
rlabel m2contact 18345 4229 18345 4229 6 PcSel[2]
rlabel m2contact 18273 3893 18273 3893 6 Op1Sel
rlabel m2contact 18273 4229 18273 4229 6 n_375
rlabel m2contact 18225 6077 18225 6077 6 n_299
rlabel m2contact 18201 5621 18201 5621 6 n_37
rlabel m2contact 18201 3893 18201 3893 6 n_37
rlabel m2contact 18177 6821 18177 6821 6 n_363
rlabel m2contact 18153 6917 18153 6917 6 n_231
rlabel m2contact 18153 6701 18153 6701 6 n_90
rlabel m2contact 18129 6101 18129 6101 6 n_257
rlabel m2contact 18105 5381 18105 5381 6 n_80
rlabel m2contact 18081 3893 18081 3893 6 n_37
rlabel m2contact 18081 4517 18081 4517 6 n_251
rlabel m2contact 18045 5501 18045 5501 6 n_221
rlabel m2contact 18045 3893 18045 3893 6 n_221
rlabel m2contact 18033 6413 18033 6413 6 n_23
rlabel m2contact 18009 3749 18009 3749 6 state[0]
rlabel m2contact 17985 7109 17985 7109 6 n_27
rlabel m2contact 17961 4037 17961 4037 6 IrWe
rlabel m2contact 17937 6293 17937 6293 6 n_178
rlabel m2contact 17913 5621 17913 5621 6 n_37
rlabel m2contact 17889 3197 17889 3197 6 n_187
rlabel m2contact 17865 7157 17865 7157 6 n_30
rlabel m2contact 17865 4037 17865 4037 6 n_30
rlabel m2contact 17841 3893 17841 3893 6 n_221
rlabel m2contact 17841 4517 17841 4517 6 n_251
rlabel m2contact 17817 5981 17817 5981 6 stateSub[2]
rlabel m2contact 17793 4037 17793 4037 6 n_30
rlabel m2contact 17793 5837 17793 5837 6 n_96
rlabel m2contact 17769 3557 17769 3557 6 state[1]
rlabel m2contact 17745 6797 17745 6797 6 n_359
rlabel m2contact 17721 5453 17721 5453 6 n_165
rlabel m2contact 17697 5261 17697 5261 6 n_107
rlabel m2contact 17697 2813 17697 2813 6 n_296
rlabel m2contact 17673 1997 17673 1997 6 n_123
rlabel m2contact 17649 7301 17649 7301 6 n_278
rlabel m2contact 17649 3725 17649 3725 6 n_278
rlabel m2contact 17625 7301 17625 7301 6 n_278
rlabel m2contact 17625 7229 17625 7229 6 n_98
rlabel m2contact 17601 2573 17601 2573 6 n_11
rlabel m2contact 17577 2693 17577 2693 6 n_270
rlabel m2contact 17529 4229 17529 4229 6 n_375
rlabel m2contact 17505 2549 17505 2549 6 n_338
rlabel m2contact 17505 2597 17505 2597 6 n_303
rlabel m2contact 17481 7325 17481 7325 6 n_339
rlabel m2contact 17481 4229 17481 4229 6 n_339
rlabel m2contact 17457 5621 17457 5621 6 n_314
rlabel m2contact 17457 5741 17457 5741 6 OpcodeCondIn[2]
rlabel m2contact 17433 6365 17433 6365 6 SysBus[0]
rlabel m2contact 17433 3677 17433 3677 6 SysBus[0]
rlabel m2contact 17409 4229 17409 4229 6 n_339
rlabel m2contact 17409 6581 17409 6581 6 n_268
rlabel m2contact 17385 2093 17385 2093 6 n_337
rlabel m2contact 17385 5045 17385 5045 6 n_266
rlabel m2contact 17361 3677 17361 3677 6 SysBus[0]
rlabel m2contact 17361 3821 17361 3821 6 n_267
rlabel m2contact 17313 7301 17313 7301 6 n_83
rlabel m2contact 17313 2549 17313 2549 6 Op2Sel[0]
rlabel m2contact 17289 3485 17289 3485 6 OpcodeCondIn[1]
rlabel m2contact 17265 5045 17265 5045 6 n_266
rlabel m2contact 17241 4661 17241 4661 6 OpcodeCondIn[7]
rlabel m2contact 17193 5213 17193 5213 6 n_167
rlabel m2contact 17169 4661 17169 4661 6 OpcodeCondIn[7]
rlabel m2contact 17145 5285 17145 5285 6 n_225
rlabel m2contact 17121 3245 17121 3245 6 n_143
rlabel m2contact 17097 6293 17097 6293 6 IRQ2
rlabel m2contact 17073 7397 17073 7397 6 n_230
rlabel m2contact 17049 5429 17049 5429 6 n_227
rlabel m2contact 17025 5093 17025 5093 6 n_228
rlabel m2contact 17001 4373 17001 4373 6 n_229
rlabel m2contact 16881 2021 16881 2021 6 n_301
rlabel m2contact 16833 4229 16833 4229 6 AluOR[0]
rlabel m2contact 16785 3893 16785 3893 6 n_352
rlabel m2contact 16761 4037 16761 4037 6 Flags[0]
rlabel m2contact 16737 7037 16737 7037 6 n_349
rlabel m2contact 16593 5981 16593 5981 6 stateSub[2]
rlabel m2contact 16545 3797 16545 3797 6 n_275
rlabel m2contact 16521 7253 16521 7253 6 n_75
rlabel m2contact 16497 5693 16497 5693 6 n_158
rlabel m2contact 16449 4037 16449 4037 6 Flags[0]
rlabel m2contact 16401 4229 16401 4229 6 AluOR[0]
rlabel m2contact 16377 2621 16377 2621 6 n_306
rlabel m2contact 16353 5453 16353 5453 6 n_284
rlabel m2contact 16305 5213 16305 5213 6 n_128
rlabel m2contact 16185 5861 16185 5861 6 n_305
rlabel m2contact 16185 5381 16185 5381 6 n_80
rlabel m2contact 16161 3341 16161 3341 6 IntReq
rlabel m2contact 16137 4253 16137 4253 6 n_162
rlabel m2contact 16113 5861 16113 5861 6 n_99
rlabel m2contact 16113 3293 16113 3293 6 n_99
rlabel m2contact 16089 5261 16089 5261 6 n_173
rlabel m2contact 16065 4613 16065 4613 6 n_197
rlabel m2contact 16041 5861 16041 5861 6 n_99
rlabel m2contact 16041 4373 16041 4373 6 n_229
rlabel m2contact 16017 6149 16017 6149 6 n_253
rlabel m2contact 16017 4253 16017 4253 6 n_253
rlabel m2contact 15993 5669 15993 5669 6 OpcodeCondIn[4]
rlabel m2contact 15969 6413 15969 6413 6 n_237
rlabel m2contact 15945 4253 15945 4253 6 n_253
rlabel m2contact 15945 5861 15945 5861 6 n_372
rlabel m2contact 15921 4229 15921 4229 6 n_330
rlabel m2contact 15897 7565 15897 7565 6 n_348
rlabel m2contact 15873 6005 15873 6005 6 n_312
rlabel m2contact 15873 4469 15873 4469 6 n_136
rlabel m2contact 15849 4013 15849 4013 6 n_60
rlabel m2contact 15753 4757 15753 4757 6 n_181
rlabel m2contact 15729 4085 15729 4085 6 StatusReg[3]
rlabel m2contact 15729 3413 15729 3413 6 n_210
rlabel m2contact 15681 5477 15681 5477 6 n_493
rlabel m2contact 15585 2765 15585 2765 6 InISR
rlabel m2contact 15537 4253 15537 4253 6 n_495
rlabel m2contact 15321 4757 15321 4757 6 n_371
rlabel m2contact 15201 5405 15201 5405 6 n_118
rlabel m2contact 15177 4109 15177 4109 6 n_364
rlabel m2contact 15153 3749 15153 3749 6 state[0]
rlabel m2contact 15129 6101 15129 6101 6 n_257
rlabel m2contact 15081 6653 15081 6653 6 n_163
rlabel m2contact 15057 5309 15057 5309 6 n_156
rlabel m2contact 15033 3485 15033 3485 6 OpcodeCondIn[1]
rlabel m2contact 15033 4589 15033 4589 6 n_174
rlabel m2contact 15009 5093 15009 5093 6 n_228
rlabel m2contact 15009 4109 15009 4109 6 n_56
rlabel m2contact 14985 5405 14985 5405 6 n_137
rlabel m2contact 14985 2045 14985 2045 6 n_137
rlabel m2contact 14961 4037 14961 4037 6 n_138
rlabel m2contact 14937 5045 14937 5045 6 n_266
rlabel m2contact 14913 5405 14913 5405 6 n_137
rlabel m2contact 14913 2909 14913 2909 6 n_34
rlabel m2contact 14865 4061 14865 4061 6 n_35
rlabel m2contact 14865 5237 14865 5237 6 n_150
rlabel m2contact 14841 6125 14841 6125 6 n_31
rlabel m2contact 14841 5501 14841 5501 6 n_221
rlabel m2contact 14817 6005 14817 6005 6 n_68
rlabel m2contact 14793 2837 14793 2837 6 n_79
rlabel m2contact 14769 3677 14769 3677 6 n_64
rlabel m2contact 14745 4565 14745 4565 6 SysBus[2]
rlabel m2contact 14721 6941 14721 6941 6 n_202
rlabel m2contact 14697 6341 14697 6341 6 n_224
rlabel m2contact 14697 4061 14697 4061 6 n_224
rlabel m2contact 14673 4061 14673 4061 6 n_224
rlabel m2contact 14673 5237 14673 5237 6 n_151
rlabel m2contact 14649 4925 14649 4925 6 n_140
rlabel m2contact 14625 6461 14625 6461 6 n_185
rlabel m2contact 14625 4061 14625 4061 6 n_185
rlabel m2contact 14601 4853 14601 4853 6 n_91
rlabel m2contact 14601 2885 14601 2885 6 StatusReg[2]
rlabel m2contact 14577 5981 14577 5981 6 stateSub[2]
rlabel m2contact 14553 4277 14553 4277 6 n_66
rlabel m2contact 14553 5405 14553 5405 6 n_51
rlabel m2contact 14529 4685 14529 4685 6 OpcodeCondIn[3]
rlabel m2contact 14505 3749 14505 3749 6 state[0]
rlabel m2contact 14505 4157 14505 4157 6 n_78
rlabel m2contact 14481 3845 14481 3845 6 n_110
rlabel m2contact 14457 5645 14457 5645 6 OpcodeCondIn[6]
rlabel m2contact 14457 4157 14457 4157 6 n_78
rlabel m2contact 14433 6461 14433 6461 6 n_185
rlabel m2contact 14409 3077 14409 3077 6 n_186
rlabel m2contact 14385 4061 14385 4061 4 n_185
rlabel m2contact 14385 4277 14385 4277 4 n_214
rlabel m2contact 14349 4853 14349 4853 4 n_275
rlabel m2contact 14349 3797 14349 3797 4 n_275
rlabel m2contact 14337 5837 14337 5837 4 n_96
rlabel m2contact 14313 3077 14313 3077 4 n_154
rlabel m2contact 14313 4853 14313 4853 4 n_275
rlabel m2contact 14289 3749 14289 3749 4 state[0]
rlabel m2contact 14265 3221 14265 3221 4 n_126
rlabel m2contact 14265 5477 14265 5477 4 n_200
rlabel m2contact 14241 4901 14241 4901 4 n_157
rlabel m2contact 14241 4061 14241 4061 4 n_157
rlabel m2contact 14217 4229 14217 4229 4 n_330
rlabel m2contact 14217 4685 14217 4685 4 OpcodeCondIn[3]
rlabel m2contact 14193 2093 14193 2093 4 n_337
rlabel m2contact 14193 2165 14193 2165 4 n_134
rlabel m2contact 14169 4565 14169 4565 4 SysBus[2]
rlabel m2contact 14145 3221 14145 3221 4 n_92
rlabel m2contact 14121 4709 14121 4709 4 n_135
rlabel m2contact 14097 4853 14097 4853 4 n_275
rlabel m2contact 14097 3845 14097 3845 4 n_110
rlabel m2contact 14073 5381 14073 5381 4 n_80
rlabel m2contact 14049 5837 14049 5837 4 n_96
rlabel m2contact 14049 2981 14049 2981 4 n_96
rlabel m2contact 14025 3533 14025 3533 4 n_323
rlabel m2contact 14025 3821 14025 3821 4 n_267
rlabel m2contact 14001 4229 14001 4229 4 n_111
rlabel m2contact 13977 3533 13977 3533 4 n_246
rlabel m2contact 13977 5789 13977 5789 4 n_15
rlabel m2contact 13953 2717 13953 2717 4 n_240
rlabel m2contact 13929 6125 13929 6125 4 n_259
rlabel m2contact 13905 4853 13905 4853 4 n_381
rlabel m2contact 13881 4925 13881 4925 4 n_131
rlabel m2contact 13857 4061 13857 4061 4 n_157
rlabel m2contact 13857 4565 13857 4565 4 n_252
rlabel m2contact 13833 7589 13833 7589 4 n_194
rlabel m2contact 13833 6677 13833 6677 4 n_55
rlabel m2contact 13809 7061 13809 7061 4 n_47
rlabel m2contact 13809 3053 13809 3053 4 n_47
rlabel m2contact 13785 7613 13785 7613 4 n_18
rlabel m2contact 13785 1949 13785 1949 4 n_18
rlabel m2contact 13761 5381 13761 5381 4 n_80
rlabel m2contact 13761 3461 13761 3461 4 n_122
rlabel m2contact 13737 5165 13737 5165 4 n_260
rlabel m2contact 13713 7109 13713 7109 4 n_27
rlabel m2contact 13713 2597 13713 2597 4 n_303
rlabel m2contact 13677 5069 13677 5069 4 n_247
rlabel m2contact 13677 4061 13677 4061 4 n_247
rlabel m2contact 13665 7157 13665 7157 4 n_30
rlabel m2contact 13641 5669 13641 5669 4 OpcodeCondIn[4]
rlabel m2contact 13617 2669 13617 2669 4 n_101
rlabel m2contact 13617 4709 13617 4709 4 n_29
rlabel m2contact 13593 2957 13593 2957 4 n_160
rlabel m2contact 13569 2621 13569 2621 4 n_306
rlabel m2contact 13545 2645 13545 2645 4 n_82
rlabel m2contact 13545 6701 13545 6701 4 n_90
rlabel m2contact 13521 2981 13521 2981 4 n_96
rlabel m2contact 13521 5093 13521 5093 4 n_228
rlabel m2contact 13497 5045 13497 5045 4 n_266
rlabel m2contact 13473 7133 13473 7133 4 n_95
rlabel m2contact 13449 5981 13449 5981 4 stateSub[2]
rlabel m2contact 13425 3053 13425 3053 4 n_47
rlabel m2contact 13425 5381 13425 5381 4 n_80
rlabel m2contact 13401 3797 13401 3797 4 n_275
rlabel m2contact 13377 2981 13377 2981 4 WdSel
rlabel m2contact 13341 6461 13341 6461 4 n_185
rlabel m2contact 13341 2645 13341 2645 4 n_185
rlabel m2contact 13329 6677 13329 6677 4 n_55
rlabel m2contact 13305 4061 13305 4061 4 n_247
rlabel m2contact 13305 4685 13305 4685 4 OpcodeCondIn[3]
rlabel m2contact 13281 6677 13281 6677 4 n_13
rlabel m2contact 13281 3053 13281 3053 4 n_233
rlabel m2contact 13257 7589 13257 7589 4 n_9
rlabel m2contact 13257 2453 13257 2453 4 n_9
rlabel m2contact 13233 7109 13233 7109 4 n_27
rlabel m2contact 13233 6965 13233 6965 4 n_170
rlabel m2contact 13209 3389 13209 3389 4 n_215
rlabel m2contact 13209 3869 13209 3869 4 stateSub[0]
rlabel m2contact 13185 2645 13185 2645 4 n_185
rlabel m2contact 13185 3101 13185 3101 4 stateSub[1]
rlabel m2contact 13161 7133 13161 7133 4 PcSel[0]
rlabel m2contact 13161 4061 13161 4061 4 PcSel[0]
rlabel m2contact 13137 7157 13137 7157 4 n_33
rlabel m2contact 13137 6485 13137 6485 4 n_205
rlabel m2contact 13113 7613 13113 7613 4 n_18
rlabel m2contact 13113 5813 13113 5813 4 n_203
rlabel m2contact 13089 7589 13089 7589 4 n_9
rlabel m2contact 13089 5285 13089 5285 4 n_225
rlabel m2contact 13065 4901 13065 4901 4 n_157
rlabel m2contact 13041 7133 13041 7133 4 PcSel[0]
rlabel m2contact 13041 5693 13041 5693 4 n_158
rlabel m2contact 12993 2981 12993 2981 4 WdSel
rlabel m2contact 12969 7589 12969 7589 4 n_365
rlabel m2contact 12969 7133 12969 7133 4 n_198
rlabel m2contact 12945 3725 12945 3725 4 n_278
rlabel m2contact 12921 3989 12921 3989 4 n_355
rlabel m2contact 12897 3269 12897 3269 4 n_206
rlabel m2contact 12873 2093 12873 2093 4 n_8
rlabel m2contact 12849 7277 12849 7277 4 OpcodeCondIn[5]
rlabel m2contact 12825 3749 12825 3749 4 state[0]
rlabel m2contact 12801 7277 12801 7277 4 Flags[2]
rlabel m2contact 12801 2645 12801 2645 4 Flags[2]
rlabel m2contact 12777 7565 12777 7565 4 n_348
rlabel m2contact 12777 3725 12777 3725 4 n_311
rlabel m2contact 12753 7277 12753 7277 4 Flags[2]
rlabel m2contact 12753 4085 12753 4085 4 StatusReg[3]
rlabel m2contact 12729 7037 12729 7037 4 n_349
rlabel m2contact 12729 6989 12729 6989 4 n_313
rlabel m2contact 12681 4061 12681 4061 4 PcSel[0]
rlabel m2contact 12657 7565 12657 7565 4 n_204
rlabel m2contact 12657 4877 12657 4877 4 n_356
rlabel m2contact 12633 2021 12633 2021 4 n_301
rlabel m2contact 12585 2645 12585 2645 4 Flags[2]
rlabel m2contact 12585 3389 12585 3389 4 n_332
rlabel m2contact 12537 6149 12537 6149 4 n_253
rlabel m2contact 12513 4301 12513 4301 4 n_297
rlabel m2contact 12513 5357 12513 5357 4 n_287
rlabel m2contact 12489 7277 12489 7277 4 n_39
rlabel m2contact 12489 3989 12489 3989 4 n_39
rlabel m2contact 12465 2525 12465 2525 4 n_335
rlabel m2contact 12465 4301 12465 4301 4 n_265
rlabel m2contact 12441 4925 12441 4925 4 n_131
rlabel m2contact 12417 2645 12417 2645 4 n_196
rlabel m2contact 12393 1949 12393 1949 4 n_18
rlabel m2contact 12393 4061 12393 4061 4 n_175
rlabel m2contact 12369 3797 12369 3797 4 n_275
rlabel m2contact 12345 6845 12345 6845 4 n_189
rlabel m2contact 12321 1997 12321 1997 4 n_123
rlabel m2contact 12321 4925 12321 4925 4 n_129
rlabel m2contact 12297 5285 12297 5285 4 n_225
rlabel m2contact 12297 3461 12297 3461 4 n_122
rlabel m2contact 12273 6917 12273 6917 4 n_231
rlabel m2contact 12249 2597 12249 2597 4 n_303
rlabel m2contact 12225 4877 12225 4877 4 n_356
rlabel m2contact 12201 7589 12201 7589 4 n_365
rlabel m2contact 12201 2909 12201 2909 4 n_34
rlabel m2contact 12177 3149 12177 3149 4 n_384
rlabel m2contact 12153 3173 12153 3173 4 n_211
rlabel m2contact 12129 4685 12129 4685 4 OpcodeCondIn[3]
rlabel m2contact 12105 7565 12105 7565 4 n_204
rlabel m2contact 12093 4997 12093 4997 4 n_40
rlabel m2contact 12093 1997 12093 1997 4 n_40
rlabel m2contact 12081 1973 12081 1973 4 n_41
rlabel m2contact 12081 5813 12081 5813 4 n_203
rlabel m2contact 12057 3989 12057 3989 4 n_39
rlabel m2contact 12057 6917 12057 6917 4 n_231
rlabel m2contact 12033 1997 12033 1997 4 n_40
rlabel m2contact 12033 3797 12033 3797 4 n_275
rlabel m2contact 12009 4613 12009 4613 4 n_197
rlabel m2contact 11985 2021 11985 2021 4 n_301
rlabel m2contact 11985 5189 11985 5189 4 n_226
rlabel m2contact 11985 3989 11985 3989 4 n_226
rlabel m2contact 11961 3989 11961 3989 4 n_226
rlabel m2contact 11961 4541 11961 4541 4 n_244
rlabel m2contact 11937 6029 11937 6029 4 n_291
rlabel m2contact 11913 4949 11913 4949 4 n_172
rlabel m2contact 11889 7469 11889 7469 4 n_32
rlabel m2contact 11841 2045 11841 2045 4 n_137
rlabel m2contact 11841 3989 11841 3989 4 n_147
rlabel m2contact 11817 5045 11817 5045 4 n_266
rlabel m2contact 11793 7541 11793 7541 4 n_54
rlabel m2contact 11793 7469 11793 7469 4 n_143
rlabel m2contact 11793 3245 11793 3245 4 n_143
rlabel m2contact 11769 2069 11769 2069 4 n_127
rlabel m2contact 11769 3317 11769 3317 4 n_88
rlabel m2contact 11745 3749 11745 3749 4 state[0]
rlabel m2contact 11721 7517 11721 7517 4 n_209
rlabel m2contact 11721 6965 11721 6965 4 n_170
rlabel m2contact 11721 3317 11721 3317 4 n_170
rlabel m2contact 11697 6845 11697 6845 4 n_189
rlabel m2contact 11673 2285 11673 2285 4 n_155
rlabel m2contact 11649 7493 11649 7493 4 n_188
rlabel m2contact 11649 4781 11649 4781 4 n_258
rlabel m2contact 11625 4541 11625 4541 4 n_244
rlabel m2contact 11601 2405 11601 2405 4 n_144
rlabel m2contact 11577 7469 11577 7469 4 n_143
rlabel m2contact 11577 4805 11577 4805 4 n_255
rlabel m2contact 11553 3317 11553 3317 4 n_170
rlabel m2contact 11553 5285 11553 5285 4 n_225
rlabel m2contact 11529 6149 11529 6149 4 n_253
rlabel m2contact 11529 2405 11529 2405 4 n_253
rlabel m2contact 11505 3365 11505 3365 4 n_293
rlabel m2contact 11481 2285 11481 2285 4 n_176
rlabel m2contact 11457 2093 11457 2093 4 n_8
rlabel m2contact 11457 4277 11457 4277 4 n_214
rlabel m2contact 11433 5837 11433 5837 4 n_96
rlabel m2contact 11433 3317 11433 3317 4 n_96
rlabel m2contact 11409 2789 11409 2789 4 n_279
rlabel m2contact 11385 2405 11385 2405 4 n_253
rlabel m2contact 11385 5309 11385 5309 4 n_156
rlabel m2contact 11361 6101 11361 6101 4 n_257
rlabel m2contact 11361 4781 11361 4781 4 n_258
rlabel m2contact 11337 3317 11337 3317 4 n_96
rlabel m2contact 11337 4517 11337 4517 4 n_251
rlabel m2contact 11313 7469 11313 7469 4 n_149
rlabel m2contact 11313 2405 11313 2405 4 n_149
rlabel m2contact 11289 2117 11289 2117 4 n_148
rlabel m2contact 11289 3317 11289 3317 4 n_208
rlabel m2contact 11265 7469 11265 7469 4 n_149
rlabel m2contact 11265 5501 11265 5501 4 n_221
rlabel m2contact 11241 7445 11241 7445 4 n_159
rlabel m2contact 11241 3437 11241 3437 4 n_119
rlabel m2contact 11193 2141 11193 2141 4 n_16
rlabel m2contact 11193 7421 11193 7421 4 n_28
rlabel m2contact 11169 5981 11169 5981 4 stateSub[2]
rlabel m2contact 11169 3845 11169 3845 4 n_110
rlabel m2contact 11145 7109 11145 7109 4 n_27
rlabel m2contact 11145 3797 11145 3797 4 n_275
rlabel m2contact 11073 7397 11073 7397 4 n_230
rlabel m2contact 11049 3005 11049 3005 4 n_282
rlabel m2contact 11025 3317 11025 3317 4 n_208
rlabel m2contact 11025 3917 11025 3917 4 n_274
rlabel m2contact 10977 5621 10977 5621 4 n_314
rlabel m2contact 10953 6437 10953 6437 4 CFlag
rlabel m2contact 10953 6341 10953 6341 4 n_224
rlabel m2contact 10929 6989 10929 6989 4 n_313
rlabel m2contact 10905 4949 10905 4949 4 n_172
rlabel m2contact 10881 4037 10881 4037 4 n_138
rlabel m2contact 10881 5621 10881 5621 4 n_46
rlabel m2contact 10857 5957 10857 5957 4 n_45
rlabel m2contact 10833 5981 10833 5981 4 stateSub[2]
rlabel m2contact 10761 2909 10761 2909 4 n_34
rlabel m2contact 10761 3005 10761 3005 4 n_325
rlabel m2contact 10713 7373 10713 7373 4 n_310
rlabel m2contact 10713 4037 10713 4037 4 ENB
rlabel m2contact 10689 6437 10689 6437 4 n_272
rlabel m2contact 10665 7277 10665 7277 4 n_39
rlabel m2contact 10665 3917 10665 3917 4 n_273
rlabel m2contact 10641 2909 10641 2909 4 n_494
rlabel m2contact 10617 4085 10617 4085 4 StatusReg[3]
rlabel m2contact 10593 2597 10593 2597 4 n_303
rlabel m2contact 10569 7349 10569 7349 4 n_374
rlabel m2contact 10569 4349 10569 4349 4 n_281
rlabel m2contact 10545 7325 10545 7325 4 n_339
rlabel m2contact 10545 4517 10545 4517 4 n_251
rlabel m2contact 10521 3893 10521 3893 4 n_352
rlabel m2contact 10497 7013 10497 7013 4 n_315
rlabel m2contact 10497 4085 10497 4085 4 nWE
rlabel m2contact 10473 4205 10473 4205 4 n_256
rlabel m2contact 10449 6437 10449 6437 4 n_272
rlabel m2contact 10425 5045 10425 5045 4 n_266
rlabel m2contact 10401 6437 10401 6437 4 n_236
rlabel m2contact 10377 3893 10377 3893 4 n_190
rlabel m2contact 10377 3317 10377 3317 4 n_190
rlabel m2contact 10353 5501 10353 5501 4 n_221
rlabel m2contact 10329 3317 10329 3317 4 n_190
rlabel m2contact 10329 3389 10329 3389 4 n_332
rlabel m2contact 10305 7013 10305 7013 4 n_387
rlabel m2contact 10281 7301 10281 7301 4 n_83
rlabel m2contact 10281 4613 10281 4613 4 n_197
rlabel m2contact 10257 3317 10257 3317 4 n_53
rlabel m2contact 10233 4469 10233 4469 4 n_136
rlabel m2contact 10209 5309 10209 5309 4 n_156
rlabel m2contact 10185 4925 10185 4925 4 n_129
rlabel m2contact 10161 2165 10161 2165 4 n_134
rlabel m2contact 10161 5309 10161 5309 4 n_156
rlabel m2contact 10161 4205 10161 4205 4 n_156
rlabel m2contact 10137 4205 10137 4205 4 n_156
rlabel m2contact 10137 4709 10137 4709 4 n_29
rlabel m2contact 10113 5093 10113 5093 4 n_228
rlabel m2contact 10089 4205 10089 4205 4 n_62
rlabel m2contact 10065 7253 10065 7253 4 n_75
rlabel m2contact 10041 2189 10041 2189 4 n_104
rlabel m2contact 10041 4997 10041 4997 4 n_40
rlabel m2contact 10017 7277 10017 7277 4 n_39
rlabel m2contact 10017 5285 10017 5285 4 n_225
rlabel m2contact 9993 7253 9993 7253 4 n_171
rlabel m2contact 9993 2741 9993 2741 4 n_171
rlabel m2contact 9969 4997 9969 4997 4 n_169
rlabel m2contact 9969 3701 9969 3701 4 n_63
rlabel m2contact 9945 7253 9945 7253 4 n_171
rlabel m2contact 9945 5501 9945 5501 4 n_221
rlabel m2contact 9921 7229 9921 7229 4 n_98
rlabel m2contact 9921 3293 9921 3293 4 n_99
rlabel m2contact 9873 2213 9873 2213 4 n_14
rlabel m2contact 9873 7205 9873 7205 4 n_65
rlabel m2contact 9849 7181 9849 7181 4 n_6
rlabel m2contact 9825 7157 9825 7157 4 n_33
rlabel m2contact 9825 4469 9825 4469 4 n_136
rlabel m2contact 9801 3869 9801 3869 4 stateSub[0]
rlabel m2contact 9753 6701 9753 6701 4 n_90
rlabel m2contact 9705 2237 9705 2237 4 n_20
rlabel m2contact 9705 5933 9705 5933 4 n_22
rlabel m2contact 9657 2957 9657 2957 4 n_160
rlabel m2contact 9633 2261 9633 2261 4 n_21
rlabel m2contact 9633 4877 9633 4877 4 n_356
rlabel m2contact 9609 3341 9609 3341 4 IntReq
rlabel m2contact 9609 2957 9609 2957 4 n_4
rlabel m2contact 9585 4373 9585 4373 4 n_229
rlabel m2contact 9561 6413 9561 6413 4 n_237
rlabel m2contact 9537 4613 9537 4613 4 n_197
rlabel m2contact 9513 2357 9513 2357 4 n_316
rlabel m2contact 9513 4781 9513 4781 4 n_258
rlabel m2contact 9489 4877 9489 4877 4 n_275
rlabel m2contact 9489 3797 9489 3797 4 n_275
rlabel m2contact 9465 7133 9465 7133 4 n_198
rlabel m2contact 9465 7037 9465 7037 4 n_349
rlabel m2contact 9441 7061 9441 7061 4 n_47
rlabel m2contact 9417 6917 9417 6917 4 n_231
rlabel m2contact 9393 4877 9393 4877 4 n_275
rlabel m2contact 9393 4469 9393 4469 4 n_136
rlabel m2contact 9369 4613 9369 4613 4 n_197
rlabel m2contact 9345 5645 9345 5645 4 OpcodeCondIn[6]
rlabel m2contact 9321 2357 9321 2357 4 n_133
rlabel m2contact 9297 2285 9297 2285 4 n_176
rlabel m2contact 9297 4901 9297 4901 4 n_157
rlabel m2contact 9273 2357 9273 2357 4 n_133
rlabel m2contact 9273 2477 9273 2477 4 n_132
rlabel m2contact 9249 4061 9249 4061 4 n_175
rlabel m2contact 9225 2357 9225 2357 4 AluEn
rlabel m2contact 9201 5093 9201 5093 4 n_228
rlabel m2contact 9201 2285 9201 2285 4 n_228
rlabel m2contact 9177 2285 9177 2285 4 n_228
rlabel m2contact 9177 4877 9177 4877 4 n_377
rlabel m2contact 9153 3797 9153 3797 4 n_275
rlabel m2contact 9129 6701 9129 6701 4 n_90
rlabel m2contact 9105 7109 9105 7109 4 n_27
rlabel m2contact 9093 7061 9093 7061 4 n_303
rlabel m2contact 9093 2597 9093 2597 4 n_303
rlabel m2contact 9081 2357 9081 2357 4 AluEn
rlabel m2contact 9057 7085 9057 7085 4 n_70
rlabel m2contact 9057 4877 9057 4877 4 n_377
rlabel m2contact 9033 6797 9033 6797 4 n_359
rlabel m2contact 9009 3005 9009 3005 4 n_325
rlabel m2contact 9009 3485 9009 3485 4 OpcodeCondIn[1]
rlabel m2contact 8985 7061 8985 7061 4 n_303
rlabel m2contact 8985 6077 8985 6077 4 n_299
rlabel m2contact 8937 6533 8937 6533 4 n_26
rlabel m2contact 8913 3101 8913 3101 4 stateSub[1]
rlabel m2contact 8889 3797 8889 3797 4 n_275
rlabel m2contact 8841 3341 8841 3341 4 IntReq
rlabel m2contact 8841 3533 8841 3533 4 n_246
rlabel m2contact 8817 4781 8817 4781 4 n_258
rlabel m2contact 8793 5477 8793 5477 4 n_200
rlabel m2contact 8745 3533 8745 3533 4 ImmSel
rlabel m2contact 8697 4229 8697 4229 4 n_111
rlabel m2contact 8673 5837 8673 5837 4 n_96
rlabel m2contact 8649 5093 8649 5093 4 n_228
rlabel m2contact 8625 3845 8625 3845 4 n_110
rlabel m2contact 8577 4733 8577 4733 4 n_328
rlabel m2contact 8553 3101 8553 3101 4 stateSub[1]
rlabel m2contact 8529 3341 8529 3341 4 n_294
rlabel m2contact 8481 4733 8481 4733 4 n_347
rlabel m2contact 8457 4229 8457 4229 4 Flags[3]
rlabel m2contact 8433 7037 8433 7037 4 n_349
rlabel m2contact 8385 2357 8385 2357 4 n_168
rlabel m2contact 8361 3005 8361 3005 4 n_125
rlabel m2contact 8337 3869 8337 3869 4 stateSub[0]
rlabel m2contact 8313 7037 8313 7037 4 n_335
rlabel m2contact 8313 2525 8313 2525 4 n_335
rlabel m2contact 8289 7037 8289 7037 4 n_335
rlabel m2contact 8289 5117 8289 5117 4 n_84
rlabel m2contact 8265 6917 8265 6917 4 n_231
rlabel m2contact 8265 3221 8265 3221 4 n_92
rlabel m2contact 8241 4541 8241 4541 4 n_244
rlabel m2contact 8217 7013 8217 7013 4 n_387
rlabel m2contact 8193 6989 8193 6989 4 n_313
rlabel m2contact 8169 2309 8169 2309 4 n_124
rlabel m2contact 8169 6965 8169 6965 4 n_170
rlabel m2contact 8145 2333 8145 2333 4 n_379
rlabel m2contact 8145 6941 8145 6941 4 n_202
rlabel m2contact 8121 6917 8121 6917 4 n_231
rlabel m2contact 8097 6893 8097 6893 4 n_115
rlabel m2contact 8049 2357 8049 2357 4 n_168
rlabel m2contact 8049 2381 8049 2381 4 n_223
rlabel m2contact 8025 3293 8025 3293 4 n_99
rlabel m2contact 8001 2405 8001 2405 4 n_149
rlabel m2contact 8001 6869 8001 6869 4 n_216
rlabel m2contact 7977 5501 7977 5501 4 n_221
rlabel m2contact 7953 2429 7953 2429 4 n_100
rlabel m2contact 7953 3893 7953 3893 4 n_190
rlabel m2contact 7905 5645 7905 5645 4 OpcodeCondIn[6]
rlabel m2contact 7905 3893 7905 3893 4 n_73
rlabel m2contact 7881 6845 7881 6845 4 n_189
rlabel m2contact 7881 6701 7881 6701 4 n_90
rlabel m2contact 7857 5045 7857 5045 4 n_266
rlabel m2contact 7809 2453 7809 2453 4 n_9
rlabel m2contact 7809 6821 7809 6821 4 n_363
rlabel m2contact 7785 6797 7785 6797 4 n_359
rlabel m2contact 7785 3869 7785 3869 4 stateSub[0]
rlabel m2contact 7761 6773 7761 6773 4 n_298
rlabel m2contact 7761 3749 7761 3749 4 state[0]
rlabel m2contact 7713 2477 7713 2477 4 n_132
rlabel m2contact 7713 6749 7713 6749 4 n_74
rlabel m2contact 7689 5381 7689 5381 4 n_80
rlabel m2contact 7665 6701 7665 6701 4 n_90
rlabel m2contact 7641 2573 7641 2573 4 n_11
rlabel m2contact 7617 6725 7617 6725 4 n_239
rlabel m2contact 7617 6701 7617 6701 4 n_275
rlabel m2contact 7617 3797 7617 3797 4 n_275
rlabel m2contact 7593 6701 7593 6701 4 n_275
rlabel m2contact 7593 4109 7593 4109 4 n_56
rlabel m2contact 7569 4637 7569 4637 4 n_232
rlabel m2contact 7545 6461 7545 6461 4 n_185
rlabel m2contact 7521 5837 7521 5837 4 n_96
rlabel m2contact 7497 6677 7497 6677 4 n_13
rlabel m2contact 7473 2501 7473 2501 4 AluOR[1]
rlabel m2contact 7449 2621 7449 2621 4 n_306
rlabel m2contact 7449 3461 7449 3461 4 n_122
rlabel m2contact 7425 5453 7425 5453 4 n_284
rlabel m2contact 7401 2525 7401 2525 4 n_335
rlabel m2contact 7401 3965 7401 3965 4 n_351
rlabel m2contact 7377 6653 7377 6653 4 n_163
rlabel m2contact 7353 6629 7353 6629 4 n_249
rlabel m2contact 7353 3965 7353 3965 4 nME
rlabel m2contact 7329 6605 7329 6605 4 n_184
rlabel m2contact 7305 6581 7305 6581 4 n_268
rlabel m2contact 7281 6557 7281 6557 4 n_120
rlabel m2contact 7257 5549 7257 5549 4 n_86
rlabel m2contact 7233 5045 7233 5045 4 n_266
rlabel m2contact 7185 6533 7185 6533 4 n_26
rlabel m2contact 7161 3197 7161 3197 4 n_187
rlabel m2contact 7137 2549 7137 2549 4 Op2Sel[0]
rlabel m2contact 7089 2573 7089 2573 4 n_11
rlabel m2contact 7065 2621 7065 2621 4 n_306
rlabel m2contact 7041 6509 7041 6509 4 n_353
rlabel m2contact 7041 4685 7041 4685 4 OpcodeCondIn[3]
rlabel m2contact 7017 4853 7017 4853 4 n_381
rlabel m2contact 6993 6485 6993 6485 4 n_205
rlabel m2contact 6993 6053 6993 6053 4 n_177
rlabel m2contact 6969 2597 6969 2597 4 n_303
rlabel m2contact 6945 2621 6945 2621 4 RwSel[0]
rlabel m2contact 6897 2741 6897 2741 4 n_171
rlabel m2contact 6849 6461 6849 6461 4 n_185
rlabel m2contact 6825 4901 6825 4901 4 n_157
rlabel m2contact 6777 2621 6777 2621 4 RwSel[0]
rlabel m2contact 6777 6437 6777 6437 4 n_236
rlabel m2contact 6753 6149 6753 6149 4 n_253
rlabel m2contact 6729 5261 6729 5261 4 n_173
rlabel m2contact 6705 4493 6705 4493 4 n_161
rlabel m2contact 6681 5261 6681 5261 4 n_254
rlabel m2contact 6681 3389 6681 3389 4 n_332
rlabel m2contact 6657 6413 6657 6413 4 n_237
rlabel m2contact 6633 6149 6633 6149 4 n_253
rlabel m2contact 6609 2645 6609 2645 4 n_196
rlabel m2contact 6609 6389 6609 6389 4 n_17
rlabel m2contact 6537 6365 6537 6365 4 SysBus[0]
rlabel m2contact 6489 3845 6489 3845 4 n_110
rlabel m2contact 6465 6341 6465 6341 4 n_224
rlabel m2contact 6465 5045 6465 5045 4 n_266
rlabel m2contact 6441 5117 6441 5117 4 n_84
rlabel m2contact 6393 6317 6393 6317 4 StatusReg[0]
rlabel m2contact 6393 4013 6393 4013 4 n_60
rlabel m2contact 6345 2669 6345 2669 4 n_101
rlabel m2contact 6321 6293 6321 6293 4 IRQ2
rlabel m2contact 6321 3293 6321 3293 4 n_99
rlabel m2contact 6297 4253 6297 4253 4 n_495
rlabel m2contact 6249 4589 6249 4589 4 n_174
rlabel m2contact 6249 4253 6249 4253 4 nWait
rlabel m2contact 6225 2693 6225 2693 4 n_270
rlabel m2contact 6201 3845 6201 3845 4 n_110
rlabel m2contact 6177 2717 6177 2717 4 n_240
rlabel m2contact 6177 4517 6177 4517 4 n_251
rlabel m2contact 6129 2741 6129 2741 4 n_171
rlabel m2contact 6129 6269 6129 6269 4 n_346
rlabel m2contact 6105 6245 6105 6245 4 n_345
rlabel m2contact 6105 4517 6105 4517 4 n_251
rlabel m2contact 6081 2765 6081 2765 4 InISR
rlabel m2contact 6057 3533 6057 3533 4 ImmSel
rlabel m2contact 6033 2789 6033 2789 4 n_279
rlabel m2contact 6033 6221 6033 6221 4 n_58
rlabel m2contact 6009 3533 6009 3533 4 n_354
rlabel m2contact 6009 3845 6009 3845 4 n_110
rlabel m2contact 5985 2813 5985 2813 4 n_296
rlabel m2contact 5985 4829 5985 4829 4 n_50
rlabel m2contact 5913 3149 5913 3149 4 n_384
rlabel m2contact 5913 4901 5913 4901 4 n_157
rlabel m2contact 5889 4661 5889 4661 4 OpcodeCondIn[7]
rlabel m2contact 5865 6197 5865 6197 4 n_105
rlabel m2contact 5865 5285 5865 5285 4 n_225
rlabel m2contact 5841 4469 5841 4469 4 n_136
rlabel m2contact 5817 6173 5817 6173 4 n_277
rlabel m2contact 5793 4829 5793 4829 4 n_243
rlabel m2contact 5769 6149 5769 6149 4 n_253
rlabel m2contact 5769 3461 5769 3461 4 n_122
rlabel m2contact 5745 3797 5745 3797 4 n_275
rlabel m2contact 5721 6125 5721 6125 4 n_259
rlabel m2contact 5721 5813 5721 5813 4 n_203
rlabel m2contact 5697 4805 5697 4805 4 n_255
rlabel m2contact 5673 2837 5673 2837 4 n_79
rlabel m2contact 5673 6101 5673 6101 4 n_257
rlabel m2contact 5649 4781 5649 4781 4 n_258
rlabel m2contact 5649 4157 5649 4157 4 n_78
rlabel m2contact 5625 5045 5625 5045 4 n_266
rlabel m2contact 5577 6029 5577 6029 4 n_291
rlabel m2contact 5529 2861 5529 2861 4 n_207
rlabel m2contact 5481 2885 5481 2885 4 StatusReg[2]
rlabel m2contact 5481 6077 5481 6077 4 n_299
rlabel m2contact 5457 6053 5457 6053 4 n_177
rlabel m2contact 5433 2909 5433 2909 4 n_494
rlabel m2contact 5433 6029 5433 6029 4 n_291
rlabel m2contact 5385 6005 5385 6005 4 n_68
rlabel m2contact 5361 5741 5361 5741 4 OpcodeCondIn[2]
rlabel m2contact 5337 5981 5337 5981 4 stateSub[2]
rlabel m2contact 5313 5957 5313 5957 4 n_45
rlabel m2contact 5289 5501 5289 5501 4 n_221
rlabel m2contact 5241 5933 5241 5933 4 n_22
rlabel m2contact 5217 5837 5217 5837 4 n_96
rlabel m2contact 5193 3557 5193 3557 4 state[1]
rlabel m2contact 5145 5909 5145 5909 4 n_24
rlabel m2contact 5121 3485 5121 3485 4 OpcodeCondIn[1]
rlabel m2contact 5097 5885 5097 5885 4 n_19
rlabel m2contact 5073 5861 5073 5861 4 n_372
rlabel m2contact 5049 2933 5049 2933 4 n_97
rlabel m2contact 5025 5837 5025 5837 4 n_96
rlabel m2contact 5001 3221 5001 3221 4 n_92
rlabel m2contact 4929 5813 4929 5813 4 n_203
rlabel m2contact 4905 4133 4905 4133 4 n_183
rlabel m2contact 4881 5789 4881 5789 4 n_15
rlabel m2contact 4857 5765 4857 5765 4 n_61
rlabel m2contact 4809 2957 4809 2957 4 n_4
rlabel m2contact 4785 4013 4785 4013 4 n_60
rlabel m2contact 4761 4253 4761 4253 4 nWait
rlabel m2contact 4713 4013 4713 4013 4 n_57
rlabel m2contact 4689 2981 4689 2981 4 WdSel
rlabel m2contact 4689 5741 4689 5741 4 OpcodeCondIn[2]
rlabel m2contact 4665 5717 4665 5717 4 n_496
rlabel m2contact 4641 5693 4641 5693 4 n_158
rlabel m2contact 4593 4061 4593 4061 4 n_175
rlabel m2contact 4569 5669 4569 5669 4 OpcodeCondIn[4]
rlabel m2contact 4545 5501 4545 5501 4 n_221
rlabel m2contact 4545 4061 4545 4061 4 nIRQ
rlabel m2contact 4521 4925 4521 4925 4 n_129
rlabel m2contact 4497 3005 4497 3005 4 n_125
rlabel m2contact 4497 5645 4497 5645 4 OpcodeCondIn[6]
rlabel m2contact 4473 5501 4473 5501 4 n_221
rlabel m2contact 4449 3029 4449 3029 4 n_71
rlabel m2contact 4449 3053 4449 3053 4 n_233
rlabel m2contact 4425 5621 4425 5621 4 n_46
rlabel m2contact 4401 3077 4401 3077 4 n_154
rlabel m2contact 4377 5597 4377 5597 4 n_164
rlabel m2contact 4353 3101 4353 3101 4 stateSub[1]
rlabel m2contact 4353 3125 4353 3125 4 n_121
rlabel m2contact 4305 5573 4305 5573 4 n_87
rlabel m2contact 4281 3845 4281 3845 4 n_110
rlabel m2contact 4257 5549 4257 5549 4 n_86
rlabel m2contact 4257 4973 4257 4973 4 n_219
rlabel m2contact 4209 3149 4209 3149 4 n_384
rlabel m2contact 4209 5525 4209 5525 4 n_222
rlabel m2contact 4185 5501 4185 5501 4 n_221
rlabel m2contact 4161 3173 4161 3173 4 n_211
rlabel m2contact 4161 4973 4161 4973 4 n_219
rlabel m2contact 4137 4709 4137 4709 4 n_29
rlabel m2contact 4113 3197 4113 3197 4 n_187
rlabel m2contact 4089 4973 4089 4973 4 n_201
rlabel m2contact 4041 5477 4041 5477 4 n_200
rlabel m2contact 4017 3221 4017 3221 4 n_92
rlabel m2contact 3993 5453 3993 5453 4 n_284
rlabel m2contact 3969 3245 3969 3245 4 n_143
rlabel m2contact 3969 5429 3969 5429 4 n_227
rlabel m2contact 3945 5285 3945 5285 4 n_225
rlabel m2contact 3921 3269 3921 3269 4 n_206
rlabel m2contact 3921 5189 3921 5189 4 n_226
rlabel m2contact 3897 3293 3897 3293 4 n_99
rlabel m2contact 3873 5405 3873 5405 4 n_51
rlabel m2contact 3849 3317 3849 3317 4 n_53
rlabel m2contact 3849 5381 3849 5381 4 n_80
rlabel m2contact 3825 5357 3825 5357 4 n_287
rlabel m2contact 3801 4109 3801 4109 4 n_56
rlabel m2contact 3777 5333 3777 5333 4 n_142
rlabel m2contact 3753 5309 3753 5309 4 n_156
rlabel m2contact 3729 5285 3729 5285 4 n_225
rlabel m2contact 3729 3797 3729 3797 4 n_275
rlabel m2contact 3705 5261 3705 5261 4 n_254
rlabel m2contact 3681 5237 3681 5237 4 n_151
rlabel m2contact 3657 3341 3657 3341 4 n_294
rlabel m2contact 3657 4661 3657 4661 4 OpcodeCondIn[7]
rlabel m2contact 3633 5213 3633 5213 4 n_128
rlabel m2contact 3633 3869 3633 3869 4 stateSub[0]
rlabel m2contact 3609 3365 3609 3365 4 n_293
rlabel m2contact 3585 3389 3585 3389 4 n_332
rlabel m2contact 3585 3413 3585 3413 4 n_210
rlabel m2contact 3561 5189 3561 5189 4 n_226
rlabel m2contact 3537 3437 3537 3437 4 n_119
rlabel m2contact 3537 5165 3537 5165 4 n_260
rlabel m2contact 3489 5141 3489 5141 4 n_77
rlabel m2contact 3489 4493 3489 4493 4 n_161
rlabel m2contact 3465 5117 3465 5117 4 n_84
rlabel m2contact 3441 3461 3441 3461 4 n_122
rlabel m2contact 3441 5093 3441 5093 4 n_228
rlabel m2contact 3393 3485 3393 3485 4 OpcodeCondIn[1]
rlabel m2contact 3393 5069 3393 5069 4 n_247
rlabel m2contact 3345 3509 3345 3509 4 n_117
rlabel m2contact 3321 4109 3321 4109 4 n_56
rlabel m2contact 3249 3533 3249 3533 4 n_354
rlabel m2contact 3225 3557 3225 3557 4 state[1]
rlabel m2contact 3201 3581 3201 3581 4 n_326
rlabel m2contact 3177 4781 3177 4781 4 n_258
rlabel m2contact 3153 3605 3153 3605 4 n_94
rlabel m2contact 3129 5045 3129 5045 4 n_266
rlabel m2contact 3105 4589 3105 4589 4 n_174
rlabel m2contact 3057 5021 3057 5021 4 n_264
rlabel m2contact 3033 4997 3033 4997 4 n_169
rlabel m2contact 3009 4973 3009 4973 4 n_201
rlabel m2contact 2961 4949 2961 4949 4 n_172
rlabel m2contact 2937 4925 2937 4925 4 n_129
rlabel m2contact 2913 4901 2913 4901 4 n_157
rlabel m2contact 2841 4877 2841 4877 4 n_377
rlabel m2contact 2817 3629 2817 3629 4 n_362
rlabel m2contact 2793 4853 2793 4853 4 n_381
rlabel m2contact 2745 4829 2745 4829 4 n_243
rlabel m2contact 2721 4805 2721 4805 4 n_255
rlabel m2contact 2697 4781 2697 4781 4 n_258
rlabel m2contact 2649 4757 2649 4757 4 n_371
rlabel m2contact 2625 3653 2625 3653 4 n_329
rlabel m2contact 2601 3677 2601 3677 4 n_64
rlabel m2contact 2601 4733 2601 4733 4 n_347
rlabel m2contact 2577 3701 2577 3701 4 n_63
rlabel m2contact 2577 3725 2577 3725 4 n_311
rlabel m2contact 2553 3797 2553 3797 4 n_275
rlabel m2contact 2529 3749 2529 3749 4 state[0]
rlabel m2contact 2529 4709 2529 4709 4 n_29
rlabel m2contact 2505 4685 2505 4685 4 OpcodeCondIn[3]
rlabel m2contact 2481 3773 2481 3773 4 n_276
rlabel m2contact 2481 4661 2481 4661 4 OpcodeCondIn[7]
rlabel m2contact 2457 3797 2457 3797 4 n_275
rlabel m2contact 2433 3821 2433 3821 4 n_267
rlabel m2contact 2433 4637 2433 4637 4 n_232
rlabel m2contact 2385 4613 2385 4613 4 n_197
rlabel m2contact 2361 4589 2361 4589 4 n_174
rlabel m2contact 2313 4565 2313 4565 4 n_252
rlabel m2contact 2289 3845 2289 3845 4 n_110
rlabel m2contact 2289 3869 2289 3869 4 stateSub[0]
rlabel m2contact 2265 4541 2265 4541 4 n_244
rlabel m2contact 2241 3869 2241 3869 4 stateSub[0]
rlabel m2contact 2241 4517 2241 4517 4 n_251
rlabel m2contact 2193 4493 2193 4493 4 n_161
rlabel m2contact 2169 4469 2169 4469 4 n_136
rlabel m2contact 2145 4109 2145 4109 4 n_56
rlabel m2contact 2097 4109 2097 4109 4 nOE
rlabel m2contact 2073 3893 2073 3893 4 n_73
rlabel m2contact 2049 4445 2049 4445 4 n_324
rlabel m2contact 2025 4421 2025 4421 4 n_366
rlabel m2contact 2001 4397 2001 4397 4 n_241
rlabel m2contact 1953 3917 1953 3917 4 n_273
rlabel m2contact 1929 4373 1929 4373 4 n_229
rlabel m2contact 1905 4349 1905 4349 4 n_281
rlabel m2contact 1881 4325 1881 4325 4 n_139
rlabel m2contact 1857 3941 1857 3941 4 n_321
rlabel m2contact 1833 4301 1833 4301 4 n_265
rlabel m2contact 1809 4277 1809 4277 4 n_214
rlabel m2contact 1761 4253 1761 4253 4 nWait
rlabel m2contact 1761 4229 1761 4229 4 Flags[3]
rlabel m2contact 1713 3965 1713 3965 4 nME
rlabel m2contact 1689 4205 1689 4205 4 n_62
rlabel m2contact 1665 3989 1665 3989 4 n_147
rlabel m2contact 1665 4181 1665 4181 4 n_182
rlabel m2contact 1641 4157 1641 4157 4 n_78
rlabel m2contact 1617 4013 1617 4013 4 n_57
rlabel m2contact 1617 4133 1617 4133 4 n_183
rlabel metal2 26271 8799 26283 8799 6 MemEn
rlabel metal2 24735 8799 24747 8799 6 IrWe
rlabel metal2 23199 8799 23211 8799 6 LrSel
rlabel metal2 21663 8799 21675 8799 6 LrWe
rlabel metal2 20127 8799 20139 8799 6 WdSel
rlabel metal2 20103 8799 20115 8799 6 LrEn
rlabel metal2 17055 8799 17067 8799 6 PcSel[0]
rlabel metal2 17031 8799 17043 8799 6 PcSel[1]
rlabel metal2 15495 8799 15507 8799 6 PcSel[2]
rlabel metal2 13947 8799 13959 8799 4 PcEn
rlabel metal2 12255 8799 12267 8799 4 PcWe
rlabel metal2 10851 8799 10863 8799 4 Op1Sel
rlabel metal2 8751 8799 8763 8799 4 ImmSel
rlabel metal2 7143 8799 7155 8799 4 Op2Sel[0]
rlabel metal2 4695 8799 4707 8799 4 Op2Sel[1]
rlabel metal2 4659 8799 4671 8799 4 AluWe
rlabel metal2 3111 8799 3123 8799 4 AluEn
rlabel metal2 28311 8584 28311 8596 6 CFlag
rlabel metal2 28311 8560 28311 8572 6 RegWe
rlabel metal2 28311 8536 28311 8548 6 RwSel[0]
rlabel metal2 28311 8512 28311 8524 6 Rs1Sel[1]
rlabel metal2 28311 8488 28311 8500 6 RwSel[1]
rlabel metal2 28311 8464 28311 8476 6 Rs1Sel[0]
rlabel metal2 28311 8440 28311 8452 6 AluOR[0]
rlabel metal2 28311 126 28311 138 8 OpcodeCondIn[0]
rlabel metal2 28311 102 28311 114 8 OpcodeCondIn[2]
rlabel metal2 28311 78 28311 90 8 OpcodeCondIn[7]
rlabel metal2 28311 54 28311 66 8 OpcodeCondIn[6]
rlabel metal2 28311 30 28311 42 8 OpcodeCondIn[4]
rlabel metal2 28311 6 28311 18 8 OpcodeCondIn[5]
rlabel metal2 28311 2495 28311 2507 6 AluOR[1]
rlabel metal2 28311 2063 28311 2075 6 SysBus[1]
rlabel metal2 28311 2039 28311 2051 6 SysBus[0]
rlabel metal2 28311 2015 28311 2027 6 SysBus[3]
rlabel metal2 28311 1991 28311 2003 6 SysBus[2]
rlabel metal2 28311 1967 28311 1979 6 OpcodeCondIn[3]
rlabel metal2 28311 1943 28311 1955 6 OpcodeCondIn[1]
rlabel metal2 27915 8799 28115 8799 5 GND!
rlabel metal2 27915 0 28115 0 1 GND!
rlabel metal2 0 78 0 90 2 Flags[1]
rlabel metal2 0 54 0 66 2 Flags[3]
rlabel metal2 0 30 0 42 2 Flags[2]
rlabel metal2 0 6 0 18 2 Flags[0]
rlabel metal2 0 4103 0 4115 4 nOE
rlabel metal2 0 4079 0 4091 4 nWE
rlabel metal2 0 4055 0 4067 4 nIRQ
rlabel metal2 0 4031 0 4043 4 ENB
rlabel metal2 0 8632 0 8644 4 ALE
rlabel metal2 0 8608 0 8620 4 nME
rlabel metal2 0 8584 0 8596 4 nWait
rlabel metal2 123 0 323 0 1 Vdd!
rlabel metal2 123 8799 323 8799 5 Vdd!
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 339 8799 351 8799 5 SDO
rlabel metal2 387 8799 399 8799 5 Clock
rlabel metal2 363 8799 375 8799 5 Test
rlabel metal2 411 8799 423 8799 5 nReset
<< end >>
