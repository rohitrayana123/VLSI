../../../Design/Implementation/verilog/behavioural/trisBuf16.sv