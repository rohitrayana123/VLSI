magic
tech c035u
timestamp 1394314552
<< metal1 >>
rect 1573 1062 3023 1072
rect 3037 1062 12360 1072
rect 0 95 2903 105
rect 2917 95 3071 105
rect 3085 95 12364 105
rect 0 73 12364 83
rect 2629 51 12364 61
rect 12109 29 12364 39
rect 12325 7 12364 17
<< m2contact >>
rect 1559 1060 1573 1074
rect 3023 1060 3037 1074
rect 2903 93 2917 107
rect 3071 93 3085 107
rect 2615 49 2629 63
rect 12095 27 12109 41
rect 12311 5 12325 19
<< metal2 >>
rect 216 1050 228 1079
rect 360 1050 372 1079
rect 576 1050 588 1079
rect 1320 1050 1332 1079
rect 1488 1050 1500 1079
rect 1560 1050 1572 1060
rect 1872 1050 1884 1079
rect 2088 1050 2100 1079
rect 2832 1050 2844 1079
rect 3000 970 3012 1079
rect 3024 970 3036 1060
rect 3096 1050 3180 1062
rect 3216 1050 3228 1079
rect 3960 1050 3972 1079
rect 4176 1050 4188 1079
rect 4368 1050 4380 1079
rect 5112 1050 5124 1079
rect 5328 1050 5340 1079
rect 5520 1050 5532 1079
rect 6264 1050 6276 1079
rect 6480 1050 6492 1079
rect 6672 1050 6684 1079
rect 7416 1050 7428 1079
rect 7632 1050 7644 1079
rect 7824 1050 7836 1079
rect 8568 1050 8580 1079
rect 8784 1050 8796 1079
rect 8976 1050 8988 1079
rect 9720 1050 9732 1079
rect 9936 1050 9948 1079
rect 10128 1050 10140 1079
rect 10872 1050 10884 1079
rect 11088 1050 11100 1079
rect 11280 1050 11292 1079
rect 12024 1050 12036 1079
rect 12240 1050 12252 1079
rect 3096 970 3108 1050
rect 216 0 228 111
rect 360 0 372 111
rect 576 0 588 111
rect 1320 0 1332 111
rect 1488 0 1500 111
rect 1872 0 1884 111
rect 2088 0 2100 111
rect 2616 63 2628 111
rect 2832 0 2844 111
rect 2904 107 2916 111
rect 3000 0 3012 171
rect 3072 107 3084 171
rect 3216 0 3228 111
rect 3960 0 3972 111
rect 4176 0 4188 111
rect 4368 0 4380 111
rect 5112 0 5124 111
rect 5328 0 5340 111
rect 5520 0 5532 111
rect 6264 0 6276 111
rect 6480 0 6492 111
rect 6672 0 6684 111
rect 7416 0 7428 111
rect 7632 0 7644 111
rect 7824 0 7836 111
rect 8568 0 8580 111
rect 8784 0 8796 111
rect 8976 0 8988 111
rect 9720 0 9732 111
rect 9936 0 9948 111
rect 10128 0 10140 111
rect 10872 0 10884 111
rect 11088 0 11100 111
rect 11280 0 11292 111
rect 12024 0 12036 111
rect 12096 41 12108 111
rect 12240 0 12252 111
rect 12312 19 12324 111
use Pc_slice Pc_slice_0
timestamp 1394294966
transform 1 0 0 0 1 111
box 0 0 2952 939
use mux2 mux2_0
timestamp 1386235218
transform 1 0 2952 0 1 171
box 0 0 192 799
use regBlock_slice regBlock_slice_0
timestamp 1394295027
transform 1 0 3144 0 1 111
box 0 0 9216 939
<< labels >>
rlabel metal1 3096 100 3096 100 1 SysBus
rlabel metal1 12358 1067 12358 1067 6 AluOut
rlabel metal1 12353 34 12353 34 1 Rd1
rlabel metal1 12355 11 12355 11 1 Rd2
rlabel metal2 216 0 228 0 1 PcIncCin
rlabel metal2 360 0 372 0 1 LrSel
rlabel metal2 576 0 588 0 1 LrWe
rlabel metal2 1320 0 1332 0 1 LrEn
rlabel metal2 1488 0 1500 0 1 PcSel[0]
rlabel metal2 1872 0 1884 0 1 PcSel[1]
rlabel metal2 2088 0 2100 0 1 PcWe
rlabel metal2 2832 0 2844 0 1 PcEn
rlabel metal2 3000 0 3012 0 1 WdSel
rlabel metal2 3960 0 3972 0 1 Rs1[0]
rlabel metal2 4368 0 4380 0 1 Rw[1]
rlabel metal2 5112 0 5124 0 1 Rs1[1]
rlabel metal2 5328 0 5340 0 1 Rs2[1]
rlabel metal2 5520 0 5532 0 1 Rw[2]
rlabel metal2 6264 0 6276 0 1 Rs1[2]
rlabel metal2 6480 0 6492 0 1 Rs2[2]
rlabel metal2 6672 0 6684 0 1 Rw[3]
rlabel metal2 7416 0 7428 0 1 Rs1[3]
rlabel metal2 7632 0 7644 0 1 Rs2[3]
rlabel metal2 7824 0 7836 0 1 Rw[4]
rlabel metal2 8568 0 8580 0 1 Rs1[4]
rlabel metal2 8784 0 8796 0 1 Rs2[4]
rlabel metal2 8976 0 8988 0 1 Rw[5]
rlabel metal2 9720 0 9732 0 1 Rs1[5]
rlabel metal2 9936 0 9948 0 1 Rs2[5]
rlabel metal2 10128 0 10140 0 1 Rw[6]
rlabel metal2 10872 0 10884 0 1 Rs1[6]
rlabel metal2 11088 0 11100 0 1 Rs2[6]
rlabel metal2 11280 0 11292 0 1 Rw[7]
rlabel metal2 12024 0 12036 0 1 Rs1[7]
rlabel metal2 12240 0 12252 0 1 Rs2[7]
rlabel metal1 12352 100 12352 100 1 SysBus
rlabel metal1 12353 78 12353 78 1 Imm
rlabel metal1 12354 56 12354 56 1 Pc
rlabel metal2 12240 1079 12252 1079 5 Rs2[7]
rlabel metal2 12024 1079 12036 1079 5 Rs1[7]
rlabel metal2 11280 1079 11292 1079 5 Rw[7]
rlabel metal2 11088 1079 11100 1079 5 Rs2[6]
rlabel metal2 10872 1079 10884 1079 5 Rs1[6]
rlabel metal2 10128 1079 10140 1079 5 Rw[6]
rlabel metal2 9720 1079 9732 1079 5 Rs1[5]
rlabel metal2 9936 1079 9948 1079 5 Rs2[5]
rlabel metal2 8976 1079 8988 1079 5 Rw[5]
rlabel metal2 8784 1079 8796 1079 5 Rs2[4]
rlabel metal2 8568 1079 8580 1079 5 Rs1[4]
rlabel metal2 7824 1079 7836 1079 5 Rw[4]
rlabel metal2 7632 1079 7644 1079 5 Rs2[3]
rlabel metal2 7416 1079 7428 1079 5 Rs1[3]
rlabel metal2 6672 1079 6684 1079 5 Rw[3]
rlabel metal2 6480 1079 6492 1079 5 Rs2[2]
rlabel metal2 6264 1079 6276 1079 5 Rs1[2]
rlabel metal2 5520 1079 5532 1079 5 Rw[2]
rlabel metal2 5328 1079 5340 1079 5 Rs2[1]
rlabel metal2 5112 1079 5124 1079 5 Rs1[1]
rlabel metal2 4368 1079 4380 1079 5 Rw[1]
rlabel metal2 4176 1079 4188 1079 5 Rs2[0]
rlabel metal2 3960 1079 3972 1079 5 Rs1[0]
rlabel metal2 3216 1079 3228 1079 5 Rw[0]
rlabel metal2 3000 1079 3012 1079 5 WdSel
rlabel metal2 2832 1079 2844 1079 5 PcEn
rlabel metal2 2088 1079 2100 1079 5 PcWe
rlabel metal2 1872 1079 1884 1079 5 PcSel[1]
rlabel metal2 1488 1079 1500 1079 5 PcSel[0]
rlabel metal2 1320 1079 1332 1079 5 LrEn
rlabel metal2 576 1079 588 1079 5 LrWe
rlabel metal2 360 1079 372 1079 5 LrSel
rlabel metal2 216 1079 228 1079 5 PcIncCout
rlabel metal2 3216 0 3228 0 1 Rw[0]
rlabel metal2 4176 0 4188 0 1 Rs2[0]
rlabel metal1 0 95 0 105 1 SysBus
rlabel metal1 0 73 0 83 1 Imm
<< end >>
