magic
tech c035u
timestamp 1394475869
<< metal1 >>
rect 1573 1159 3023 1169
rect 3037 1159 12360 1169
rect 0 95 2903 105
rect 2917 95 3071 105
rect 3085 95 12364 105
rect 0 73 12364 83
rect 2629 51 12364 61
rect 12109 29 12364 39
rect 12325 7 12364 17
<< m2contact >>
rect 1559 1157 1573 1171
rect 3023 1157 3037 1171
rect 2903 93 2917 107
rect 3071 93 3085 107
rect 2615 49 2629 63
rect 12095 27 12109 41
rect 12311 5 12325 19
<< metal2 >>
rect 216 1153 228 1176
rect 360 1153 372 1176
rect 576 1153 588 1176
rect 1320 1153 1332 1176
rect 1488 1153 1500 1176
rect 1560 1153 1572 1157
rect 1872 1153 1884 1176
rect 2088 1153 2100 1176
rect 2832 1153 2844 1176
rect 3000 976 3012 1176
rect 3024 976 3036 1157
rect 3096 1153 3180 1165
rect 3216 1153 3228 1176
rect 3960 1153 3972 1176
rect 4176 1153 4188 1176
rect 4368 1153 4380 1176
rect 5112 1153 5124 1176
rect 5328 1153 5340 1176
rect 5520 1153 5532 1176
rect 6264 1153 6276 1176
rect 6480 1153 6492 1176
rect 6672 1153 6684 1176
rect 7416 1153 7428 1176
rect 7632 1153 7644 1176
rect 7824 1153 7836 1176
rect 8568 1153 8580 1176
rect 8784 1153 8796 1176
rect 8976 1153 8988 1176
rect 9720 1153 9732 1176
rect 9936 1153 9948 1176
rect 10128 1153 10140 1176
rect 10872 1153 10884 1176
rect 11088 1153 11100 1176
rect 11280 1153 11292 1176
rect 12024 1153 12036 1176
rect 12240 1153 12252 1176
rect 3096 976 3108 1153
rect 216 0 228 111
rect 360 0 372 111
rect 576 0 588 111
rect 1320 0 1332 111
rect 1488 0 1500 111
rect 1872 0 1884 111
rect 2088 0 2100 111
rect 2616 63 2628 111
rect 2832 0 2844 111
rect 2904 107 2916 111
rect 3000 0 3012 177
rect 3072 107 3084 177
rect 3216 0 3228 111
rect 3960 0 3972 111
rect 4176 0 4188 111
rect 4368 0 4380 111
rect 5112 0 5124 111
rect 5328 0 5340 111
rect 5520 0 5532 111
rect 6264 0 6276 111
rect 6480 0 6492 111
rect 6672 0 6684 111
rect 7416 0 7428 111
rect 7632 0 7644 111
rect 7824 0 7836 111
rect 8568 0 8580 111
rect 8784 0 8796 111
rect 8976 0 8988 111
rect 9720 0 9732 111
rect 9936 0 9948 111
rect 10128 0 10140 111
rect 10872 0 10884 111
rect 11088 0 11100 111
rect 11280 0 11292 111
rect 12024 0 12036 111
rect 12096 41 12108 111
rect 12240 0 12252 111
rect 12312 19 12324 111
use Pc_slice  Pc_slice_0
timestamp 1394475379
transform 1 0 0 0 1 111
box 0 0 2952 1042
use mux2  mux2_0
timestamp 1386235218
transform 1 0 2952 0 1 177
box 0 0 192 799
use regBlock_slice  regBlock_slice_0
timestamp 1394475337
transform 1 0 3144 0 1 111
box 0 0 9216 1042
<< labels >>
rlabel metal1 3096 100 3096 100 1 SysBus
rlabel metal1 12353 34 12353 34 1 Rd1
rlabel metal1 12355 11 12355 11 1 Rd2
rlabel metal2 216 0 228 0 1 PcIncCin
rlabel metal2 360 0 372 0 1 LrSel
rlabel metal2 576 0 588 0 1 LrWe
rlabel metal2 1320 0 1332 0 1 LrEn
rlabel metal2 1488 0 1500 0 1 PcSel[0]
rlabel metal2 1872 0 1884 0 1 PcSel[1]
rlabel metal2 2088 0 2100 0 1 PcWe
rlabel metal2 2832 0 2844 0 1 PcEn
rlabel metal2 3000 0 3012 0 1 WdSel
rlabel metal2 3960 0 3972 0 1 Rs1[0]
rlabel metal2 4368 0 4380 0 1 Rw[1]
rlabel metal2 5112 0 5124 0 1 Rs1[1]
rlabel metal2 5328 0 5340 0 1 Rs2[1]
rlabel metal2 5520 0 5532 0 1 Rw[2]
rlabel metal2 6264 0 6276 0 1 Rs1[2]
rlabel metal2 6480 0 6492 0 1 Rs2[2]
rlabel metal2 6672 0 6684 0 1 Rw[3]
rlabel metal2 7416 0 7428 0 1 Rs1[3]
rlabel metal2 7632 0 7644 0 1 Rs2[3]
rlabel metal2 7824 0 7836 0 1 Rw[4]
rlabel metal2 8568 0 8580 0 1 Rs1[4]
rlabel metal2 8784 0 8796 0 1 Rs2[4]
rlabel metal2 8976 0 8988 0 1 Rw[5]
rlabel metal2 9720 0 9732 0 1 Rs1[5]
rlabel metal2 9936 0 9948 0 1 Rs2[5]
rlabel metal2 10128 0 10140 0 1 Rw[6]
rlabel metal2 10872 0 10884 0 1 Rs1[6]
rlabel metal2 11088 0 11100 0 1 Rs2[6]
rlabel metal2 11280 0 11292 0 1 Rw[7]
rlabel metal2 12024 0 12036 0 1 Rs1[7]
rlabel metal2 12240 0 12252 0 1 Rs2[7]
rlabel metal1 12352 100 12352 100 1 SysBus
rlabel metal1 12353 78 12353 78 1 Imm
rlabel metal1 12354 56 12354 56 1 Pc
rlabel metal2 3216 0 3228 0 1 Rw[0]
rlabel metal2 4176 0 4188 0 1 Rs2[0]
rlabel metal1 0 95 0 105 1 SysBus
rlabel metal1 0 73 0 83 1 Imm
rlabel metal1 12358 1164 12358 1164 6 AluOut
rlabel metal2 12240 1176 12252 1176 5 Rs2[7]
rlabel metal2 12024 1176 12036 1176 5 Rs1[7]
rlabel metal2 11280 1176 11292 1176 5 Rw[7]
rlabel metal2 11088 1176 11100 1176 5 Rs2[6]
rlabel metal2 10872 1176 10884 1176 5 Rs1[6]
rlabel metal2 10128 1176 10140 1176 5 Rw[6]
rlabel metal2 9720 1176 9732 1176 5 Rs1[5]
rlabel metal2 9936 1176 9948 1176 5 Rs2[5]
rlabel metal2 8976 1176 8988 1176 5 Rw[5]
rlabel metal2 8784 1176 8796 1176 5 Rs2[4]
rlabel metal2 8568 1176 8580 1176 5 Rs1[4]
rlabel metal2 7824 1176 7836 1176 5 Rw[4]
rlabel metal2 7632 1176 7644 1176 5 Rs2[3]
rlabel metal2 7416 1176 7428 1176 5 Rs1[3]
rlabel metal2 6672 1176 6684 1176 5 Rw[3]
rlabel metal2 6480 1176 6492 1176 5 Rs2[2]
rlabel metal2 6264 1176 6276 1176 5 Rs1[2]
rlabel metal2 5520 1176 5532 1176 5 Rw[2]
rlabel metal2 5328 1176 5340 1176 5 Rs2[1]
rlabel metal2 5112 1176 5124 1176 5 Rs1[1]
rlabel metal2 4368 1176 4380 1176 5 Rw[1]
rlabel metal2 4176 1176 4188 1176 5 Rs2[0]
rlabel metal2 3960 1176 3972 1176 5 Rs1[0]
rlabel metal2 3216 1176 3228 1176 5 Rw[0]
rlabel metal2 3000 1176 3012 1176 5 WdSel
rlabel metal2 2832 1176 2844 1176 5 PcEn
rlabel metal2 2088 1176 2100 1176 5 PcWe
rlabel metal2 1872 1176 1884 1176 5 PcSel[1]
rlabel metal2 1488 1176 1500 1176 5 PcSel[0]
rlabel metal2 1320 1176 1332 1176 5 LrEn
rlabel metal2 576 1176 588 1176 5 LrWe
rlabel metal2 360 1176 372 1176 5 LrSel
rlabel metal2 216 1176 228 1176 5 PcIncCout
<< end >>
