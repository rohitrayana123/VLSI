magic
tech c035u
timestamp 1395701949
<< metal1 >>
rect 9544 7964 9562 7978
rect 9496 7942 12206 7952
rect 9280 7918 21062 7928
rect 9160 7894 13826 7904
rect 17836 7894 17882 7904
rect 19444 7894 23354 7904
rect 5416 7868 5434 7882
rect 7288 7870 10058 7880
rect 10384 7868 10402 7882
rect 13816 7870 14330 7880
rect 17032 7870 21890 7880
rect 22660 7870 24482 7880
rect 4744 7846 14630 7856
rect 16228 7846 24410 7856
rect 3736 7822 19454 7832
rect 22168 7822 23474 7832
rect 24016 7822 25826 7832
rect 2584 7798 11390 7808
rect 12040 7798 12602 7808
rect 12616 7798 16850 7808
rect 16864 7798 25778 7808
rect 84 7774 1730 7784
rect 2392 7774 6098 7784
rect 6736 7774 25754 7784
rect 25792 7774 26451 7784
rect 84 7750 11162 7760
rect 12664 7750 22670 7760
rect 25696 7748 25714 7762
rect 25744 7750 25778 7760
rect 25816 7750 26451 7760
rect 3208 7726 6002 7736
rect 7720 7726 17846 7736
rect 19144 7726 25802 7736
rect 25840 7726 26451 7736
rect 4024 7702 5786 7712
rect 5920 7700 5938 7714
rect 8008 7702 10574 7712
rect 14152 7702 24278 7712
rect 25792 7702 26451 7712
rect 4840 7678 5762 7688
rect 8080 7676 8098 7690
rect 8920 7678 12986 7688
rect 17728 7678 20258 7688
rect 25768 7678 26451 7688
rect 25755 7649 26091 7659
rect 25755 7626 26091 7636
rect 25755 7588 26091 7613
rect 25755 6943 26091 6968
rect 13336 6845 23282 6855
rect 12520 6821 13322 6831
rect 13336 6821 20018 6831
rect 12328 6797 12578 6807
rect 13264 6797 13346 6807
rect 13408 6797 21554 6807
rect 12064 6773 24866 6783
rect 12040 6749 22322 6759
rect 11848 6725 19346 6735
rect 11392 6701 19874 6711
rect 11128 6677 16106 6687
rect 11104 6653 17258 6663
rect 17272 6653 20738 6663
rect 11080 6629 17858 6639
rect 17872 6629 25298 6639
rect 9640 6605 18458 6615
rect 9544 6581 20234 6591
rect 9400 6557 18818 6567
rect 23776 6557 24290 6567
rect 9208 6533 10346 6543
rect 10360 6533 17618 6543
rect 17632 6533 19442 6543
rect 19456 6533 23762 6543
rect 9112 6509 9434 6519
rect 9448 6509 15050 6519
rect 8944 6485 9266 6495
rect 9328 6485 11426 6495
rect 11440 6485 16178 6495
rect 16192 6485 22010 6495
rect 8920 6461 9650 6471
rect 9664 6461 15530 6471
rect 15544 6461 18842 6471
rect 18856 6461 22058 6471
rect 22072 6461 25442 6471
rect 25456 6461 25922 6471
rect 8680 6437 25418 6447
rect 8512 6413 11882 6423
rect 11896 6413 12146 6423
rect 12280 6413 14378 6423
rect 14392 6413 23522 6423
rect 8392 6389 9554 6399
rect 9568 6389 10586 6399
rect 10600 6389 11186 6399
rect 11200 6389 12290 6399
rect 12304 6389 19010 6399
rect 19024 6389 21410 6399
rect 21424 6389 23594 6399
rect 8248 6365 12530 6375
rect 13216 6365 23906 6375
rect 8224 6341 8234 6351
rect 8344 6341 10274 6351
rect 10288 6341 22682 6351
rect 8152 6317 13970 6327
rect 7984 6293 24890 6303
rect 7816 6269 10154 6279
rect 10168 6269 13538 6279
rect 7768 6245 10394 6255
rect 10408 6245 14546 6255
rect 14560 6245 15218 6255
rect 15232 6245 19754 6255
rect 7648 6221 9698 6231
rect 9712 6221 19250 6231
rect 7528 6197 9026 6207
rect 9088 6197 23378 6207
rect 7504 6173 19202 6183
rect 19216 6173 21722 6183
rect 7384 6149 12602 6159
rect 13096 6149 15074 6159
rect 15088 6149 23642 6159
rect 7192 6125 17186 6135
rect 17200 6125 19202 6135
rect 6880 6101 15794 6111
rect 17968 6101 19346 6111
rect 6712 6077 7922 6087
rect 7936 6077 13826 6087
rect 13840 6077 19106 6087
rect 19120 6077 23522 6087
rect 23536 6077 23978 6087
rect 6664 6053 19178 6063
rect 19312 6053 21914 6063
rect 6568 6029 21146 6039
rect 6472 6005 9818 6015
rect 9880 6005 21482 6015
rect 22984 6005 23258 6015
rect 24496 6005 24650 6015
rect 6448 5981 12482 5991
rect 12784 5981 21338 5991
rect 21352 5981 22034 5991
rect 22048 5981 24482 5991
rect 6400 5957 8210 5967
rect 8224 5957 13394 5967
rect 15520 5957 24530 5967
rect 6208 5933 8570 5943
rect 8584 5933 23042 5943
rect 6184 5909 6290 5919
rect 6304 5909 12362 5919
rect 12376 5909 19970 5919
rect 19984 5909 22970 5919
rect 6160 5885 8522 5895
rect 8632 5885 23210 5895
rect 6112 5861 6314 5871
rect 6328 5861 6914 5871
rect 6928 5861 14690 5871
rect 14704 5861 21554 5871
rect 21568 5861 22394 5871
rect 22408 5861 23546 5871
rect 23560 5861 24794 5871
rect 6040 5837 7490 5847
rect 7576 5837 14138 5847
rect 14152 5837 23018 5847
rect 6016 5813 6122 5823
rect 6136 5813 12338 5823
rect 12352 5813 14666 5823
rect 14680 5813 20114 5823
rect 20128 5813 21578 5823
rect 21592 5813 22802 5823
rect 22816 5813 24218 5823
rect 5944 5789 9842 5799
rect 9904 5789 20378 5799
rect 5824 5765 6410 5775
rect 6424 5765 19730 5775
rect 19744 5765 20354 5775
rect 20368 5765 21842 5775
rect 5800 5741 8018 5751
rect 8032 5741 8090 5751
rect 8104 5741 14474 5751
rect 14488 5741 19298 5751
rect 19312 5741 24098 5751
rect 5680 5717 12650 5727
rect 12664 5717 20162 5727
rect 5632 5693 23882 5703
rect 5536 5669 15842 5679
rect 17392 5669 24914 5679
rect 5368 5645 14186 5655
rect 14200 5645 21818 5655
rect 5296 5621 6650 5631
rect 6664 5621 24386 5631
rect 5296 5597 19370 5607
rect 5200 5573 7610 5583
rect 7624 5573 22490 5583
rect 5176 5549 6530 5559
rect 6544 5549 7658 5559
rect 7672 5549 10898 5559
rect 10912 5549 19010 5559
rect 5128 5525 6026 5535
rect 6040 5525 19538 5535
rect 5008 5501 10706 5511
rect 10792 5501 16610 5511
rect 17056 5501 23306 5511
rect 4936 5477 20114 5487
rect 4888 5453 9890 5463
rect 10024 5453 11546 5463
rect 11632 5453 25010 5463
rect 4888 5429 24362 5439
rect 4816 5405 8930 5415
rect 8944 5405 10730 5415
rect 10744 5405 16250 5415
rect 16264 5405 22538 5415
rect 22552 5405 24554 5415
rect 24568 5405 25874 5415
rect 4696 5381 9122 5391
rect 9136 5381 13514 5391
rect 13528 5381 14306 5391
rect 14320 5381 24314 5391
rect 4648 5357 17978 5367
rect 4648 5333 21074 5343
rect 4528 5309 15170 5319
rect 15184 5309 15314 5319
rect 15328 5309 20954 5319
rect 4432 5285 16826 5295
rect 16840 5285 21218 5295
rect 4384 5261 6890 5271
rect 6904 5261 16298 5271
rect 16312 5261 17498 5271
rect 17560 5261 18506 5271
rect 21760 5261 22730 5271
rect 4312 5237 6434 5247
rect 6448 5237 7778 5247
rect 7792 5237 9122 5247
rect 9184 5237 13610 5247
rect 15400 5237 15674 5247
rect 16456 5237 24938 5247
rect 4264 5213 21674 5223
rect 21688 5213 21746 5223
rect 4216 5189 12506 5199
rect 12736 5189 12842 5199
rect 12928 5189 13586 5199
rect 15376 5189 18026 5199
rect 18112 5189 19130 5199
rect 4168 5165 6410 5175
rect 6424 5165 7850 5175
rect 7864 5165 10898 5175
rect 10912 5165 14618 5175
rect 14632 5165 20546 5175
rect 4120 5141 6986 5151
rect 7000 5141 7850 5151
rect 7864 5141 8354 5151
rect 8368 5141 12194 5151
rect 12208 5141 15578 5151
rect 15592 5141 18722 5151
rect 21976 5141 22130 5151
rect 4096 5117 4106 5127
rect 4168 5117 9506 5127
rect 9520 5117 17570 5127
rect 17584 5117 17738 5127
rect 17752 5117 24602 5127
rect 4072 5093 5834 5103
rect 5848 5093 5930 5103
rect 5944 5093 10538 5103
rect 10552 5093 22850 5103
rect 22864 5093 25370 5103
rect 25384 5093 25610 5103
rect 4024 5069 9362 5079
rect 9472 5069 13442 5079
rect 15352 5069 23978 5079
rect 3976 5045 5978 5055
rect 5992 5045 7370 5055
rect 7384 5045 8474 5055
rect 8488 5045 14810 5055
rect 14824 5045 17210 5055
rect 17224 5045 19970 5055
rect 19984 5045 21962 5055
rect 21976 5045 23402 5055
rect 23416 5045 24674 5055
rect 3928 5021 15122 5031
rect 15136 5021 15650 5031
rect 16216 5021 22082 5031
rect 25240 5021 25250 5031
rect 3904 4997 11258 5007
rect 11320 4997 23642 5007
rect 23656 4997 25226 5007
rect 3880 4973 8450 4983
rect 8464 4973 10226 4983
rect 10336 4973 21098 4983
rect 3808 4949 4754 4959
rect 4768 4949 7346 4959
rect 7360 4949 13034 4959
rect 13048 4949 25490 4959
rect 3688 4925 25274 4935
rect 3664 4901 18434 4911
rect 3640 4877 9770 4887
rect 9784 4877 12386 4887
rect 12400 4877 14354 4887
rect 14368 4877 18338 4887
rect 18352 4877 21098 4887
rect 21112 4877 23714 4887
rect 3568 4853 11210 4863
rect 11224 4853 13178 4863
rect 13192 4853 19226 4863
rect 19696 4853 20762 4863
rect 3520 4829 12458 4839
rect 12472 4829 15554 4839
rect 15880 4829 18146 4839
rect 19672 4829 20882 4839
rect 3472 4805 12890 4815
rect 12904 4805 24074 4815
rect 3424 4781 11978 4791
rect 11992 4781 21194 4791
rect 21208 4781 23474 4791
rect 3400 4757 6290 4767
rect 6304 4757 18674 4767
rect 19504 4757 26090 4767
rect 3328 4733 3602 4743
rect 3616 4733 5906 4743
rect 5920 4733 7634 4743
rect 7648 4733 8810 4743
rect 8824 4733 10082 4743
rect 10096 4733 14882 4743
rect 14896 4733 19034 4743
rect 19048 4733 22874 4743
rect 3304 4709 16994 4719
rect 17008 4709 23570 4719
rect 3232 4685 9386 4695
rect 9400 4685 10514 4695
rect 10528 4685 10922 4695
rect 10936 4685 15194 4695
rect 15208 4685 18410 4695
rect 18424 4685 24410 4695
rect 3184 4661 4274 4671
rect 4288 4661 6218 4671
rect 6232 4661 8426 4671
rect 8440 4661 8498 4671
rect 8512 4661 13562 4671
rect 14104 4661 14150 4671
rect 15256 4661 15626 4671
rect 15832 4661 17714 4671
rect 17896 4661 22922 4671
rect 3112 4637 19562 4647
rect 19576 4637 21794 4647
rect 3064 4613 5066 4623
rect 5080 4613 7250 4623
rect 7264 4613 15386 4623
rect 15400 4613 16946 4623
rect 16960 4613 20042 4623
rect 3064 4589 21122 4599
rect 21448 4589 21530 4599
rect 3016 4565 3770 4575
rect 3784 4565 5042 4575
rect 5056 4565 5474 4575
rect 5488 4565 6674 4575
rect 6688 4565 8138 4575
rect 8200 4565 11018 4575
rect 11032 4565 19946 4575
rect 21256 4565 24122 4575
rect 24136 4565 25130 4575
rect 2968 4541 10946 4551
rect 10960 4541 13610 4551
rect 13624 4541 16322 4551
rect 16336 4541 18602 4551
rect 18616 4541 20978 4551
rect 20992 4541 23066 4551
rect 23944 4541 24434 4551
rect 2944 4517 4058 4527
rect 4072 4517 6626 4527
rect 6640 4517 8906 4527
rect 8920 4517 14090 4527
rect 14104 4517 17114 4527
rect 17128 4517 17282 4527
rect 17296 4517 20330 4527
rect 20344 4517 22610 4527
rect 22624 4517 23930 4527
rect 2896 4493 14282 4503
rect 15208 4493 15530 4503
rect 15712 4493 22130 4503
rect 2872 4469 7226 4479
rect 7240 4469 9746 4479
rect 9760 4469 15002 4479
rect 15160 4469 18554 4479
rect 18880 4469 23858 4479
rect 2800 4445 13730 4455
rect 15040 4445 17882 4455
rect 17896 4445 23042 4455
rect 2752 4421 19154 4431
rect 19432 4421 22274 4431
rect 2728 4397 7586 4407
rect 7720 4397 21434 4407
rect 2704 4373 10610 4383
rect 10672 4373 17666 4383
rect 17776 4373 18350 4383
rect 18784 4373 18938 4383
rect 19336 4373 24026 4383
rect 2680 4349 10418 4359
rect 10480 4349 13730 4359
rect 14464 4349 21386 4359
rect 23128 4349 23486 4359
rect 23848 4349 24626 4359
rect 2656 4325 22898 4335
rect 23104 4325 23126 4335
rect 23176 4325 24002 4335
rect 2608 4301 20282 4311
rect 20704 4301 22778 4311
rect 22792 4301 24650 4311
rect 25096 4301 26451 4311
rect 2560 4277 14234 4287
rect 14320 4277 14378 4287
rect 14440 4277 19274 4287
rect 19288 4277 24266 4287
rect 25072 4277 25094 4287
rect 25384 4277 25442 4287
rect 2560 4253 6746 4263
rect 6808 4253 6866 4263
rect 6976 4253 9002 4263
rect 9016 4253 19994 4263
rect 20008 4253 20090 4263
rect 20104 4253 24194 4263
rect 25408 4253 26114 4263
rect 2536 4229 7274 4239
rect 7288 4229 7946 4239
rect 8176 4229 10634 4239
rect 10648 4229 10670 4239
rect 10684 4229 20282 4239
rect 20296 4229 22202 4239
rect 22216 4229 23954 4239
rect 24088 4229 24530 4239
rect 2464 4205 3698 4215
rect 3760 4205 15602 4215
rect 16792 4205 17930 4215
rect 18136 4205 23786 4215
rect 24112 4205 24722 4215
rect 2416 4181 5114 4191
rect 5128 4181 9026 4191
rect 9040 4181 15242 4191
rect 15304 4181 21986 4191
rect 2344 4157 12866 4167
rect 12880 4157 14738 4167
rect 14752 4157 16730 4167
rect 16744 4157 17450 4167
rect 17464 4157 23426 4167
rect 2320 4133 4514 4143
rect 4528 4133 6170 4143
rect 6184 4133 6362 4143
rect 6376 4133 19610 4143
rect 19624 4133 21170 4143
rect 21184 4133 25466 4143
rect 2248 4109 13250 4119
rect 13432 4109 24530 4119
rect 2200 4085 4466 4095
rect 4480 4085 8282 4095
rect 8296 4085 11474 4095
rect 11488 4085 22514 4095
rect 2128 4061 3818 4071
rect 3832 4061 12866 4071
rect 12880 4061 15506 4071
rect 17680 4061 19922 4071
rect 20008 4061 20018 4071
rect 20176 4061 22106 4071
rect 22120 4061 22946 4071
rect 2104 4037 22994 4047
rect 2056 4013 18578 4023
rect 18592 4013 21938 4023
rect 23008 4013 23546 4023
rect 1984 3989 3458 3999
rect 3472 3989 4490 3999
rect 4504 3989 7130 3999
rect 7144 3989 10298 3999
rect 10312 3989 18314 3999
rect 20584 3989 23690 3999
rect 1936 3965 4562 3975
rect 4624 3965 15266 3975
rect 18256 3965 23330 3975
rect 1912 3941 2234 3951
rect 2248 3941 4610 3951
rect 4624 3941 4826 3951
rect 4840 3941 5138 3951
rect 5152 3941 6314 3951
rect 6328 3941 9626 3951
rect 9640 3941 10874 3951
rect 10888 3941 13946 3951
rect 14344 3941 18218 3951
rect 18328 3941 18578 3951
rect 21088 3941 21146 3951
rect 21208 3941 24146 3951
rect 1888 3917 10202 3927
rect 10288 3917 10346 3927
rect 10528 3917 10586 3927
rect 10840 3917 21674 3927
rect 23344 3917 24122 3927
rect 1864 3893 17834 3903
rect 21184 3893 21218 3903
rect 21352 3893 22466 3903
rect 1840 3869 17786 3879
rect 21256 3869 24338 3879
rect 1816 3845 2210 3855
rect 2224 3845 2258 3855
rect 2272 3845 4082 3855
rect 4096 3845 4946 3855
rect 4960 3845 5450 3855
rect 5464 3845 6626 3855
rect 6640 3845 7874 3855
rect 7888 3845 10730 3855
rect 10744 3845 11138 3855
rect 11152 3845 13082 3855
rect 13096 3845 13154 3855
rect 13168 3845 22538 3855
rect 84 3821 6842 3831
rect 6856 3821 20834 3831
rect 21376 3821 23858 3831
rect 23872 3821 24986 3831
rect 84 3797 15410 3807
rect 17800 3797 21458 3807
rect 1624 3773 6794 3783
rect 6856 3773 6890 3783
rect 7072 3773 17930 3783
rect 1624 3749 3074 3759
rect 3088 3749 6506 3759
rect 6520 3749 7322 3759
rect 7336 3749 9146 3759
rect 9160 3749 9530 3759
rect 9544 3749 10610 3759
rect 10624 3749 11690 3759
rect 11704 3749 13274 3759
rect 13288 3749 15410 3759
rect 15424 3749 15962 3759
rect 15976 3749 18914 3759
rect 18928 3749 22178 3759
rect 22192 3749 22226 3759
rect 22240 3749 24386 3759
rect 1648 3725 5402 3735
rect 5416 3725 8570 3735
rect 8584 3725 10178 3735
rect 10192 3725 12722 3735
rect 12736 3725 17114 3735
rect 17128 3725 17546 3735
rect 17560 3725 24170 3735
rect 1672 3701 2426 3711
rect 2488 3701 10370 3711
rect 10840 3701 17354 3711
rect 1696 3677 4346 3687
rect 4360 3677 7418 3687
rect 7432 3677 12218 3687
rect 12232 3677 18098 3687
rect 18112 3677 18194 3687
rect 1744 3653 22586 3663
rect 1744 3629 9578 3639
rect 9688 3629 18050 3639
rect 18064 3629 22706 3639
rect 22720 3629 23810 3639
rect 1792 3605 20786 3615
rect 22720 3605 22922 3615
rect 2008 3581 20906 3591
rect 2152 3557 26066 3567
rect 2224 3533 2234 3543
rect 2296 3533 3434 3543
rect 3448 3533 4178 3543
rect 4192 3533 6050 3543
rect 6064 3533 6482 3543
rect 6496 3533 15434 3543
rect 15448 3533 17426 3543
rect 17440 3533 17906 3543
rect 17920 3533 18530 3543
rect 18544 3533 23306 3543
rect 23320 3533 25154 3543
rect 2368 3509 12530 3519
rect 12928 3509 12986 3519
rect 13192 3509 14150 3519
rect 14464 3509 20642 3519
rect 2464 3485 9194 3495
rect 9208 3485 9242 3495
rect 9256 3485 17690 3495
rect 2536 3461 24506 3471
rect 2632 3437 24242 3447
rect 24520 3437 24530 3447
rect 2656 3413 12818 3423
rect 13000 3413 22658 3423
rect 2680 3389 7898 3399
rect 7912 3389 12074 3399
rect 12136 3389 12158 3399
rect 12208 3389 12290 3399
rect 12472 3389 12602 3399
rect 13528 3389 15674 3399
rect 15688 3389 17810 3399
rect 17824 3389 22562 3399
rect 2776 3365 20690 3375
rect 2824 3341 10970 3351
rect 10984 3341 14114 3351
rect 14128 3341 20834 3351
rect 2848 3317 11090 3327
rect 11344 3317 16994 3327
rect 17368 3317 17858 3327
rect 2872 3293 8306 3303
rect 8320 3293 13490 3303
rect 13504 3293 14066 3303
rect 14080 3293 16490 3303
rect 16504 3293 17090 3303
rect 17104 3293 22754 3303
rect 2896 3269 4946 3279
rect 4960 3269 7394 3279
rect 7408 3269 10418 3279
rect 10432 3269 16274 3279
rect 16288 3269 20066 3279
rect 20080 3269 20186 3279
rect 20200 3269 21986 3279
rect 22000 3269 23090 3279
rect 23104 3269 25010 3279
rect 2944 3245 6602 3255
rect 6616 3245 18290 3255
rect 18304 3245 22418 3255
rect 22768 3245 23018 3255
rect 3136 3221 23690 3231
rect 3352 3197 6746 3207
rect 6832 3197 15554 3207
rect 17104 3197 17498 3207
rect 18304 3197 18554 3207
rect 22432 3197 22778 3207
rect 3424 3173 4922 3183
rect 4936 3173 17234 3183
rect 17248 3173 18626 3183
rect 18640 3173 19634 3183
rect 19648 3173 20042 3183
rect 20056 3173 22442 3183
rect 3664 3149 4298 3159
rect 4312 3149 7010 3159
rect 7024 3149 9986 3159
rect 10000 3149 10154 3159
rect 10168 3149 11354 3159
rect 11368 3149 11714 3159
rect 11728 3149 16850 3159
rect 16864 3149 17018 3159
rect 17032 3149 17522 3159
rect 17536 3149 18746 3159
rect 22456 3149 22802 3159
rect 3736 3125 5594 3135
rect 5608 3125 6266 3135
rect 6280 3125 7034 3135
rect 7048 3125 7154 3135
rect 7168 3125 12746 3135
rect 12760 3125 13370 3135
rect 13384 3125 14570 3135
rect 14584 3125 17306 3135
rect 17320 3125 17426 3135
rect 17440 3125 18074 3135
rect 18088 3125 20306 3135
rect 20320 3125 23906 3135
rect 23920 3125 24578 3135
rect 24592 3125 25058 3135
rect 25072 3125 25202 3135
rect 3784 3101 16058 3111
rect 3832 3077 7442 3087
rect 7456 3077 14810 3087
rect 14824 3077 20474 3087
rect 3856 3053 5882 3063
rect 5896 3053 14786 3063
rect 14800 3053 17594 3063
rect 17608 3053 19034 3063
rect 19048 3053 19850 3063
rect 3880 3029 4106 3039
rect 4120 3029 8066 3039
rect 8080 3029 10442 3039
rect 10456 3029 11138 3039
rect 11152 3029 12434 3039
rect 12448 3029 12770 3039
rect 12784 3029 15482 3039
rect 15496 3029 16250 3039
rect 16264 3029 23126 3039
rect 23140 3029 24770 3039
rect 3952 3005 12314 3015
rect 12328 3005 25178 3015
rect 3976 2981 5690 2991
rect 5704 2981 6866 2991
rect 6880 2981 8066 2991
rect 8080 2981 10850 2991
rect 10864 2981 12578 2991
rect 12592 2981 12842 2991
rect 12856 2981 23354 2991
rect 4000 2957 6554 2967
rect 6616 2957 6674 2967
rect 6784 2957 25514 2967
rect 4024 2933 8258 2943
rect 8272 2933 11786 2943
rect 11800 2933 17330 2943
rect 17344 2933 20642 2943
rect 4120 2909 13274 2919
rect 13288 2909 21290 2919
rect 4216 2885 5210 2895
rect 5224 2885 6506 2895
rect 6520 2885 8378 2895
rect 8392 2885 8402 2895
rect 8416 2885 12098 2895
rect 12112 2885 13298 2895
rect 13504 2885 13538 2895
rect 13720 2885 22370 2895
rect 4288 2861 5858 2871
rect 5872 2861 10634 2871
rect 10648 2861 11666 2871
rect 11680 2861 12242 2871
rect 12256 2861 13346 2871
rect 13360 2861 24698 2871
rect 4384 2837 4682 2847
rect 4696 2837 5306 2847
rect 5320 2837 10562 2847
rect 10576 2837 17450 2847
rect 4408 2813 5762 2823
rect 5776 2813 5954 2823
rect 5968 2813 8594 2823
rect 8608 2813 12794 2823
rect 12808 2813 14906 2823
rect 14920 2813 16274 2823
rect 16288 2813 16370 2823
rect 16384 2813 19826 2823
rect 19840 2813 21650 2823
rect 21664 2813 22250 2823
rect 22264 2813 23114 2823
rect 23128 2813 23570 2823
rect 4456 2789 5498 2799
rect 5512 2789 17138 2799
rect 17152 2789 21506 2799
rect 22264 2789 22490 2799
rect 4504 2765 4514 2775
rect 4600 2765 19586 2775
rect 4528 2741 13058 2751
rect 13072 2741 14858 2751
rect 14872 2741 15098 2751
rect 15112 2741 16442 2751
rect 16456 2741 17762 2751
rect 17776 2741 18266 2751
rect 18280 2741 23186 2751
rect 23200 2741 23834 2751
rect 4552 2717 15914 2727
rect 15928 2717 17522 2727
rect 4600 2693 12554 2703
rect 15016 2693 23738 2703
rect 23752 2693 24194 2703
rect 4720 2669 4850 2679
rect 4864 2669 9434 2679
rect 9448 2669 12242 2679
rect 12256 2669 12410 2679
rect 12424 2669 13634 2679
rect 13648 2669 15626 2679
rect 15640 2669 19874 2679
rect 19888 2669 22322 2679
rect 4840 2645 18962 2655
rect 5056 2621 16466 2631
rect 16480 2621 25094 2631
rect 25108 2621 25322 2631
rect 5248 2597 9290 2607
rect 9424 2597 12122 2607
rect 12136 2597 18386 2607
rect 5584 2573 9938 2583
rect 10000 2573 18170 2583
rect 18184 2573 23234 2583
rect 5704 2549 13154 2559
rect 13168 2549 21890 2559
rect 21904 2549 22154 2559
rect 5728 2525 22298 2535
rect 6112 2501 25682 2511
rect 6256 2477 7538 2487
rect 7552 2477 12002 2487
rect 12016 2477 21866 2487
rect 21880 2477 24458 2487
rect 6352 2453 7538 2463
rect 7672 2453 15770 2463
rect 17344 2453 17738 2463
rect 6544 2429 24818 2439
rect 6712 2405 21770 2415
rect 7048 2381 8234 2391
rect 8632 2381 18506 2391
rect 18520 2381 22826 2391
rect 7096 2357 16514 2367
rect 7096 2333 8834 2343
rect 8896 2333 13466 2343
rect 13480 2333 21002 2343
rect 7192 2309 7442 2319
rect 7456 2309 8978 2319
rect 8992 2309 15314 2319
rect 15328 2309 25346 2319
rect 7288 2285 16034 2295
rect 16048 2285 23486 2295
rect 7336 2261 9962 2271
rect 10048 2261 19466 2271
rect 7576 2237 15458 2247
rect 7720 2213 24434 2223
rect 7792 2189 25034 2199
rect 7888 2165 8786 2175
rect 8872 2165 18482 2175
rect 18496 2165 23666 2175
rect 7960 2141 25730 2151
rect 8704 2117 23162 2127
rect 8752 2093 24050 2103
rect 8776 2069 9338 2079
rect 9352 2069 16154 2079
rect 8824 2045 10490 2055
rect 10504 2045 11234 2055
rect 11248 2045 11930 2055
rect 11944 2045 21626 2055
rect 21640 2045 22346 2055
rect 22360 2045 23234 2055
rect 8968 2021 18350 2031
rect 18364 2021 19706 2031
rect 22360 2021 22730 2031
rect 9016 1997 9914 2007
rect 10072 1997 10130 2007
rect 10144 1997 12158 2007
rect 12172 1997 21530 2007
rect 21544 1997 23618 2007
rect 23632 1997 24218 2007
rect 24232 1997 24290 2007
rect 24304 1997 25562 2007
rect 9088 1973 9218 1983
rect 9328 1973 17162 1983
rect 9472 1949 17642 1959
rect 9856 1925 19058 1935
rect 9928 1901 10106 1911
rect 10120 1901 20426 1911
rect 10120 1877 10130 1887
rect 10216 1877 10226 1887
rect 10336 1877 19658 1887
rect 19672 1877 24002 1887
rect 10360 1853 26451 1863
rect 10576 1829 10670 1839
rect 11056 1829 18002 1839
rect 11584 1805 12794 1815
rect 15112 1805 17402 1815
rect 17416 1805 17474 1815
rect 11752 1781 23450 1791
rect 11824 1757 17042 1767
rect 17488 1757 22634 1767
rect 22648 1757 23258 1767
rect 12016 1733 13418 1743
rect 13432 1733 14210 1743
rect 14224 1733 19778 1743
rect 26128 1733 26451 1743
rect 12568 1709 25250 1719
rect 26104 1709 26451 1719
rect 16912 876 17642 886
rect 18160 876 23498 886
rect 16408 852 19394 862
rect 19552 852 24434 862
rect 15352 828 21290 838
rect 13360 804 25514 814
rect 13312 780 16658 790
rect 16720 780 24338 790
rect 12976 756 13562 766
rect 13576 756 22514 766
rect 12640 732 13202 742
rect 13216 732 24290 742
rect 11320 708 21122 718
rect 22144 708 25346 718
rect 11272 684 16538 694
rect 16600 684 21026 694
rect 22072 684 24122 694
rect 11080 660 12674 670
rect 12856 660 24530 670
rect 11032 636 22466 646
rect 22648 636 22898 646
rect 10720 612 25250 622
rect 9736 588 12338 598
rect 12352 588 15458 598
rect 15712 588 18866 598
rect 19240 588 24650 598
rect 9592 564 23474 574
rect 9352 540 22850 550
rect 9256 516 10442 526
rect 10672 516 14282 526
rect 14392 516 26090 526
rect 7744 492 10778 502
rect 10840 490 10858 504
rect 11008 492 14498 502
rect 14848 492 23426 502
rect 7708 468 8282 478
rect 8488 468 23258 478
rect 7312 444 13658 454
rect 13888 444 22658 454
rect 7240 420 19154 430
rect 19432 420 20594 430
rect 20680 418 20698 432
rect 7144 396 18218 406
rect 18352 396 20954 406
rect 6208 372 13778 382
rect 14152 372 21314 382
rect 5992 348 7826 358
rect 8416 348 20858 358
rect 5896 324 7106 334
rect 7216 324 8522 334
rect 8704 324 17834 334
rect 5872 300 6890 310
rect 6904 300 8834 310
rect 8848 300 10130 310
rect 10144 300 16970 310
rect 16984 300 19058 310
rect 19072 300 22202 310
rect 5656 276 22778 286
rect 5176 252 9746 262
rect 9760 252 10250 262
rect 10264 252 12362 262
rect 12424 252 26114 262
rect 4816 228 19082 238
rect 4336 204 9866 214
rect 10312 204 19466 214
rect 3904 180 6722 190
rect 6976 180 17138 190
rect 2776 156 16106 166
rect 16360 156 19562 166
rect 2752 132 11834 142
rect 12616 132 22802 142
rect 22816 132 24314 142
rect 2584 108 8306 118
rect 8728 108 14018 118
rect 15136 108 19634 118
rect 84 84 13010 94
rect 13120 84 24026 94
rect 26104 84 26451 94
rect 84 60 1730 70
rect 2416 60 10946 70
rect 10960 60 19514 70
rect 26104 60 26451 70
rect 9808 36 26090 46
rect 26128 36 26451 46
rect 17056 10 17074 24
rect 26080 12 26451 22
<< m2contact >>
rect 9530 7964 9544 7978
rect 9482 7940 9496 7954
rect 12206 7940 12220 7954
rect 9266 7916 9280 7930
rect 21062 7916 21076 7930
rect 9146 7892 9160 7906
rect 13826 7892 13840 7906
rect 17822 7892 17836 7906
rect 17882 7892 17896 7906
rect 19430 7892 19444 7906
rect 23354 7892 23368 7906
rect 5402 7868 5416 7882
rect 7274 7868 7288 7882
rect 10058 7868 10072 7882
rect 10370 7868 10384 7882
rect 13802 7868 13816 7882
rect 14330 7868 14344 7882
rect 17018 7868 17032 7882
rect 21890 7868 21904 7882
rect 22646 7868 22660 7882
rect 24482 7868 24496 7882
rect 4730 7844 4744 7858
rect 14630 7844 14644 7858
rect 16214 7844 16228 7858
rect 24410 7844 24424 7858
rect 3722 7820 3736 7834
rect 19454 7820 19468 7834
rect 22154 7820 22168 7834
rect 23474 7820 23488 7834
rect 24002 7820 24016 7834
rect 25826 7820 25840 7834
rect 2570 7796 2584 7810
rect 11390 7796 11404 7810
rect 12026 7796 12040 7810
rect 12602 7796 12616 7810
rect 16850 7796 16864 7810
rect 25778 7796 25792 7810
rect 70 7772 84 7786
rect 1730 7772 1744 7786
rect 2378 7772 2392 7786
rect 6098 7772 6112 7786
rect 6722 7772 6736 7786
rect 25754 7772 25768 7786
rect 25778 7772 25792 7786
rect 26451 7772 26465 7786
rect 70 7748 84 7762
rect 11162 7748 11176 7762
rect 12650 7748 12664 7762
rect 22670 7748 22684 7762
rect 25682 7748 25696 7762
rect 25730 7748 25744 7762
rect 25778 7748 25792 7762
rect 25802 7748 25816 7762
rect 26451 7748 26465 7762
rect 3194 7724 3208 7738
rect 6002 7724 6016 7738
rect 7706 7724 7720 7738
rect 17846 7724 17860 7738
rect 19130 7724 19144 7738
rect 25802 7724 25816 7738
rect 25826 7724 25840 7738
rect 26451 7724 26465 7738
rect 4010 7700 4024 7714
rect 5786 7700 5800 7714
rect 5906 7700 5920 7714
rect 7994 7700 8008 7714
rect 10574 7700 10588 7714
rect 14138 7700 14152 7714
rect 24278 7700 24292 7714
rect 25778 7700 25792 7714
rect 26451 7700 26465 7714
rect 4826 7676 4840 7690
rect 5762 7676 5776 7690
rect 8066 7676 8080 7690
rect 8906 7676 8920 7690
rect 12986 7676 13000 7690
rect 17714 7676 17728 7690
rect 20258 7676 20272 7690
rect 25754 7676 25768 7690
rect 26451 7676 26465 7690
rect 13322 6843 13336 6857
rect 23282 6843 23296 6857
rect 12506 6819 12520 6833
rect 13322 6819 13336 6833
rect 20018 6819 20032 6833
rect 12314 6795 12328 6809
rect 12578 6795 12592 6809
rect 13250 6795 13264 6809
rect 13346 6795 13360 6809
rect 13394 6795 13408 6809
rect 21554 6795 21568 6809
rect 12050 6771 12064 6785
rect 24866 6771 24880 6785
rect 12026 6747 12040 6761
rect 22322 6747 22336 6761
rect 11834 6723 11848 6737
rect 19346 6723 19360 6737
rect 11378 6699 11392 6713
rect 19874 6699 19888 6713
rect 11114 6675 11128 6689
rect 16106 6675 16120 6689
rect 11090 6651 11104 6665
rect 17258 6651 17272 6665
rect 20738 6651 20752 6665
rect 11066 6627 11080 6641
rect 17858 6627 17872 6641
rect 25298 6627 25312 6641
rect 9626 6603 9640 6617
rect 18458 6603 18472 6617
rect 9530 6579 9544 6593
rect 20234 6579 20248 6593
rect 9386 6555 9400 6569
rect 18818 6555 18832 6569
rect 23762 6555 23776 6569
rect 24290 6555 24304 6569
rect 9194 6531 9208 6545
rect 10346 6531 10360 6545
rect 17618 6531 17632 6545
rect 19442 6531 19456 6545
rect 23762 6531 23776 6545
rect 9098 6507 9112 6521
rect 9434 6507 9448 6521
rect 15050 6507 15064 6521
rect 8930 6483 8944 6497
rect 9266 6483 9280 6497
rect 9314 6483 9328 6497
rect 11426 6483 11440 6497
rect 16178 6483 16192 6497
rect 22010 6483 22024 6497
rect 8906 6459 8920 6473
rect 9650 6459 9664 6473
rect 15530 6459 15544 6473
rect 18842 6459 18856 6473
rect 22058 6459 22072 6473
rect 25442 6459 25456 6473
rect 25922 6459 25936 6473
rect 8666 6435 8680 6449
rect 25418 6435 25432 6449
rect 8498 6411 8512 6425
rect 11882 6411 11896 6425
rect 12146 6411 12160 6425
rect 12266 6411 12280 6425
rect 14378 6411 14392 6425
rect 23522 6411 23536 6425
rect 8378 6387 8392 6401
rect 9554 6387 9568 6401
rect 10586 6387 10600 6401
rect 11186 6387 11200 6401
rect 12290 6387 12304 6401
rect 19010 6387 19024 6401
rect 21410 6387 21424 6401
rect 23594 6387 23608 6401
rect 8234 6363 8248 6377
rect 12530 6363 12544 6377
rect 13202 6363 13216 6377
rect 23906 6363 23920 6377
rect 8210 6339 8224 6353
rect 8234 6339 8248 6353
rect 8330 6339 8344 6353
rect 10274 6339 10288 6353
rect 22682 6339 22696 6353
rect 8138 6315 8152 6329
rect 13970 6315 13984 6329
rect 7970 6291 7984 6305
rect 24890 6291 24904 6305
rect 7802 6267 7816 6281
rect 10154 6267 10168 6281
rect 13538 6267 13552 6281
rect 7754 6243 7768 6257
rect 10394 6243 10408 6257
rect 14546 6243 14560 6257
rect 15218 6243 15232 6257
rect 19754 6243 19768 6257
rect 7634 6219 7648 6233
rect 9698 6219 9712 6233
rect 19250 6219 19264 6233
rect 7514 6195 7528 6209
rect 9026 6195 9040 6209
rect 9074 6195 9088 6209
rect 23378 6195 23392 6209
rect 7490 6171 7504 6185
rect 19202 6171 19216 6185
rect 21722 6171 21736 6185
rect 7370 6147 7384 6161
rect 12602 6147 12616 6161
rect 13082 6147 13096 6161
rect 15074 6147 15088 6161
rect 23642 6147 23656 6161
rect 7178 6123 7192 6137
rect 17186 6123 17200 6137
rect 19202 6123 19216 6137
rect 6866 6099 6880 6113
rect 15794 6099 15808 6113
rect 17954 6099 17968 6113
rect 19346 6099 19360 6113
rect 6698 6075 6712 6089
rect 7922 6075 7936 6089
rect 13826 6075 13840 6089
rect 19106 6075 19120 6089
rect 23522 6075 23536 6089
rect 23978 6075 23992 6089
rect 6650 6051 6664 6065
rect 19178 6051 19192 6065
rect 19298 6051 19312 6065
rect 21914 6051 21928 6065
rect 6554 6027 6568 6041
rect 21146 6027 21160 6041
rect 6458 6003 6472 6017
rect 9818 6003 9832 6017
rect 9866 6003 9880 6017
rect 21482 6003 21496 6017
rect 22970 6003 22984 6017
rect 23258 6003 23272 6017
rect 24482 6003 24496 6017
rect 24650 6003 24664 6017
rect 6434 5979 6448 5993
rect 12482 5979 12496 5993
rect 12770 5979 12784 5993
rect 21338 5979 21352 5993
rect 22034 5979 22048 5993
rect 24482 5979 24496 5993
rect 6386 5955 6400 5969
rect 8210 5955 8224 5969
rect 13394 5955 13408 5969
rect 15506 5955 15520 5969
rect 24530 5955 24544 5969
rect 6194 5931 6208 5945
rect 8570 5931 8584 5945
rect 23042 5931 23056 5945
rect 6170 5907 6184 5921
rect 6290 5907 6304 5921
rect 12362 5907 12376 5921
rect 19970 5907 19984 5921
rect 22970 5907 22984 5921
rect 6146 5883 6160 5897
rect 8522 5883 8536 5897
rect 8618 5883 8632 5897
rect 23210 5883 23224 5897
rect 6098 5859 6112 5873
rect 6314 5859 6328 5873
rect 6914 5859 6928 5873
rect 14690 5859 14704 5873
rect 21554 5859 21568 5873
rect 22394 5859 22408 5873
rect 23546 5859 23560 5873
rect 24794 5859 24808 5873
rect 6026 5835 6040 5849
rect 7490 5835 7504 5849
rect 7562 5835 7576 5849
rect 14138 5835 14152 5849
rect 23018 5835 23032 5849
rect 6002 5811 6016 5825
rect 6122 5811 6136 5825
rect 12338 5811 12352 5825
rect 14666 5811 14680 5825
rect 20114 5811 20128 5825
rect 21578 5811 21592 5825
rect 22802 5811 22816 5825
rect 24218 5811 24232 5825
rect 5930 5787 5944 5801
rect 9842 5787 9856 5801
rect 9890 5787 9904 5801
rect 20378 5787 20392 5801
rect 5810 5763 5824 5777
rect 6410 5763 6424 5777
rect 19730 5763 19744 5777
rect 20354 5763 20368 5777
rect 21842 5763 21856 5777
rect 5786 5739 5800 5753
rect 8018 5739 8032 5753
rect 8090 5739 8104 5753
rect 14474 5739 14488 5753
rect 19298 5739 19312 5753
rect 24098 5739 24112 5753
rect 5666 5715 5680 5729
rect 12650 5715 12664 5729
rect 20162 5715 20176 5729
rect 5618 5691 5632 5705
rect 23882 5691 23896 5705
rect 5522 5667 5536 5681
rect 15842 5667 15856 5681
rect 17378 5667 17392 5681
rect 24914 5667 24928 5681
rect 5354 5643 5368 5657
rect 14186 5643 14200 5657
rect 21818 5643 21832 5657
rect 5282 5619 5296 5633
rect 6650 5619 6664 5633
rect 24386 5619 24400 5633
rect 5282 5595 5296 5609
rect 19370 5595 19384 5609
rect 5186 5571 5200 5585
rect 7610 5571 7624 5585
rect 22490 5571 22504 5585
rect 5162 5547 5176 5561
rect 6530 5547 6544 5561
rect 7658 5547 7672 5561
rect 10898 5547 10912 5561
rect 19010 5547 19024 5561
rect 5114 5523 5128 5537
rect 6026 5523 6040 5537
rect 19538 5523 19552 5537
rect 4994 5499 5008 5513
rect 10706 5499 10720 5513
rect 10778 5499 10792 5513
rect 16610 5499 16624 5513
rect 17042 5499 17056 5513
rect 23306 5499 23320 5513
rect 4922 5475 4936 5489
rect 20114 5475 20128 5489
rect 4874 5451 4888 5465
rect 9890 5451 9904 5465
rect 10010 5451 10024 5465
rect 11546 5451 11560 5465
rect 11618 5451 11632 5465
rect 25010 5451 25024 5465
rect 4874 5427 4888 5441
rect 24362 5427 24376 5441
rect 4802 5403 4816 5417
rect 8930 5403 8944 5417
rect 10730 5403 10744 5417
rect 16250 5403 16264 5417
rect 22538 5403 22552 5417
rect 24554 5403 24568 5417
rect 25874 5403 25888 5417
rect 4682 5379 4696 5393
rect 9122 5379 9136 5393
rect 13514 5379 13528 5393
rect 14306 5379 14320 5393
rect 24314 5379 24328 5393
rect 4634 5355 4648 5369
rect 17978 5355 17992 5369
rect 4634 5331 4648 5345
rect 21074 5331 21088 5345
rect 4514 5307 4528 5321
rect 15170 5307 15184 5321
rect 15314 5307 15328 5321
rect 20954 5307 20968 5321
rect 4418 5283 4432 5297
rect 16826 5283 16840 5297
rect 21218 5283 21232 5297
rect 4370 5259 4384 5273
rect 6890 5259 6904 5273
rect 16298 5259 16312 5273
rect 17498 5259 17512 5273
rect 17546 5259 17560 5273
rect 18506 5259 18520 5273
rect 21746 5259 21760 5273
rect 22730 5259 22744 5273
rect 4298 5235 4312 5249
rect 6434 5235 6448 5249
rect 7778 5235 7792 5249
rect 9122 5235 9136 5249
rect 9170 5235 9184 5249
rect 13610 5235 13624 5249
rect 15386 5235 15400 5249
rect 15674 5235 15688 5249
rect 16442 5235 16456 5249
rect 24938 5235 24952 5249
rect 4250 5211 4264 5225
rect 21674 5211 21688 5225
rect 21746 5211 21760 5225
rect 4202 5187 4216 5201
rect 12506 5187 12520 5201
rect 12722 5187 12736 5201
rect 12842 5187 12856 5201
rect 12914 5187 12928 5201
rect 13586 5187 13600 5201
rect 15362 5187 15376 5201
rect 18026 5187 18040 5201
rect 18098 5187 18112 5201
rect 19130 5187 19144 5201
rect 4154 5163 4168 5177
rect 6410 5163 6424 5177
rect 7850 5163 7864 5177
rect 10898 5163 10912 5177
rect 14618 5163 14632 5177
rect 20546 5163 20560 5177
rect 4106 5139 4120 5153
rect 6986 5139 7000 5153
rect 7850 5139 7864 5153
rect 8354 5139 8368 5153
rect 12194 5139 12208 5153
rect 15578 5139 15592 5153
rect 18722 5139 18736 5153
rect 21962 5139 21976 5153
rect 22130 5139 22144 5153
rect 4082 5115 4096 5129
rect 4106 5115 4120 5129
rect 4154 5115 4168 5129
rect 9506 5115 9520 5129
rect 17570 5115 17584 5129
rect 17738 5115 17752 5129
rect 24602 5115 24616 5129
rect 4058 5091 4072 5105
rect 5834 5091 5848 5105
rect 5930 5091 5944 5105
rect 10538 5091 10552 5105
rect 22850 5091 22864 5105
rect 25370 5091 25384 5105
rect 25610 5091 25624 5105
rect 4010 5067 4024 5081
rect 9362 5067 9376 5081
rect 9458 5067 9472 5081
rect 13442 5067 13456 5081
rect 15338 5067 15352 5081
rect 23978 5067 23992 5081
rect 3962 5043 3976 5057
rect 5978 5043 5992 5057
rect 7370 5043 7384 5057
rect 8474 5043 8488 5057
rect 14810 5043 14824 5057
rect 17210 5043 17224 5057
rect 19970 5043 19984 5057
rect 21962 5043 21976 5057
rect 23402 5043 23416 5057
rect 24674 5043 24688 5057
rect 3914 5019 3928 5033
rect 15122 5019 15136 5033
rect 15650 5019 15664 5033
rect 16202 5019 16216 5033
rect 22082 5019 22096 5033
rect 25226 5019 25240 5033
rect 25250 5019 25264 5033
rect 3890 4995 3904 5009
rect 11258 4995 11272 5009
rect 11306 4995 11320 5009
rect 23642 4995 23656 5009
rect 25226 4995 25240 5009
rect 3866 4971 3880 4985
rect 8450 4971 8464 4985
rect 10226 4971 10240 4985
rect 10322 4971 10336 4985
rect 21098 4971 21112 4985
rect 3794 4947 3808 4961
rect 4754 4947 4768 4961
rect 7346 4947 7360 4961
rect 13034 4947 13048 4961
rect 25490 4947 25504 4961
rect 3674 4923 3688 4937
rect 25274 4923 25288 4937
rect 3650 4899 3664 4913
rect 18434 4899 18448 4913
rect 3626 4875 3640 4889
rect 9770 4875 9784 4889
rect 12386 4875 12400 4889
rect 14354 4875 14368 4889
rect 18338 4875 18352 4889
rect 21098 4875 21112 4889
rect 23714 4875 23728 4889
rect 3554 4851 3568 4865
rect 11210 4851 11224 4865
rect 13178 4851 13192 4865
rect 19226 4851 19240 4865
rect 19682 4851 19696 4865
rect 20762 4851 20776 4865
rect 3506 4827 3520 4841
rect 12458 4827 12472 4841
rect 15554 4827 15568 4841
rect 15866 4827 15880 4841
rect 18146 4827 18160 4841
rect 19658 4827 19672 4841
rect 20882 4827 20896 4841
rect 3458 4803 3472 4817
rect 12890 4803 12904 4817
rect 24074 4803 24088 4817
rect 3410 4779 3424 4793
rect 11978 4779 11992 4793
rect 21194 4779 21208 4793
rect 23474 4779 23488 4793
rect 3386 4755 3400 4769
rect 6290 4755 6304 4769
rect 18674 4755 18688 4769
rect 19490 4755 19504 4769
rect 26090 4755 26104 4769
rect 3314 4731 3328 4745
rect 3602 4731 3616 4745
rect 5906 4731 5920 4745
rect 7634 4731 7648 4745
rect 8810 4731 8824 4745
rect 10082 4731 10096 4745
rect 14882 4731 14896 4745
rect 19034 4731 19048 4745
rect 22874 4731 22888 4745
rect 3290 4707 3304 4721
rect 16994 4707 17008 4721
rect 23570 4707 23584 4721
rect 3218 4683 3232 4697
rect 9386 4683 9400 4697
rect 10514 4683 10528 4697
rect 10922 4683 10936 4697
rect 15194 4683 15208 4697
rect 18410 4683 18424 4697
rect 24410 4683 24424 4697
rect 3170 4659 3184 4673
rect 4274 4659 4288 4673
rect 6218 4659 6232 4673
rect 8426 4659 8440 4673
rect 8498 4659 8512 4673
rect 13562 4659 13576 4673
rect 14090 4659 14104 4673
rect 14150 4659 14164 4673
rect 15242 4659 15256 4673
rect 15626 4659 15640 4673
rect 15818 4659 15832 4673
rect 17714 4659 17728 4673
rect 17882 4659 17896 4673
rect 22922 4659 22936 4673
rect 3098 4635 3112 4649
rect 19562 4635 19576 4649
rect 21794 4635 21808 4649
rect 3050 4611 3064 4625
rect 5066 4611 5080 4625
rect 7250 4611 7264 4625
rect 15386 4611 15400 4625
rect 16946 4611 16960 4625
rect 20042 4611 20056 4625
rect 3050 4587 3064 4601
rect 21122 4587 21136 4601
rect 21434 4587 21448 4601
rect 21530 4587 21544 4601
rect 3002 4563 3016 4577
rect 3770 4563 3784 4577
rect 5042 4563 5056 4577
rect 5474 4563 5488 4577
rect 6674 4563 6688 4577
rect 8138 4563 8152 4577
rect 8186 4563 8200 4577
rect 11018 4563 11032 4577
rect 19946 4563 19960 4577
rect 21242 4563 21256 4577
rect 24122 4563 24136 4577
rect 25130 4563 25144 4577
rect 2954 4539 2968 4553
rect 10946 4539 10960 4553
rect 13610 4539 13624 4553
rect 16322 4539 16336 4553
rect 18602 4539 18616 4553
rect 20978 4539 20992 4553
rect 23066 4539 23080 4553
rect 23930 4539 23944 4553
rect 24434 4539 24448 4553
rect 2930 4515 2944 4529
rect 4058 4515 4072 4529
rect 6626 4515 6640 4529
rect 8906 4515 8920 4529
rect 14090 4515 14104 4529
rect 17114 4515 17128 4529
rect 17282 4515 17296 4529
rect 20330 4515 20344 4529
rect 22610 4515 22624 4529
rect 23930 4515 23944 4529
rect 2882 4491 2896 4505
rect 14282 4491 14296 4505
rect 15194 4491 15208 4505
rect 15530 4491 15544 4505
rect 15698 4491 15712 4505
rect 22130 4491 22144 4505
rect 2858 4467 2872 4481
rect 7226 4467 7240 4481
rect 9746 4467 9760 4481
rect 15002 4467 15016 4481
rect 15146 4467 15160 4481
rect 18554 4467 18568 4481
rect 18866 4467 18880 4481
rect 23858 4467 23872 4481
rect 2786 4443 2800 4457
rect 13730 4443 13744 4457
rect 15026 4443 15040 4457
rect 17882 4443 17896 4457
rect 23042 4443 23056 4457
rect 2738 4419 2752 4433
rect 19154 4419 19168 4433
rect 19418 4419 19432 4433
rect 22274 4419 22288 4433
rect 2714 4395 2728 4409
rect 7586 4395 7600 4409
rect 7706 4395 7720 4409
rect 21434 4395 21448 4409
rect 2690 4371 2704 4385
rect 10610 4371 10624 4385
rect 10658 4371 10672 4385
rect 17666 4371 17680 4385
rect 17762 4371 17776 4385
rect 18350 4371 18364 4385
rect 18770 4371 18784 4385
rect 18938 4371 18952 4385
rect 19322 4371 19336 4385
rect 24026 4371 24040 4385
rect 2666 4347 2680 4361
rect 10418 4347 10432 4361
rect 10466 4347 10480 4361
rect 13730 4347 13744 4361
rect 14450 4347 14464 4361
rect 21386 4347 21400 4361
rect 23114 4347 23128 4361
rect 23486 4347 23500 4361
rect 23834 4347 23848 4361
rect 24626 4347 24640 4361
rect 2642 4323 2656 4337
rect 22898 4323 22912 4337
rect 23090 4323 23104 4337
rect 23126 4323 23140 4337
rect 23162 4323 23176 4337
rect 24002 4323 24016 4337
rect 2594 4299 2608 4313
rect 20282 4299 20296 4313
rect 20690 4299 20704 4313
rect 22778 4299 22792 4313
rect 24650 4299 24664 4313
rect 25082 4299 25096 4313
rect 26451 4299 26465 4313
rect 2546 4275 2560 4289
rect 14234 4275 14248 4289
rect 14306 4275 14320 4289
rect 14378 4275 14392 4289
rect 14426 4275 14440 4289
rect 19274 4275 19288 4289
rect 24266 4275 24280 4289
rect 25058 4275 25072 4289
rect 25094 4275 25108 4289
rect 25370 4275 25384 4289
rect 25442 4275 25456 4289
rect 2546 4251 2560 4265
rect 6746 4251 6760 4265
rect 6794 4251 6808 4265
rect 6866 4251 6880 4265
rect 6962 4251 6976 4265
rect 9002 4251 9016 4265
rect 19994 4251 20008 4265
rect 20090 4251 20104 4265
rect 24194 4251 24208 4265
rect 25394 4251 25408 4265
rect 26114 4251 26128 4265
rect 2522 4227 2536 4241
rect 7274 4227 7288 4241
rect 7946 4227 7960 4241
rect 8162 4227 8176 4241
rect 10634 4227 10648 4241
rect 10670 4227 10684 4241
rect 20282 4227 20296 4241
rect 22202 4227 22216 4241
rect 23954 4227 23968 4241
rect 24074 4227 24088 4241
rect 24530 4227 24544 4241
rect 2450 4203 2464 4217
rect 3698 4203 3712 4217
rect 3746 4203 3760 4217
rect 15602 4203 15616 4217
rect 16778 4203 16792 4217
rect 17930 4203 17944 4217
rect 18122 4203 18136 4217
rect 23786 4203 23800 4217
rect 24098 4203 24112 4217
rect 24722 4203 24736 4217
rect 2402 4179 2416 4193
rect 5114 4179 5128 4193
rect 9026 4179 9040 4193
rect 15242 4179 15256 4193
rect 15290 4179 15304 4193
rect 21986 4179 22000 4193
rect 2330 4155 2344 4169
rect 12866 4155 12880 4169
rect 14738 4155 14752 4169
rect 16730 4155 16744 4169
rect 17450 4155 17464 4169
rect 23426 4155 23440 4169
rect 2306 4131 2320 4145
rect 4514 4131 4528 4145
rect 6170 4131 6184 4145
rect 6362 4131 6376 4145
rect 19610 4131 19624 4145
rect 21170 4131 21184 4145
rect 25466 4131 25480 4145
rect 2234 4107 2248 4121
rect 13250 4107 13264 4121
rect 13418 4107 13432 4121
rect 24530 4107 24544 4121
rect 2186 4083 2200 4097
rect 4466 4083 4480 4097
rect 8282 4083 8296 4097
rect 11474 4083 11488 4097
rect 22514 4083 22528 4097
rect 2114 4059 2128 4073
rect 3818 4059 3832 4073
rect 12866 4059 12880 4073
rect 15506 4059 15520 4073
rect 17666 4059 17680 4073
rect 19922 4059 19936 4073
rect 19994 4059 20008 4073
rect 20018 4059 20032 4073
rect 20162 4059 20176 4073
rect 22106 4059 22120 4073
rect 22946 4059 22960 4073
rect 2090 4035 2104 4049
rect 22994 4035 23008 4049
rect 2042 4011 2056 4025
rect 18578 4011 18592 4025
rect 21938 4011 21952 4025
rect 22994 4011 23008 4025
rect 23546 4011 23560 4025
rect 1970 3987 1984 4001
rect 3458 3987 3472 4001
rect 4490 3987 4504 4001
rect 7130 3987 7144 4001
rect 10298 3987 10312 4001
rect 18314 3987 18328 4001
rect 20570 3987 20584 4001
rect 23690 3987 23704 4001
rect 1922 3963 1936 3977
rect 4562 3963 4576 3977
rect 4610 3963 4624 3977
rect 15266 3963 15280 3977
rect 18242 3963 18256 3977
rect 23330 3963 23344 3977
rect 1898 3939 1912 3953
rect 2234 3939 2248 3953
rect 4610 3939 4624 3953
rect 4826 3939 4840 3953
rect 5138 3939 5152 3953
rect 6314 3939 6328 3953
rect 9626 3939 9640 3953
rect 10874 3939 10888 3953
rect 13946 3939 13960 3953
rect 14330 3939 14344 3953
rect 18218 3939 18232 3953
rect 18314 3939 18328 3953
rect 18578 3939 18592 3953
rect 21074 3939 21088 3953
rect 21146 3939 21160 3953
rect 21194 3939 21208 3953
rect 24146 3939 24160 3953
rect 1874 3915 1888 3929
rect 10202 3915 10216 3929
rect 10274 3915 10288 3929
rect 10346 3915 10360 3929
rect 10514 3915 10528 3929
rect 10586 3915 10600 3929
rect 10826 3915 10840 3929
rect 21674 3915 21688 3929
rect 23330 3915 23344 3929
rect 24122 3915 24136 3929
rect 1850 3891 1864 3905
rect 17834 3891 17848 3905
rect 21170 3891 21184 3905
rect 21218 3891 21232 3905
rect 21338 3891 21352 3905
rect 22466 3891 22480 3905
rect 1826 3867 1840 3881
rect 17786 3867 17800 3881
rect 21242 3867 21256 3881
rect 24338 3867 24352 3881
rect 1802 3843 1816 3857
rect 2210 3843 2224 3857
rect 2258 3843 2272 3857
rect 4082 3843 4096 3857
rect 4946 3843 4960 3857
rect 5450 3843 5464 3857
rect 6626 3843 6640 3857
rect 7874 3843 7888 3857
rect 10730 3843 10744 3857
rect 11138 3843 11152 3857
rect 13082 3843 13096 3857
rect 13154 3843 13168 3857
rect 22538 3843 22552 3857
rect 70 3819 84 3833
rect 6842 3819 6856 3833
rect 20834 3819 20848 3833
rect 21362 3819 21376 3833
rect 23858 3819 23872 3833
rect 24986 3819 25000 3833
rect 70 3795 84 3809
rect 15410 3795 15424 3809
rect 17786 3795 17800 3809
rect 21458 3795 21472 3809
rect 1610 3771 1624 3785
rect 6794 3771 6808 3785
rect 6842 3771 6856 3785
rect 6890 3771 6904 3785
rect 7058 3771 7072 3785
rect 17930 3771 17944 3785
rect 1610 3747 1624 3761
rect 3074 3747 3088 3761
rect 6506 3747 6520 3761
rect 7322 3747 7336 3761
rect 9146 3747 9160 3761
rect 9530 3747 9544 3761
rect 10610 3747 10624 3761
rect 11690 3747 11704 3761
rect 13274 3747 13288 3761
rect 15410 3747 15424 3761
rect 15962 3747 15976 3761
rect 18914 3747 18928 3761
rect 22178 3747 22192 3761
rect 22226 3747 22240 3761
rect 24386 3747 24400 3761
rect 1634 3723 1648 3737
rect 5402 3723 5416 3737
rect 8570 3723 8584 3737
rect 10178 3723 10192 3737
rect 12722 3723 12736 3737
rect 17114 3723 17128 3737
rect 17546 3723 17560 3737
rect 24170 3723 24184 3737
rect 1658 3699 1672 3713
rect 2426 3699 2440 3713
rect 2474 3699 2488 3713
rect 10370 3699 10384 3713
rect 10826 3699 10840 3713
rect 17354 3699 17368 3713
rect 1682 3675 1696 3689
rect 4346 3675 4360 3689
rect 7418 3675 7432 3689
rect 12218 3675 12232 3689
rect 18098 3675 18112 3689
rect 18194 3675 18208 3689
rect 1730 3651 1744 3665
rect 22586 3651 22600 3665
rect 1730 3627 1744 3641
rect 9578 3627 9592 3641
rect 9674 3627 9688 3641
rect 18050 3627 18064 3641
rect 22706 3627 22720 3641
rect 23810 3627 23824 3641
rect 1778 3603 1792 3617
rect 20786 3603 20800 3617
rect 22706 3603 22720 3617
rect 22922 3603 22936 3617
rect 1994 3579 2008 3593
rect 20906 3579 20920 3593
rect 2138 3555 2152 3569
rect 26066 3555 26080 3569
rect 2210 3531 2224 3545
rect 2234 3531 2248 3545
rect 2282 3531 2296 3545
rect 3434 3531 3448 3545
rect 4178 3531 4192 3545
rect 6050 3531 6064 3545
rect 6482 3531 6496 3545
rect 15434 3531 15448 3545
rect 17426 3531 17440 3545
rect 17906 3531 17920 3545
rect 18530 3531 18544 3545
rect 23306 3531 23320 3545
rect 25154 3531 25168 3545
rect 2354 3507 2368 3521
rect 12530 3507 12544 3521
rect 12914 3507 12928 3521
rect 12986 3507 13000 3521
rect 13178 3507 13192 3521
rect 14150 3507 14164 3521
rect 14450 3507 14464 3521
rect 20642 3507 20656 3521
rect 2450 3483 2464 3497
rect 9194 3483 9208 3497
rect 9242 3483 9256 3497
rect 17690 3483 17704 3497
rect 2522 3459 2536 3473
rect 24506 3459 24520 3473
rect 2618 3435 2632 3449
rect 24242 3435 24256 3449
rect 24506 3435 24520 3449
rect 24530 3435 24544 3449
rect 2642 3411 2656 3425
rect 12818 3411 12832 3425
rect 12986 3411 13000 3425
rect 22658 3411 22672 3425
rect 2666 3387 2680 3401
rect 7898 3387 7912 3401
rect 12074 3387 12088 3401
rect 12122 3387 12136 3401
rect 12158 3387 12172 3401
rect 12194 3387 12208 3401
rect 12290 3387 12304 3401
rect 12458 3387 12472 3401
rect 12602 3387 12616 3401
rect 13514 3387 13528 3401
rect 15674 3387 15688 3401
rect 17810 3387 17824 3401
rect 22562 3387 22576 3401
rect 2762 3363 2776 3377
rect 20690 3363 20704 3377
rect 2810 3339 2824 3353
rect 10970 3339 10984 3353
rect 14114 3339 14128 3353
rect 20834 3339 20848 3353
rect 2834 3315 2848 3329
rect 11090 3315 11104 3329
rect 11330 3315 11344 3329
rect 16994 3315 17008 3329
rect 17354 3315 17368 3329
rect 17858 3315 17872 3329
rect 2858 3291 2872 3305
rect 8306 3291 8320 3305
rect 13490 3291 13504 3305
rect 14066 3291 14080 3305
rect 16490 3291 16504 3305
rect 17090 3291 17104 3305
rect 22754 3291 22768 3305
rect 2882 3267 2896 3281
rect 4946 3267 4960 3281
rect 7394 3267 7408 3281
rect 10418 3267 10432 3281
rect 16274 3267 16288 3281
rect 20066 3267 20080 3281
rect 20186 3267 20200 3281
rect 21986 3267 22000 3281
rect 23090 3267 23104 3281
rect 25010 3267 25024 3281
rect 2930 3243 2944 3257
rect 6602 3243 6616 3257
rect 18290 3243 18304 3257
rect 22418 3243 22432 3257
rect 22754 3243 22768 3257
rect 23018 3243 23032 3257
rect 3122 3219 3136 3233
rect 23690 3219 23704 3233
rect 3338 3195 3352 3209
rect 6746 3195 6760 3209
rect 6818 3195 6832 3209
rect 15554 3195 15568 3209
rect 17090 3195 17104 3209
rect 17498 3195 17512 3209
rect 18290 3195 18304 3209
rect 18554 3195 18568 3209
rect 22418 3195 22432 3209
rect 22778 3195 22792 3209
rect 3410 3171 3424 3185
rect 4922 3171 4936 3185
rect 17234 3171 17248 3185
rect 18626 3171 18640 3185
rect 19634 3171 19648 3185
rect 20042 3171 20056 3185
rect 22442 3171 22456 3185
rect 3650 3147 3664 3161
rect 4298 3147 4312 3161
rect 7010 3147 7024 3161
rect 9986 3147 10000 3161
rect 10154 3147 10168 3161
rect 11354 3147 11368 3161
rect 11714 3147 11728 3161
rect 16850 3147 16864 3161
rect 17018 3147 17032 3161
rect 17522 3147 17536 3161
rect 18746 3147 18760 3161
rect 22442 3147 22456 3161
rect 22802 3147 22816 3161
rect 3722 3123 3736 3137
rect 5594 3123 5608 3137
rect 6266 3123 6280 3137
rect 7034 3123 7048 3137
rect 7154 3123 7168 3137
rect 12746 3123 12760 3137
rect 13370 3123 13384 3137
rect 14570 3123 14584 3137
rect 17306 3123 17320 3137
rect 17426 3123 17440 3137
rect 18074 3123 18088 3137
rect 20306 3123 20320 3137
rect 23906 3123 23920 3137
rect 24578 3123 24592 3137
rect 25058 3123 25072 3137
rect 25202 3123 25216 3137
rect 3770 3099 3784 3113
rect 16058 3099 16072 3113
rect 3818 3075 3832 3089
rect 7442 3075 7456 3089
rect 14810 3075 14824 3089
rect 20474 3075 20488 3089
rect 3842 3051 3856 3065
rect 5882 3051 5896 3065
rect 14786 3051 14800 3065
rect 17594 3051 17608 3065
rect 19034 3051 19048 3065
rect 19850 3051 19864 3065
rect 3866 3027 3880 3041
rect 4106 3027 4120 3041
rect 8066 3027 8080 3041
rect 10442 3027 10456 3041
rect 11138 3027 11152 3041
rect 12434 3027 12448 3041
rect 12770 3027 12784 3041
rect 15482 3027 15496 3041
rect 16250 3027 16264 3041
rect 23126 3027 23140 3041
rect 24770 3027 24784 3041
rect 3938 3003 3952 3017
rect 12314 3003 12328 3017
rect 25178 3003 25192 3017
rect 3962 2979 3976 2993
rect 5690 2979 5704 2993
rect 6866 2979 6880 2993
rect 8066 2979 8080 2993
rect 10850 2979 10864 2993
rect 12578 2979 12592 2993
rect 12842 2979 12856 2993
rect 23354 2979 23368 2993
rect 3986 2955 4000 2969
rect 6554 2955 6568 2969
rect 6602 2955 6616 2969
rect 6674 2955 6688 2969
rect 6770 2955 6784 2969
rect 25514 2955 25528 2969
rect 4010 2931 4024 2945
rect 8258 2931 8272 2945
rect 11786 2931 11800 2945
rect 17330 2931 17344 2945
rect 20642 2931 20656 2945
rect 4106 2907 4120 2921
rect 13274 2907 13288 2921
rect 21290 2907 21304 2921
rect 4202 2883 4216 2897
rect 5210 2883 5224 2897
rect 6506 2883 6520 2897
rect 8378 2883 8392 2897
rect 8402 2883 8416 2897
rect 12098 2883 12112 2897
rect 13298 2883 13312 2897
rect 13490 2883 13504 2897
rect 13538 2883 13552 2897
rect 13706 2883 13720 2897
rect 22370 2883 22384 2897
rect 4274 2859 4288 2873
rect 5858 2859 5872 2873
rect 10634 2859 10648 2873
rect 11666 2859 11680 2873
rect 12242 2859 12256 2873
rect 13346 2859 13360 2873
rect 24698 2859 24712 2873
rect 4370 2835 4384 2849
rect 4682 2835 4696 2849
rect 5306 2835 5320 2849
rect 10562 2835 10576 2849
rect 17450 2835 17464 2849
rect 4394 2811 4408 2825
rect 5762 2811 5776 2825
rect 5954 2811 5968 2825
rect 8594 2811 8608 2825
rect 12794 2811 12808 2825
rect 14906 2811 14920 2825
rect 16274 2811 16288 2825
rect 16370 2811 16384 2825
rect 19826 2811 19840 2825
rect 21650 2811 21664 2825
rect 22250 2811 22264 2825
rect 23114 2811 23128 2825
rect 23570 2811 23584 2825
rect 4442 2787 4456 2801
rect 5498 2787 5512 2801
rect 17138 2787 17152 2801
rect 21506 2787 21520 2801
rect 22250 2787 22264 2801
rect 22490 2787 22504 2801
rect 4490 2763 4504 2777
rect 4514 2763 4528 2777
rect 4586 2763 4600 2777
rect 19586 2763 19600 2777
rect 4514 2739 4528 2753
rect 13058 2739 13072 2753
rect 14858 2739 14872 2753
rect 15098 2739 15112 2753
rect 16442 2739 16456 2753
rect 17762 2739 17776 2753
rect 18266 2739 18280 2753
rect 23186 2739 23200 2753
rect 23834 2739 23848 2753
rect 4538 2715 4552 2729
rect 15914 2715 15928 2729
rect 17522 2715 17536 2729
rect 4586 2691 4600 2705
rect 12554 2691 12568 2705
rect 15002 2691 15016 2705
rect 23738 2691 23752 2705
rect 24194 2691 24208 2705
rect 4706 2667 4720 2681
rect 4850 2667 4864 2681
rect 9434 2667 9448 2681
rect 12242 2667 12256 2681
rect 12410 2667 12424 2681
rect 13634 2667 13648 2681
rect 15626 2667 15640 2681
rect 19874 2667 19888 2681
rect 22322 2667 22336 2681
rect 4826 2643 4840 2657
rect 18962 2643 18976 2657
rect 5042 2619 5056 2633
rect 16466 2619 16480 2633
rect 25094 2619 25108 2633
rect 25322 2619 25336 2633
rect 5234 2595 5248 2609
rect 9290 2595 9304 2609
rect 9410 2595 9424 2609
rect 12122 2595 12136 2609
rect 18386 2595 18400 2609
rect 5570 2571 5584 2585
rect 9938 2571 9952 2585
rect 9986 2571 10000 2585
rect 18170 2571 18184 2585
rect 23234 2571 23248 2585
rect 5690 2547 5704 2561
rect 13154 2547 13168 2561
rect 21890 2547 21904 2561
rect 22154 2547 22168 2561
rect 5714 2523 5728 2537
rect 22298 2523 22312 2537
rect 6098 2499 6112 2513
rect 25682 2499 25696 2513
rect 6242 2475 6256 2489
rect 7538 2475 7552 2489
rect 12002 2475 12016 2489
rect 21866 2475 21880 2489
rect 24458 2475 24472 2489
rect 6338 2451 6352 2465
rect 7538 2451 7552 2465
rect 7658 2451 7672 2465
rect 15770 2451 15784 2465
rect 17330 2451 17344 2465
rect 17738 2451 17752 2465
rect 6530 2427 6544 2441
rect 24818 2427 24832 2441
rect 6698 2403 6712 2417
rect 21770 2403 21784 2417
rect 7034 2379 7048 2393
rect 8234 2379 8248 2393
rect 8618 2379 8632 2393
rect 18506 2379 18520 2393
rect 22826 2379 22840 2393
rect 7082 2355 7096 2369
rect 16514 2355 16528 2369
rect 7082 2331 7096 2345
rect 8834 2331 8848 2345
rect 8882 2331 8896 2345
rect 13466 2331 13480 2345
rect 21002 2331 21016 2345
rect 7178 2307 7192 2321
rect 7442 2307 7456 2321
rect 8978 2307 8992 2321
rect 15314 2307 15328 2321
rect 25346 2307 25360 2321
rect 7274 2283 7288 2297
rect 16034 2283 16048 2297
rect 23486 2283 23500 2297
rect 7322 2259 7336 2273
rect 9962 2259 9976 2273
rect 10034 2259 10048 2273
rect 19466 2259 19480 2273
rect 7562 2235 7576 2249
rect 15458 2235 15472 2249
rect 7706 2211 7720 2225
rect 24434 2211 24448 2225
rect 7778 2187 7792 2201
rect 25034 2187 25048 2201
rect 7874 2163 7888 2177
rect 8786 2163 8800 2177
rect 8858 2163 8872 2177
rect 18482 2163 18496 2177
rect 23666 2163 23680 2177
rect 7946 2139 7960 2153
rect 25730 2139 25744 2153
rect 8690 2115 8704 2129
rect 23162 2115 23176 2129
rect 8738 2091 8752 2105
rect 24050 2091 24064 2105
rect 8762 2067 8776 2081
rect 9338 2067 9352 2081
rect 16154 2067 16168 2081
rect 8810 2043 8824 2057
rect 10490 2043 10504 2057
rect 11234 2043 11248 2057
rect 11930 2043 11944 2057
rect 21626 2043 21640 2057
rect 22346 2043 22360 2057
rect 23234 2043 23248 2057
rect 8954 2019 8968 2033
rect 18350 2019 18364 2033
rect 19706 2019 19720 2033
rect 22346 2019 22360 2033
rect 22730 2019 22744 2033
rect 9002 1995 9016 2009
rect 9914 1995 9928 2009
rect 10058 1995 10072 2009
rect 10130 1995 10144 2009
rect 12158 1995 12172 2009
rect 21530 1995 21544 2009
rect 23618 1995 23632 2009
rect 24218 1995 24232 2009
rect 24290 1995 24304 2009
rect 25562 1995 25576 2009
rect 9074 1971 9088 1985
rect 9218 1971 9232 1985
rect 9314 1971 9328 1985
rect 17162 1971 17176 1985
rect 9458 1947 9472 1961
rect 17642 1947 17656 1961
rect 9842 1923 9856 1937
rect 19058 1923 19072 1937
rect 9914 1899 9928 1913
rect 10106 1899 10120 1913
rect 20426 1899 20440 1913
rect 10106 1875 10120 1889
rect 10130 1875 10144 1889
rect 10202 1875 10216 1889
rect 10226 1875 10240 1889
rect 10322 1875 10336 1889
rect 19658 1875 19672 1889
rect 24002 1875 24016 1889
rect 10346 1851 10360 1865
rect 26451 1851 26465 1865
rect 10562 1827 10576 1841
rect 10670 1827 10684 1841
rect 11042 1827 11056 1841
rect 18002 1827 18016 1841
rect 11570 1803 11584 1817
rect 12794 1803 12808 1817
rect 15098 1803 15112 1817
rect 17402 1803 17416 1817
rect 17474 1803 17488 1817
rect 11738 1779 11752 1793
rect 23450 1779 23464 1793
rect 11810 1755 11824 1769
rect 17042 1755 17056 1769
rect 17474 1755 17488 1769
rect 22634 1755 22648 1769
rect 23258 1755 23272 1769
rect 12002 1731 12016 1745
rect 13418 1731 13432 1745
rect 14210 1731 14224 1745
rect 19778 1731 19792 1745
rect 26114 1731 26128 1745
rect 26451 1731 26465 1745
rect 12554 1707 12568 1721
rect 25250 1707 25264 1721
rect 26090 1707 26104 1721
rect 26451 1707 26465 1721
rect 16898 874 16912 888
rect 17642 874 17656 888
rect 18146 874 18160 888
rect 23498 874 23512 888
rect 16394 850 16408 864
rect 19394 850 19408 864
rect 19538 850 19552 864
rect 24434 850 24448 864
rect 15338 826 15352 840
rect 21290 826 21304 840
rect 13346 802 13360 816
rect 25514 802 25528 816
rect 13298 778 13312 792
rect 16658 778 16672 792
rect 16706 778 16720 792
rect 24338 778 24352 792
rect 12962 754 12976 768
rect 13562 754 13576 768
rect 22514 754 22528 768
rect 12626 730 12640 744
rect 13202 730 13216 744
rect 24290 730 24304 744
rect 11306 706 11320 720
rect 21122 706 21136 720
rect 22130 706 22144 720
rect 25346 706 25360 720
rect 11258 682 11272 696
rect 16538 682 16552 696
rect 16586 682 16600 696
rect 21026 682 21040 696
rect 22058 682 22072 696
rect 24122 682 24136 696
rect 11066 658 11080 672
rect 12674 658 12688 672
rect 12842 658 12856 672
rect 24530 658 24544 672
rect 11018 634 11032 648
rect 22466 634 22480 648
rect 22634 634 22648 648
rect 22898 634 22912 648
rect 10706 610 10720 624
rect 25250 610 25264 624
rect 9722 586 9736 600
rect 12338 586 12352 600
rect 15458 586 15472 600
rect 15698 586 15712 600
rect 18866 586 18880 600
rect 19226 586 19240 600
rect 24650 586 24664 600
rect 9578 562 9592 576
rect 23474 562 23488 576
rect 9338 538 9352 552
rect 22850 538 22864 552
rect 9242 514 9256 528
rect 10442 514 10456 528
rect 10658 514 10672 528
rect 14282 514 14296 528
rect 14378 514 14392 528
rect 26090 514 26104 528
rect 7730 490 7744 504
rect 10778 490 10792 504
rect 10826 490 10840 504
rect 10994 490 11008 504
rect 14498 490 14512 504
rect 14834 490 14848 504
rect 23426 490 23440 504
rect 7694 466 7708 480
rect 8282 466 8296 480
rect 8474 466 8488 480
rect 23258 466 23272 480
rect 7298 442 7312 456
rect 13658 442 13672 456
rect 13874 442 13888 456
rect 22658 442 22672 456
rect 7226 418 7240 432
rect 19154 418 19168 432
rect 19418 418 19432 432
rect 20594 418 20608 432
rect 20666 418 20680 432
rect 7130 394 7144 408
rect 18218 394 18232 408
rect 18338 394 18352 408
rect 20954 394 20968 408
rect 6194 370 6208 384
rect 13778 370 13792 384
rect 14138 370 14152 384
rect 21314 370 21328 384
rect 5978 346 5992 360
rect 7826 346 7840 360
rect 8402 346 8416 360
rect 20858 346 20872 360
rect 5882 322 5896 336
rect 7106 322 7120 336
rect 7202 322 7216 336
rect 8522 322 8536 336
rect 8690 322 8704 336
rect 17834 322 17848 336
rect 5858 298 5872 312
rect 6890 298 6904 312
rect 8834 298 8848 312
rect 10130 298 10144 312
rect 16970 298 16984 312
rect 19058 298 19072 312
rect 22202 298 22216 312
rect 5642 274 5656 288
rect 22778 274 22792 288
rect 5162 250 5176 264
rect 9746 250 9760 264
rect 10250 250 10264 264
rect 12362 250 12376 264
rect 12410 250 12424 264
rect 26114 250 26128 264
rect 4802 226 4816 240
rect 19082 226 19096 240
rect 4322 202 4336 216
rect 9866 202 9880 216
rect 10298 202 10312 216
rect 19466 202 19480 216
rect 3890 178 3904 192
rect 6722 178 6736 192
rect 6962 178 6976 192
rect 17138 178 17152 192
rect 2762 154 2776 168
rect 16106 154 16120 168
rect 16346 154 16360 168
rect 19562 154 19576 168
rect 2738 130 2752 144
rect 11834 130 11848 144
rect 12602 130 12616 144
rect 22802 130 22816 144
rect 24314 130 24328 144
rect 2570 106 2584 120
rect 8306 106 8320 120
rect 8714 106 8728 120
rect 14018 106 14032 120
rect 15122 106 15136 120
rect 19634 106 19648 120
rect 70 82 84 96
rect 13010 82 13024 96
rect 13106 82 13120 96
rect 24026 82 24040 96
rect 26090 82 26104 96
rect 26451 82 26465 96
rect 70 58 84 72
rect 1730 58 1744 72
rect 2402 58 2416 72
rect 10946 58 10960 72
rect 19514 58 19528 72
rect 26090 58 26104 72
rect 26451 58 26465 72
rect 9794 34 9808 48
rect 26090 34 26104 48
rect 26114 34 26128 48
rect 26451 34 26465 48
rect 17042 10 17056 24
rect 26066 10 26080 24
rect 26451 10 26465 24
<< metal2 >>
rect 0 7773 70 7785
rect 0 7749 70 7761
rect 123 7666 323 7988
rect 339 7666 351 7988
rect 363 7666 375 7988
rect 387 7666 399 7988
rect 411 7666 423 7988
rect 2379 7786 2391 7988
rect 1731 7666 1743 7772
rect 2571 7666 2583 7796
rect 3195 7738 3207 7988
rect 3723 7666 3735 7820
rect 4011 7714 4023 7988
rect 4731 7666 4743 7844
rect 4827 7690 4839 7988
rect 5415 7882 5427 7988
rect 5416 7868 5434 7882
rect 5403 7666 5415 7868
rect 5919 7714 5931 7988
rect 7275 7882 7287 7988
rect 5920 7700 5938 7714
rect 5763 7666 5775 7676
rect 5787 7666 5799 7700
rect 5907 7666 5919 7700
rect 6003 7666 6015 7724
rect 6099 7666 6111 7772
rect 6723 7666 6735 7772
rect 7707 7666 7719 7724
rect 7995 7666 8007 7700
rect 8079 7690 8091 7988
rect 8907 7690 8919 7988
rect 9543 7978 9555 7988
rect 9544 7964 9562 7978
rect 8080 7676 8098 7690
rect 8067 7666 8079 7676
rect 9147 7666 9159 7892
rect 9267 7666 9279 7916
rect 9483 7666 9495 7940
rect 9531 7666 9543 7964
rect 10383 7882 10395 7988
rect 10384 7868 10402 7882
rect 10059 7666 10071 7868
rect 10371 7666 10383 7868
rect 10575 7714 10587 7988
rect 11391 7810 11403 7988
rect 12207 7954 12219 7988
rect 13803 7882 13815 7988
rect 13827 7906 13839 7988
rect 11163 7666 11175 7748
rect 12027 7666 12039 7796
rect 12603 7666 12615 7796
rect 12651 7666 12663 7748
rect 12987 7666 12999 7676
rect 14139 7666 14151 7700
rect 14331 7666 14343 7868
rect 14631 7858 14643 7988
rect 16215 7858 16227 7988
rect 17019 7882 17031 7988
rect 17823 7906 17835 7988
rect 16851 7666 16863 7796
rect 17847 7738 17859 7988
rect 19431 7906 19443 7988
rect 17715 7666 17727 7676
rect 17883 7666 17895 7892
rect 19455 7834 19467 7988
rect 19131 7666 19143 7724
rect 20259 7690 20271 7988
rect 21063 7930 21075 7988
rect 22647 7882 22659 7988
rect 21891 7666 21903 7868
rect 22155 7666 22167 7820
rect 22671 7762 22683 7988
rect 23355 7666 23367 7892
rect 23475 7834 23487 7988
rect 24003 7666 24015 7820
rect 24279 7714 24291 7988
rect 24411 7666 24423 7844
rect 24483 7666 24495 7868
rect 25695 7762 25707 7988
rect 26211 7914 26412 7988
rect 25779 7786 25791 7796
rect 25696 7748 25714 7762
rect 25683 7666 25695 7748
rect 25731 7666 25743 7748
rect 25755 7690 25767 7772
rect 25779 7714 25791 7748
rect 25803 7738 25815 7748
rect 25827 7738 25839 7820
rect 26211 7666 26411 7914
rect 26465 7773 26535 7785
rect 26465 7749 26535 7761
rect 26465 7725 26535 7737
rect 26465 7701 26535 7713
rect 26465 7677 26535 7689
rect 0 3820 70 3832
rect 0 3796 70 3808
rect 123 1697 323 6867
rect 339 1697 351 6867
rect 363 1697 375 6867
rect 387 1697 399 6867
rect 411 1697 423 6867
rect 1611 3785 1623 6867
rect 1611 1697 1623 3747
rect 1635 1697 1647 3723
rect 1659 3713 1671 6867
rect 1683 1697 1695 3675
rect 1731 3665 1743 6867
rect 1731 1697 1743 3627
rect 1779 3617 1791 6867
rect 1803 3857 1815 6867
rect 1827 3881 1839 6867
rect 1875 3929 1887 6867
rect 1899 3953 1911 6867
rect 1923 3977 1935 6867
rect 1971 4001 1983 6867
rect 1851 1697 1863 3891
rect 1995 3593 2007 6867
rect 2043 4025 2055 6867
rect 2091 4049 2103 6867
rect 2115 4073 2127 6867
rect 2139 3569 2151 6867
rect 2187 4097 2199 6867
rect 2211 3857 2223 6867
rect 2235 4121 2247 6867
rect 2235 3545 2247 3939
rect 2211 1697 2223 3531
rect 2259 1697 2271 3843
rect 2283 3545 2295 6867
rect 2307 4145 2319 6867
rect 2331 4169 2343 6867
rect 2355 3521 2367 6867
rect 2403 4193 2415 6867
rect 2451 4217 2463 6867
rect 2523 4241 2535 6867
rect 2547 4289 2559 6867
rect 2427 1697 2439 3699
rect 2451 1697 2463 3483
rect 2475 1697 2487 3699
rect 2523 1697 2535 3459
rect 2547 1697 2559 4251
rect 2595 1697 2607 4299
rect 2619 3449 2631 6867
rect 2643 4337 2655 6867
rect 2667 4361 2679 6867
rect 2715 4409 2727 6867
rect 2739 4433 2751 6867
rect 2643 1697 2655 3411
rect 2667 1697 2679 3387
rect 2691 1697 2703 4371
rect 2763 3377 2775 6867
rect 2787 4457 2799 6867
rect 2811 1697 2823 3339
rect 2835 3329 2847 6867
rect 2859 4481 2871 6867
rect 2883 4505 2895 6867
rect 2931 4529 2943 6867
rect 2955 4553 2967 6867
rect 3003 4577 3015 6867
rect 3051 4625 3063 6867
rect 2859 1697 2871 3291
rect 2883 1697 2895 3267
rect 2931 1697 2943 3243
rect 3051 1697 3063 4587
rect 3075 3761 3087 6867
rect 3099 4649 3111 6867
rect 3123 3233 3135 6867
rect 3171 4673 3183 6867
rect 3219 4697 3231 6867
rect 3291 4721 3303 6867
rect 3315 4745 3327 6867
rect 3339 3209 3351 6867
rect 3387 4769 3399 6867
rect 3411 4793 3423 6867
rect 3435 3545 3447 6867
rect 3459 4817 3471 6867
rect 3507 4841 3519 6867
rect 3555 4865 3567 6867
rect 3627 4889 3639 6867
rect 3651 4913 3663 6867
rect 3675 4937 3687 6867
rect 3411 1697 3423 3171
rect 3459 1697 3471 3987
rect 3603 1697 3615 4731
rect 3699 4217 3711 6867
rect 3771 4577 3783 6867
rect 3795 4961 3807 6867
rect 3651 1697 3663 3147
rect 3723 1697 3735 3123
rect 3747 1697 3759 4203
rect 3819 4073 3831 6867
rect 3867 4985 3879 6867
rect 3891 5009 3903 6867
rect 3915 5033 3927 6867
rect 3963 5057 3975 6867
rect 3771 1697 3783 3099
rect 3819 1697 3831 3075
rect 3843 1697 3855 3051
rect 3867 1697 3879 3027
rect 3939 1697 3951 3003
rect 3963 1697 3975 2979
rect 3987 2969 3999 6867
rect 4011 5081 4023 6867
rect 4059 5105 4071 6867
rect 4083 5129 4095 6867
rect 4107 5153 4119 6867
rect 4155 5177 4167 6867
rect 4011 1697 4023 2931
rect 4059 1697 4071 4515
rect 4083 1697 4095 3843
rect 4107 3041 4119 5115
rect 4107 1697 4119 2907
rect 4155 1697 4167 5115
rect 4179 3545 4191 6867
rect 4203 5201 4215 6867
rect 4251 5225 4263 6867
rect 4275 4673 4287 6867
rect 4299 5249 4311 6867
rect 4347 3689 4359 6867
rect 4371 5273 4383 6867
rect 4419 5297 4431 6867
rect 4467 4097 4479 6867
rect 4491 4001 4503 6867
rect 4515 5321 4527 6867
rect 4203 1697 4215 2883
rect 4275 1697 4287 2859
rect 4299 1697 4311 3147
rect 4371 1697 4383 2835
rect 4395 1697 4407 2811
rect 4443 1697 4455 2787
rect 4515 2777 4527 4131
rect 4563 3977 4575 6867
rect 4587 2777 4599 6867
rect 4611 3977 4623 6867
rect 4635 5369 4647 6867
rect 4683 5393 4695 6867
rect 4803 5417 4815 6867
rect 4491 1697 4503 2763
rect 4515 1697 4527 2739
rect 4539 1697 4551 2715
rect 4587 1697 4599 2691
rect 4611 1697 4623 3939
rect 4635 1697 4647 5331
rect 4683 1697 4695 2835
rect 4707 1697 4719 2667
rect 4755 1697 4767 4947
rect 4827 3953 4839 6867
rect 4851 2681 4863 6867
rect 4875 5465 4887 6867
rect 4923 5489 4935 6867
rect 4827 1697 4839 2643
rect 4875 1697 4887 5427
rect 4947 3857 4959 6867
rect 4995 5513 5007 6867
rect 5043 4577 5055 6867
rect 5067 4625 5079 6867
rect 5115 5537 5127 6867
rect 5163 5561 5175 6867
rect 5187 5585 5199 6867
rect 4923 1697 4935 3171
rect 4947 1697 4959 3267
rect 5043 1697 5055 2619
rect 5115 1697 5127 4179
rect 5139 1697 5151 3939
rect 5211 2897 5223 6867
rect 5235 2609 5247 6867
rect 5283 5633 5295 6867
rect 5283 1697 5295 5595
rect 5307 2849 5319 6867
rect 5355 5657 5367 6867
rect 5403 3737 5415 6867
rect 5451 3857 5463 6867
rect 5475 4577 5487 6867
rect 5499 2801 5511 6867
rect 5523 5681 5535 6867
rect 5571 2585 5583 6867
rect 5595 3137 5607 6867
rect 5619 5705 5631 6867
rect 5667 5729 5679 6867
rect 5691 2993 5703 6867
rect 5691 1697 5703 2547
rect 5715 2537 5727 6867
rect 5763 2825 5775 6867
rect 5787 5753 5799 6867
rect 5811 5777 5823 6867
rect 5835 1697 5847 5091
rect 5859 2873 5871 6867
rect 5883 3065 5895 6867
rect 5907 4745 5919 6867
rect 5931 5801 5943 6867
rect 5931 1697 5943 5091
rect 5979 5057 5991 6867
rect 6003 5825 6015 6867
rect 6027 5849 6039 6867
rect 6099 5873 6111 6867
rect 6123 5825 6135 6867
rect 6171 5921 6183 6867
rect 6195 5945 6207 6867
rect 5955 1697 5967 2811
rect 6027 1697 6039 5523
rect 6051 1697 6063 3531
rect 6099 1697 6111 2499
rect 6147 1697 6159 5883
rect 6171 1697 6183 4131
rect 6219 1697 6231 4659
rect 6267 3137 6279 6867
rect 6291 5921 6303 6867
rect 6315 5873 6327 6867
rect 6243 1697 6255 2475
rect 6291 1697 6303 4755
rect 6315 1697 6327 3939
rect 6339 2465 6351 6867
rect 6387 5969 6399 6867
rect 6411 5777 6423 6867
rect 6435 5993 6447 6867
rect 6363 1697 6375 4131
rect 6411 1697 6423 5163
rect 6435 1697 6447 5235
rect 6459 1697 6471 6003
rect 6483 3545 6495 6867
rect 6507 3761 6519 6867
rect 6531 5561 6543 6867
rect 6555 6041 6567 6867
rect 6603 3257 6615 6867
rect 6627 4529 6639 6867
rect 6651 6065 6663 6867
rect 6699 6089 6711 6867
rect 6507 1697 6519 2883
rect 6531 1697 6543 2427
rect 6555 1697 6567 2955
rect 6603 1697 6615 2955
rect 6627 1697 6639 3843
rect 6651 1697 6663 5619
rect 6675 2969 6687 4563
rect 6747 4265 6759 6867
rect 6795 4265 6807 6867
rect 6699 1697 6711 2403
rect 6747 1697 6759 3195
rect 6771 1697 6783 2955
rect 6795 1697 6807 3771
rect 6819 3209 6831 6867
rect 6843 3833 6855 6867
rect 6867 6113 6879 6867
rect 6915 5873 6927 6867
rect 6843 1697 6855 3771
rect 6867 2993 6879 4251
rect 6891 3785 6903 5259
rect 6963 4265 6975 6867
rect 6987 1697 6999 5139
rect 7011 1697 7023 3147
rect 7035 3137 7047 6867
rect 7059 3785 7071 6867
rect 7035 1697 7047 2379
rect 7083 2369 7095 6867
rect 7131 4001 7143 6867
rect 7155 3137 7167 6867
rect 7179 6137 7191 6867
rect 7227 4481 7239 6867
rect 7251 4625 7263 6867
rect 7275 4241 7287 6867
rect 7323 3761 7335 6867
rect 7347 4961 7359 6867
rect 7371 6161 7383 6867
rect 7083 1697 7095 2331
rect 7179 1697 7191 2307
rect 7275 1697 7287 2283
rect 7323 1697 7335 2259
rect 7371 1697 7383 5043
rect 7419 3689 7431 6867
rect 7395 1697 7407 3267
rect 7443 3089 7455 6867
rect 7491 6185 7503 6867
rect 7443 1697 7455 2307
rect 7491 1697 7503 5835
rect 7515 1697 7527 6195
rect 7539 2489 7551 6867
rect 7563 5849 7575 6867
rect 7587 4409 7599 6867
rect 7635 6233 7647 6867
rect 7539 1697 7551 2451
rect 7563 1697 7575 2235
rect 7611 1697 7623 5571
rect 7659 5561 7671 6867
rect 7635 1697 7647 4731
rect 7707 4409 7719 6867
rect 7755 6257 7767 6867
rect 7779 5249 7791 6867
rect 7803 6281 7815 6867
rect 7851 5177 7863 6867
rect 7659 1697 7671 2451
rect 7707 1697 7719 2211
rect 7779 1697 7791 2187
rect 7851 1697 7863 5139
rect 7875 3857 7887 6867
rect 7899 3401 7911 6867
rect 7875 1697 7887 2163
rect 7923 1697 7935 6075
rect 7947 4241 7959 6867
rect 7947 1697 7959 2139
rect 7971 1697 7983 6291
rect 8019 1697 8031 5739
rect 8067 3041 8079 6867
rect 8091 5753 8103 6867
rect 8139 6329 8151 6867
rect 8187 4577 8199 6867
rect 8211 6353 8223 6867
rect 8235 6377 8247 6867
rect 8067 1697 8079 2979
rect 8139 1697 8151 4563
rect 8163 1697 8175 4227
rect 8211 1697 8223 5955
rect 8235 2393 8247 6339
rect 8283 4097 8295 6867
rect 8307 3305 8319 6867
rect 8331 6353 8343 6867
rect 8379 6401 8391 6867
rect 8259 1697 8271 2931
rect 8355 1697 8367 5139
rect 8403 2897 8415 6867
rect 8427 4673 8439 6867
rect 8475 5057 8487 6867
rect 8499 6425 8511 6867
rect 8523 5897 8535 6867
rect 8571 5945 8583 6867
rect 8379 1697 8391 2883
rect 8451 1697 8463 4971
rect 8499 1697 8511 4659
rect 8571 1697 8583 3723
rect 8595 2825 8607 6867
rect 8619 5897 8631 6867
rect 8667 6449 8679 6867
rect 8619 1697 8631 2379
rect 8691 2129 8703 6867
rect 8739 2105 8751 6867
rect 8787 2177 8799 6867
rect 8811 4745 8823 6867
rect 8835 2345 8847 6867
rect 8883 2345 8895 6867
rect 8907 6473 8919 6867
rect 8931 6497 8943 6867
rect 8763 1697 8775 2067
rect 8811 1697 8823 2043
rect 8859 1697 8871 2163
rect 8907 1697 8919 4515
rect 8931 1697 8943 5403
rect 8979 2321 8991 6867
rect 9003 4265 9015 6867
rect 9027 6209 9039 6867
rect 9075 6209 9087 6867
rect 9099 6521 9111 6867
rect 9123 5393 9135 6867
rect 9195 6545 9207 6867
rect 8955 1697 8967 2019
rect 9003 1697 9015 1995
rect 9027 1697 9039 4179
rect 9075 1697 9087 1971
rect 9123 1697 9135 5235
rect 9147 1697 9159 3747
rect 9171 1697 9183 5235
rect 9195 1697 9207 3483
rect 9219 1985 9231 6867
rect 9243 3497 9255 6867
rect 9315 6497 9327 6867
rect 9267 1697 9279 6483
rect 9291 1697 9303 2595
rect 9339 2081 9351 6867
rect 9363 5081 9375 6867
rect 9387 6569 9399 6867
rect 9435 6521 9447 6867
rect 9459 5081 9471 6867
rect 9531 6593 9543 6867
rect 9315 1697 9327 1971
rect 9387 1697 9399 4683
rect 9411 1697 9423 2595
rect 9435 1697 9447 2667
rect 9459 1697 9471 1947
rect 9507 1697 9519 5115
rect 9531 1697 9543 3747
rect 9555 1697 9567 6387
rect 9579 3641 9591 6867
rect 9627 6617 9639 6867
rect 9627 1697 9639 3939
rect 9651 1697 9663 6459
rect 9699 6233 9711 6867
rect 9747 4481 9759 6867
rect 9819 6017 9831 6867
rect 9843 5801 9855 6867
rect 9867 6017 9879 6867
rect 9891 5801 9903 6867
rect 9675 1697 9687 3627
rect 9771 1697 9783 4875
rect 9843 1697 9855 1923
rect 9891 1697 9903 5451
rect 9915 2009 9927 6867
rect 9915 1697 9927 1899
rect 9939 1697 9951 2571
rect 9963 2273 9975 6867
rect 9987 3161 9999 6867
rect 10011 5465 10023 6867
rect 9987 1697 9999 2571
rect 10035 1697 10047 2259
rect 10059 2009 10071 6867
rect 10083 4745 10095 6867
rect 10107 1913 10119 6867
rect 10155 6281 10167 6867
rect 10203 3929 10215 6867
rect 10275 6353 10287 6867
rect 10131 1889 10143 1995
rect 10107 1697 10119 1875
rect 10155 1697 10167 3147
rect 10179 1697 10191 3723
rect 10227 1889 10239 4971
rect 10299 4001 10311 6867
rect 10323 4985 10335 6867
rect 10347 3929 10359 6531
rect 10203 1697 10215 1875
rect 10275 1697 10287 3915
rect 10371 3713 10383 6867
rect 10323 1697 10335 1875
rect 10347 1697 10359 1851
rect 10395 1697 10407 6243
rect 10419 4361 10431 6867
rect 10419 1697 10431 3267
rect 10443 3041 10455 6867
rect 10467 4361 10479 6867
rect 10515 4697 10527 6867
rect 10539 5105 10551 6867
rect 10491 1697 10503 2043
rect 10515 1697 10527 3915
rect 10563 2849 10575 6867
rect 10587 3929 10599 6387
rect 10611 4385 10623 6867
rect 10635 4241 10647 6867
rect 10659 4385 10671 6867
rect 10707 5513 10719 6867
rect 10731 5417 10743 6867
rect 10779 5513 10791 6867
rect 10563 1697 10575 1827
rect 10611 1697 10623 3747
rect 10635 1697 10647 2859
rect 10671 1841 10683 4227
rect 10827 3929 10839 6867
rect 10731 1697 10743 3843
rect 10827 1697 10839 3699
rect 10851 2993 10863 6867
rect 10899 5561 10911 6867
rect 10875 1697 10887 3939
rect 10899 1697 10911 5163
rect 10923 1697 10935 4683
rect 10947 4553 10959 6867
rect 10971 3353 10983 6867
rect 11019 4577 11031 6867
rect 11067 6641 11079 6867
rect 11091 6665 11103 6867
rect 11115 6689 11127 6867
rect 11139 3857 11151 6867
rect 11043 1697 11055 1827
rect 11091 1697 11103 3315
rect 11139 1697 11151 3027
rect 11187 1697 11199 6387
rect 11211 4865 11223 6867
rect 11235 2057 11247 6867
rect 11259 5009 11271 6867
rect 11307 5009 11319 6867
rect 11331 3329 11343 6867
rect 11355 3161 11367 6867
rect 11379 6713 11391 6867
rect 11427 6497 11439 6867
rect 11475 4097 11487 6867
rect 11547 5465 11559 6867
rect 11571 1817 11583 6867
rect 11619 5465 11631 6867
rect 11667 2873 11679 6867
rect 11691 3761 11703 6867
rect 11715 3161 11727 6867
rect 11739 1793 11751 6867
rect 11787 2945 11799 6867
rect 11811 1769 11823 6867
rect 11835 6737 11847 6867
rect 11883 6425 11895 6867
rect 11931 2057 11943 6867
rect 11979 1697 11991 4779
rect 12003 2489 12015 6867
rect 12051 6785 12063 6867
rect 12003 1697 12015 1731
rect 12027 1697 12039 6747
rect 12075 1697 12087 3387
rect 12099 2897 12111 6867
rect 12123 3401 12135 6867
rect 12147 6425 12159 6867
rect 12195 5153 12207 6867
rect 12123 1697 12135 2595
rect 12159 2009 12171 3387
rect 12195 1697 12207 3387
rect 12219 1697 12231 3675
rect 12243 2873 12255 6867
rect 12315 6809 12327 6867
rect 12243 1697 12255 2667
rect 12267 1697 12279 6411
rect 12291 3401 12303 6387
rect 12339 5825 12351 6867
rect 12363 5921 12375 6867
rect 12315 1697 12327 3003
rect 12387 1697 12399 4875
rect 12411 2681 12423 6867
rect 12435 3041 12447 6867
rect 12459 4841 12471 6867
rect 12507 6833 12519 6867
rect 12531 6377 12543 6867
rect 12459 1697 12471 3387
rect 12483 1697 12495 5979
rect 12507 1697 12519 5187
rect 12531 1697 12543 3507
rect 12555 2705 12567 6867
rect 12579 2993 12591 6795
rect 12603 3401 12615 6147
rect 12555 1697 12567 1707
rect 12651 1697 12663 5715
rect 12723 5201 12735 6867
rect 12723 1697 12735 3723
rect 12747 3137 12759 6867
rect 12771 5993 12783 6867
rect 12747 1697 12759 3123
rect 12771 1697 12783 3027
rect 12795 2825 12807 6867
rect 12819 3425 12831 6867
rect 12843 2993 12855 5187
rect 12867 4169 12879 6867
rect 12915 5201 12927 6867
rect 12795 1697 12807 1803
rect 12867 1697 12879 4059
rect 12891 1697 12903 4803
rect 12987 3521 12999 6867
rect 13035 4961 13047 6867
rect 13083 6161 13095 6867
rect 13155 3857 13167 6867
rect 13179 4865 13191 6867
rect 13203 6377 13215 6867
rect 13251 6809 13263 6867
rect 12915 1697 12927 3507
rect 12987 1697 12999 3411
rect 13059 1697 13071 2739
rect 13083 1697 13095 3843
rect 13155 1697 13167 2547
rect 13179 1697 13191 3507
rect 13251 1697 13263 4107
rect 13275 3761 13287 6867
rect 13275 1697 13287 2907
rect 13299 2897 13311 6867
rect 13323 6857 13335 6867
rect 13323 1697 13335 6819
rect 13347 2873 13359 6795
rect 13371 3137 13383 6867
rect 13395 6809 13407 6867
rect 13395 1697 13407 5955
rect 13419 4121 13431 6867
rect 13419 1697 13431 1731
rect 13443 1697 13455 5067
rect 13467 2345 13479 6867
rect 13491 3305 13503 6867
rect 13515 5393 13527 6867
rect 13491 1697 13503 2883
rect 13515 1697 13527 3387
rect 13539 2897 13551 6267
rect 13563 4673 13575 6867
rect 13587 5201 13599 6867
rect 13611 5249 13623 6867
rect 13611 1697 13623 4539
rect 13731 4457 13743 6867
rect 13635 1697 13647 2667
rect 13707 1697 13719 2883
rect 13731 1697 13743 4347
rect 13827 1697 13839 6075
rect 13947 1697 13959 3939
rect 13971 1697 13983 6315
rect 14091 4673 14103 6867
rect 14139 5849 14151 6867
rect 14067 1697 14079 3291
rect 14091 1697 14103 4515
rect 14151 3521 14163 4659
rect 14115 1697 14127 3339
rect 14187 1697 14199 5643
rect 14283 4505 14295 6867
rect 14307 5393 14319 6867
rect 14211 1697 14223 1731
rect 14235 1697 14247 4275
rect 14307 1697 14319 4275
rect 14331 1697 14343 3939
rect 14355 1697 14367 4875
rect 14379 4289 14391 6411
rect 14451 4361 14463 6867
rect 14427 1697 14439 4275
rect 14451 1697 14463 3507
rect 14475 1697 14487 5739
rect 14547 1697 14559 6243
rect 14571 1697 14583 3123
rect 14619 1697 14631 5163
rect 14667 1697 14679 5811
rect 14691 1697 14703 5859
rect 14811 5057 14823 6867
rect 14739 1697 14751 4155
rect 14787 1697 14799 3051
rect 14811 1697 14823 3075
rect 14859 2753 14871 6867
rect 14883 1697 14895 4731
rect 15003 4481 15015 6867
rect 15027 4457 15039 6867
rect 15051 6521 15063 6867
rect 14907 1697 14919 2811
rect 15003 1697 15015 2691
rect 15075 1697 15087 6147
rect 15099 2753 15111 6867
rect 15123 5033 15135 6867
rect 15147 4481 15159 6867
rect 15099 1697 15111 1803
rect 15171 1697 15183 5307
rect 15195 4697 15207 6867
rect 15219 6257 15231 6867
rect 15243 4673 15255 6867
rect 15195 1697 15207 4491
rect 15243 1697 15255 4179
rect 15267 3977 15279 6867
rect 15315 5321 15327 6867
rect 15339 5081 15351 6867
rect 15363 5201 15375 6867
rect 15387 5249 15399 6867
rect 15291 1697 15303 4179
rect 15315 1697 15327 2307
rect 15387 1697 15399 4611
rect 15411 3809 15423 6867
rect 15411 1697 15423 3747
rect 15435 1697 15447 3531
rect 15459 2249 15471 6867
rect 15483 3041 15495 6867
rect 15507 5969 15519 6867
rect 15531 4505 15543 6459
rect 15555 4841 15567 6867
rect 15579 5153 15591 6867
rect 15603 4217 15615 6867
rect 15651 5033 15663 6867
rect 15507 1697 15519 4059
rect 15555 1697 15567 3195
rect 15627 2681 15639 4659
rect 15675 3401 15687 5235
rect 15699 4505 15711 6867
rect 15771 2465 15783 6867
rect 15795 6113 15807 6867
rect 15819 4673 15831 6867
rect 15843 5681 15855 6867
rect 15867 4841 15879 6867
rect 15915 2729 15927 6867
rect 15963 3761 15975 6867
rect 16035 2297 16047 6867
rect 16059 3113 16071 6867
rect 16107 6689 16119 6867
rect 16155 2081 16167 6867
rect 16179 6497 16191 6867
rect 16203 5033 16215 6867
rect 16251 5417 16263 6867
rect 16275 3281 16287 6867
rect 16251 1697 16263 3027
rect 16275 1697 16287 2811
rect 16299 1697 16311 5259
rect 16323 4553 16335 6867
rect 16443 5249 16455 6867
rect 16371 1697 16383 2811
rect 16443 1697 16455 2739
rect 16467 1697 16479 2619
rect 16491 1697 16503 3291
rect 16515 1697 16527 2355
rect 16611 1697 16623 5499
rect 16731 1697 16743 4155
rect 16779 1697 16791 4203
rect 16827 1697 16839 5283
rect 16995 4721 17007 6867
rect 16851 1697 16863 3147
rect 16947 1697 16959 4611
rect 16995 1697 17007 3315
rect 17019 3161 17031 6867
rect 17043 5513 17055 6867
rect 17091 3305 17103 6867
rect 17115 4529 17127 6867
rect 17043 1697 17055 1755
rect 17091 1697 17103 3195
rect 17115 1697 17127 3723
rect 17139 2801 17151 6867
rect 17163 1985 17175 6867
rect 17187 1697 17199 6123
rect 17211 5057 17223 6867
rect 17211 1697 17223 5043
rect 17235 3185 17247 6867
rect 17259 1697 17271 6651
rect 17283 4529 17295 6867
rect 17307 1697 17319 3123
rect 17331 2945 17343 6867
rect 17355 3713 17367 6867
rect 17379 5681 17391 6867
rect 17427 3545 17439 6867
rect 17451 4169 17463 6867
rect 17331 1697 17343 2451
rect 17355 1697 17367 3315
rect 17403 1697 17415 1803
rect 17427 1697 17439 3123
rect 17451 1697 17463 2835
rect 17475 1817 17487 6867
rect 17499 3209 17511 5259
rect 17523 3161 17535 6867
rect 17547 5273 17559 6867
rect 17571 5129 17583 6867
rect 17619 6545 17631 6867
rect 17475 1697 17487 1755
rect 17523 1697 17535 2715
rect 17547 1697 17559 3723
rect 17595 1697 17607 3051
rect 17643 1961 17655 6867
rect 17667 4385 17679 6867
rect 17667 1697 17679 4059
rect 17691 3497 17703 6867
rect 17715 1697 17727 4659
rect 17739 2465 17751 5115
rect 17763 4385 17775 6867
rect 17787 3881 17799 6867
rect 17763 1697 17775 2739
rect 17787 1697 17799 3795
rect 17811 3401 17823 6867
rect 17835 3905 17847 6867
rect 17859 3329 17871 6627
rect 17883 4673 17895 6867
rect 17883 1697 17895 4443
rect 17931 4217 17943 6867
rect 17955 6113 17967 6867
rect 17907 1697 17919 3531
rect 17931 1697 17943 3771
rect 17979 1697 17991 5355
rect 18003 1841 18015 6867
rect 18027 1697 18039 5187
rect 18051 3641 18063 6867
rect 18075 3137 18087 6867
rect 18099 5201 18111 6867
rect 18147 4841 18159 6867
rect 18099 1697 18111 3675
rect 18123 1697 18135 4203
rect 18171 2585 18183 6867
rect 18219 3953 18231 6867
rect 18195 1697 18207 3675
rect 18243 1697 18255 3963
rect 18267 2753 18279 6867
rect 18291 3257 18303 6867
rect 18315 4001 18327 6867
rect 18339 4889 18351 6867
rect 18291 1697 18303 3195
rect 18315 1697 18327 3939
rect 18351 2033 18363 4371
rect 18387 2609 18399 6867
rect 18411 4697 18423 6867
rect 18435 4913 18447 6867
rect 18459 1697 18471 6603
rect 18483 2177 18495 6867
rect 18507 2393 18519 5259
rect 18531 3545 18543 6867
rect 18603 4553 18615 6867
rect 18555 3209 18567 4467
rect 18579 3953 18591 4011
rect 18627 3185 18639 6867
rect 18675 4769 18687 6867
rect 18723 5153 18735 6867
rect 18747 3161 18759 6867
rect 18771 4385 18783 6867
rect 18819 6569 18831 6867
rect 18843 6473 18855 6867
rect 18867 4481 18879 6867
rect 18915 3761 18927 6867
rect 18939 4385 18951 6867
rect 18963 2657 18975 6867
rect 19011 6401 19023 6867
rect 19011 1697 19023 5547
rect 19035 4745 19047 6867
rect 19035 1697 19047 3051
rect 19059 1937 19071 6867
rect 19107 6089 19119 6867
rect 19131 1697 19143 5187
rect 19155 4433 19167 6867
rect 19203 6185 19215 6867
rect 19179 1697 19191 6051
rect 19203 1697 19215 6123
rect 19227 4865 19239 6867
rect 19251 6233 19263 6867
rect 19299 6065 19311 6867
rect 19275 1697 19287 4275
rect 19299 1697 19311 5739
rect 19323 4385 19335 6867
rect 19347 6737 19359 6867
rect 19347 1697 19359 6099
rect 19371 5609 19383 6867
rect 19419 4433 19431 6867
rect 19443 6545 19455 6867
rect 19467 2273 19479 6867
rect 19491 4769 19503 6867
rect 19539 5537 19551 6867
rect 19563 4649 19575 6867
rect 19587 2777 19599 6867
rect 19611 1697 19623 4131
rect 19635 3185 19647 6867
rect 19659 4841 19671 6867
rect 19683 4865 19695 6867
rect 19731 5777 19743 6867
rect 19659 1697 19671 1875
rect 19707 1697 19719 2019
rect 19755 1697 19767 6243
rect 19779 1745 19791 6867
rect 19851 3065 19863 6867
rect 19875 6713 19887 6867
rect 19923 4073 19935 6867
rect 19971 5921 19983 6867
rect 19827 1697 19839 2811
rect 19875 1697 19887 2667
rect 19947 1697 19959 4563
rect 19971 1697 19983 5043
rect 19995 4265 20007 6867
rect 20019 4073 20031 6819
rect 20043 4625 20055 6867
rect 20091 4265 20103 6867
rect 20115 5825 20127 6867
rect 20163 5729 20175 6867
rect 19995 1697 20007 4059
rect 20043 1697 20055 3171
rect 20067 1697 20079 3267
rect 20115 1697 20127 5475
rect 20163 1697 20175 4059
rect 20187 1697 20199 3267
rect 20235 1697 20247 6579
rect 20283 4313 20295 6867
rect 20283 1697 20295 4227
rect 20307 1697 20319 3123
rect 20331 1697 20343 4515
rect 20355 1697 20367 5763
rect 20379 1697 20391 5787
rect 20427 1697 20439 1899
rect 20475 1697 20487 3075
rect 20547 1697 20559 5163
rect 20571 1697 20583 3987
rect 20643 3521 20655 6867
rect 20691 4313 20703 6867
rect 20643 1697 20655 2931
rect 20691 1697 20703 3363
rect 20739 1697 20751 6651
rect 20763 1697 20775 4851
rect 20835 3833 20847 6867
rect 20883 4841 20895 6867
rect 20955 5321 20967 6867
rect 20787 1697 20799 3603
rect 20835 1697 20847 3339
rect 20907 1697 20919 3579
rect 20979 1697 20991 4539
rect 21003 2345 21015 6867
rect 21075 5345 21087 6867
rect 21099 4985 21111 6867
rect 21075 1697 21087 3939
rect 21099 1697 21111 4875
rect 21123 4601 21135 6867
rect 21147 3953 21159 6027
rect 21171 4145 21183 6867
rect 21195 4793 21207 6867
rect 21171 1697 21183 3891
rect 21195 1697 21207 3939
rect 21219 3905 21231 5283
rect 21243 4577 21255 6867
rect 21243 1697 21255 3867
rect 21291 2921 21303 6867
rect 21339 5993 21351 6867
rect 21411 6401 21423 6867
rect 21435 4601 21447 6867
rect 21339 1697 21351 3891
rect 21363 1697 21375 3819
rect 21387 1697 21399 4347
rect 21435 1697 21447 4395
rect 21459 3809 21471 6867
rect 21483 1697 21495 6003
rect 21507 2801 21519 6867
rect 21555 6809 21567 6867
rect 21531 2009 21543 4587
rect 21555 1697 21567 5859
rect 21579 1697 21591 5811
rect 21627 2057 21639 6867
rect 21651 2825 21663 6867
rect 21675 5225 21687 6867
rect 21723 6185 21735 6867
rect 21747 5273 21759 6867
rect 21675 1697 21687 3915
rect 21747 1697 21759 5211
rect 21771 2417 21783 6867
rect 21819 5657 21831 6867
rect 21843 5777 21855 6867
rect 21795 1697 21807 4635
rect 21867 1697 21879 2475
rect 21891 1697 21903 2547
rect 21915 1697 21927 6051
rect 21939 4025 21951 6867
rect 21963 5153 21975 6867
rect 21963 1697 21975 5043
rect 21987 4193 21999 6867
rect 21987 1697 21999 3267
rect 22011 1697 22023 6483
rect 22035 5993 22047 6867
rect 22059 6473 22071 6867
rect 22083 1697 22095 5019
rect 22107 4073 22119 6867
rect 22131 4505 22143 5139
rect 22155 2561 22167 6867
rect 22203 4241 22215 6867
rect 22227 3761 22239 6867
rect 22179 1697 22191 3747
rect 22251 2825 22263 6867
rect 22275 4433 22287 6867
rect 22323 6761 22335 6867
rect 22251 1697 22263 2787
rect 22299 1697 22311 2523
rect 22323 1697 22335 2667
rect 22347 2057 22359 6867
rect 22371 2897 22383 6867
rect 22347 1697 22359 2019
rect 22395 1697 22407 5859
rect 22419 3257 22431 6867
rect 22419 1697 22431 3195
rect 22443 3185 22455 6867
rect 22467 3905 22479 6867
rect 22443 1697 22455 3147
rect 22491 2801 22503 5571
rect 22515 4097 22527 6867
rect 22539 5417 22551 6867
rect 22539 1697 22551 3843
rect 22563 3401 22575 6867
rect 22611 4529 22623 6867
rect 22587 1697 22599 3651
rect 22635 1769 22647 6867
rect 22659 3425 22671 6867
rect 22683 1697 22695 6339
rect 22707 3641 22719 6867
rect 22707 1697 22719 3603
rect 22731 2033 22743 5259
rect 22755 3305 22767 6867
rect 22755 1697 22767 3243
rect 22779 3209 22791 4299
rect 22803 3161 22815 5811
rect 22827 2393 22839 6867
rect 22851 5105 22863 6867
rect 22875 4745 22887 6867
rect 22899 4337 22911 6867
rect 22923 3617 22935 4659
rect 22947 4073 22959 6867
rect 22971 6017 22983 6867
rect 22971 1697 22983 5907
rect 22995 4049 23007 6867
rect 23043 5945 23055 6867
rect 22995 1697 23007 4011
rect 23019 3257 23031 5835
rect 23067 4553 23079 6867
rect 23043 1697 23055 4443
rect 23091 4337 23103 6867
rect 23115 4361 23127 6867
rect 23163 4337 23175 6867
rect 23091 1697 23103 3267
rect 23127 3041 23139 4323
rect 23115 1697 23127 2811
rect 23187 2753 23199 6867
rect 23163 1697 23175 2115
rect 23211 1697 23223 5883
rect 23235 2585 23247 6867
rect 23283 6857 23295 6867
rect 23235 1697 23247 2043
rect 23259 1769 23271 6003
rect 23307 5513 23319 6867
rect 23331 3977 23343 6867
rect 23307 1697 23319 3531
rect 23331 1697 23343 3915
rect 23355 1697 23367 2979
rect 23379 1697 23391 6195
rect 23403 5057 23415 6867
rect 23427 4169 23439 6867
rect 23475 4793 23487 6867
rect 23523 6425 23535 6867
rect 23487 2297 23499 4347
rect 23451 1697 23463 1779
rect 23523 1697 23535 6075
rect 23547 4025 23559 5859
rect 23571 4721 23583 6867
rect 23571 1697 23583 2811
rect 23595 1697 23607 6387
rect 23643 6161 23655 6867
rect 23619 1697 23631 1995
rect 23643 1697 23655 4995
rect 23667 2177 23679 6867
rect 23691 4001 23703 6867
rect 23691 1697 23703 3219
rect 23715 1697 23727 4875
rect 23739 2705 23751 6867
rect 23763 6569 23775 6867
rect 23763 1697 23775 6531
rect 23787 4217 23799 6867
rect 23835 4361 23847 6867
rect 23859 4481 23871 6867
rect 23883 5705 23895 6867
rect 23907 6377 23919 6867
rect 23931 4553 23943 6867
rect 23979 6089 23991 6867
rect 23811 1697 23823 3627
rect 23835 1697 23847 2739
rect 23859 1697 23871 3819
rect 23907 1697 23919 3123
rect 23931 1697 23943 4515
rect 23955 1697 23967 4227
rect 23979 1697 23991 5067
rect 24027 4385 24039 6867
rect 24075 4817 24087 6867
rect 24099 5753 24111 6867
rect 24003 1889 24015 4323
rect 24051 1697 24063 2091
rect 24075 1697 24087 4227
rect 24099 1697 24111 4203
rect 24123 3929 24135 4563
rect 24147 3953 24159 6867
rect 24195 4265 24207 6867
rect 24219 5825 24231 6867
rect 24267 4289 24279 6867
rect 24171 1697 24183 3723
rect 24195 1697 24207 2691
rect 24219 1697 24231 1995
rect 24243 1697 24255 3435
rect 24291 2009 24303 6555
rect 24315 5393 24327 6867
rect 24339 3881 24351 6867
rect 24363 5441 24375 6867
rect 24387 5633 24399 6867
rect 24387 1697 24399 3747
rect 24411 1697 24423 4683
rect 24435 2225 24447 4539
rect 24459 2489 24471 6867
rect 24483 6017 24495 6867
rect 24483 1697 24495 5979
rect 24507 3473 24519 6867
rect 24531 4241 24543 5955
rect 24555 5417 24567 6867
rect 24531 3449 24543 4107
rect 24507 1697 24519 3435
rect 24579 3137 24591 6867
rect 24603 5129 24615 6867
rect 24627 4361 24639 6867
rect 24651 4313 24663 6003
rect 24675 5057 24687 6867
rect 24699 2873 24711 6867
rect 24723 4217 24735 6867
rect 24771 3041 24783 6867
rect 24795 5873 24807 6867
rect 24819 2441 24831 6867
rect 24867 6785 24879 6867
rect 24891 6305 24903 6867
rect 24915 5681 24927 6867
rect 24939 5249 24951 6867
rect 24987 3833 24999 6867
rect 25011 5465 25023 6867
rect 25011 1697 25023 3267
rect 25035 2201 25047 6867
rect 25059 4289 25071 6867
rect 25083 4313 25095 6867
rect 25131 4577 25143 6867
rect 25059 1697 25071 3123
rect 25095 2633 25107 4275
rect 25155 3545 25167 6867
rect 25179 3017 25191 6867
rect 25227 5033 25239 6867
rect 25203 1697 25215 3123
rect 25227 1697 25239 4995
rect 25251 1721 25263 5019
rect 25275 4937 25287 6867
rect 25299 1697 25311 6627
rect 25323 1697 25335 2619
rect 25347 2321 25359 6867
rect 25371 5105 25383 6867
rect 25419 6449 25431 6867
rect 25443 4289 25455 6459
rect 25371 1697 25383 4275
rect 25395 1697 25407 4251
rect 25467 4145 25479 6867
rect 25491 4961 25503 6867
rect 25515 2969 25527 6867
rect 25563 2009 25575 6867
rect 25611 5105 25623 6867
rect 25683 2513 25695 6867
rect 25731 2153 25743 6867
rect 25875 1697 25887 5403
rect 25923 1697 25935 6459
rect 26067 1697 26079 3555
rect 26091 1721 26103 4755
rect 26115 1745 26127 4251
rect 26211 1697 26411 6867
rect 26465 4300 26535 4312
rect 26465 1852 26535 1864
rect 26465 1732 26535 1744
rect 26465 1708 26535 1720
rect 0 83 70 95
rect 0 59 70 71
rect 123 0 323 898
rect 339 0 351 898
rect 363 0 375 898
rect 387 0 399 898
rect 411 0 423 898
rect 1731 72 1743 898
rect 2403 72 2415 898
rect 2571 120 2583 898
rect 2739 144 2751 898
rect 2763 168 2775 898
rect 3891 192 3903 898
rect 4323 216 4335 898
rect 4803 240 4815 898
rect 5163 264 5175 898
rect 5643 288 5655 898
rect 5859 312 5871 898
rect 5883 336 5895 898
rect 5979 360 5991 898
rect 6195 384 6207 898
rect 6723 192 6735 898
rect 6891 312 6903 898
rect 6963 192 6975 898
rect 7107 336 7119 898
rect 7131 408 7143 898
rect 7203 336 7215 898
rect 7227 432 7239 898
rect 7299 456 7311 898
rect 7731 504 7743 898
rect 7695 0 7707 466
rect 7827 360 7839 898
rect 8283 480 8295 898
rect 8307 120 8319 898
rect 8403 360 8415 898
rect 8475 480 8487 898
rect 8523 336 8535 898
rect 8691 336 8703 898
rect 8715 120 8727 898
rect 8835 312 8847 898
rect 9243 528 9255 898
rect 9339 552 9351 898
rect 9579 576 9591 898
rect 9723 600 9735 898
rect 9747 264 9759 898
rect 9795 48 9807 898
rect 9867 216 9879 898
rect 10131 312 10143 898
rect 10251 264 10263 898
rect 10299 216 10311 898
rect 10443 528 10455 898
rect 10659 528 10671 898
rect 10707 624 10719 898
rect 10779 504 10791 898
rect 10827 504 10839 898
rect 10840 490 10858 504
rect 10839 0 10851 490
rect 10947 72 10959 898
rect 10995 504 11007 898
rect 11019 648 11031 898
rect 11067 672 11079 898
rect 11259 696 11271 898
rect 11307 720 11319 898
rect 11835 144 11847 898
rect 12339 600 12351 898
rect 12363 264 12375 898
rect 12411 264 12423 898
rect 12603 144 12615 898
rect 12627 744 12639 898
rect 12675 672 12687 898
rect 12843 672 12855 898
rect 12963 768 12975 898
rect 13011 96 13023 898
rect 13107 96 13119 898
rect 13203 744 13215 898
rect 13299 792 13311 898
rect 13347 816 13359 898
rect 13563 768 13575 898
rect 13659 456 13671 898
rect 13779 384 13791 898
rect 13875 456 13887 898
rect 14019 120 14031 898
rect 14139 384 14151 898
rect 14283 528 14295 898
rect 14379 528 14391 898
rect 14499 504 14511 898
rect 14835 504 14847 898
rect 15123 120 15135 898
rect 15339 840 15351 898
rect 15459 600 15471 898
rect 15699 600 15711 898
rect 16107 168 16119 898
rect 16347 168 16359 898
rect 16395 864 16407 898
rect 16539 696 16551 898
rect 16587 696 16599 898
rect 16659 792 16671 898
rect 16707 792 16719 898
rect 16899 888 16911 898
rect 16971 312 16983 898
rect 17043 24 17055 898
rect 17139 192 17151 898
rect 17643 888 17655 898
rect 17835 336 17847 898
rect 18147 888 18159 898
rect 18219 408 18231 898
rect 18339 408 18351 898
rect 18867 600 18879 898
rect 19059 312 19071 898
rect 19083 240 19095 898
rect 19155 432 19167 898
rect 19227 600 19239 898
rect 19395 864 19407 898
rect 19419 432 19431 898
rect 19467 216 19479 898
rect 19515 72 19527 898
rect 19539 864 19551 898
rect 19563 168 19575 898
rect 19635 120 19647 898
rect 20595 432 20607 898
rect 20667 432 20679 898
rect 20680 418 20698 432
rect 17056 10 17074 24
rect 17055 0 17067 10
rect 20679 0 20691 418
rect 20859 360 20871 898
rect 20955 408 20967 898
rect 21027 696 21039 898
rect 21123 720 21135 898
rect 21291 840 21303 898
rect 21315 384 21327 898
rect 22059 696 22071 898
rect 22131 720 22143 898
rect 22203 312 22215 898
rect 22467 648 22479 898
rect 22515 768 22527 898
rect 22635 648 22647 898
rect 22659 456 22671 898
rect 22779 288 22791 898
rect 22803 144 22815 898
rect 22851 552 22863 898
rect 22899 648 22911 898
rect 23259 480 23271 898
rect 23427 504 23439 898
rect 23475 576 23487 898
rect 23499 888 23511 898
rect 24027 96 24039 898
rect 24123 696 24135 898
rect 24291 744 24303 898
rect 24315 144 24327 898
rect 24339 792 24351 898
rect 24435 864 24447 898
rect 24531 672 24543 898
rect 24651 600 24663 898
rect 25251 624 25263 898
rect 25347 720 25359 898
rect 25515 816 25527 898
rect 26067 24 26079 898
rect 26091 96 26103 514
rect 26091 48 26103 58
rect 26115 48 26127 250
rect 26211 0 26411 898
rect 26465 83 26535 95
rect 26465 59 26535 71
rect 26465 35 26535 47
rect 26465 11 26535 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 6867
box 0 0 1464 799
use inv g8075
timestamp 1386238110
transform 1 0 1587 0 1 6867
box 0 0 120 799
use rowcrosser StatusRegEn
timestamp 1386086759
transform 1 0 1707 0 1 6867
box 0 0 48 799
use nand2 g7994
timestamp 1386234792
transform 1 0 1755 0 1 6867
box 0 0 96 799
use nand2 g8032
timestamp 1386234792
transform 1 0 1851 0 1 6867
box 0 0 96 799
use nor2 g7941
timestamp 1386235306
transform 1 0 1947 0 1 6867
box 0 0 120 799
use nand2 g8197
timestamp 1386234792
transform 1 0 2067 0 1 6867
box 0 0 96 799
use nand2 g8043
timestamp 1386234792
transform 1 0 2163 0 1 6867
box 0 0 96 799
use nand3 g8112
timestamp 1386234893
transform 1 0 2259 0 1 6867
box 0 0 120 799
use inv g7923
timestamp 1386238110
transform 1 0 2379 0 1 6867
box 0 0 120 799
use nand2 g8060
timestamp 1386234792
transform 1 0 2499 0 1 6867
box 0 0 96 799
use nand2 g7895
timestamp 1386234792
transform 1 0 2595 0 1 6867
box 0 0 96 799
use nand3 g7942
timestamp 1386234893
transform 1 0 2691 0 1 6867
box 0 0 120 799
use nand2 g8182
timestamp 1386234792
transform 1 0 2811 0 1 6867
box 0 0 96 799
use and2 g8066
timestamp 1386234845
transform 1 0 2907 0 1 6867
box 0 0 120 799
use nand3 g8169
timestamp 1386234893
transform 1 0 3027 0 1 6867
box 0 0 120 799
use inv g7934
timestamp 1386238110
transform 1 0 3147 0 1 6867
box 0 0 120 799
use nand2 g8107
timestamp 1386234792
transform 1 0 3267 0 1 6867
box 0 0 96 799
use nand3 g8229
timestamp 1386234893
transform 1 0 3363 0 1 6867
box 0 0 120 799
use inv g7912
timestamp 1386238110
transform 1 0 3483 0 1 6867
box 0 0 120 799
use nand4 g8039
timestamp 1386234936
transform 1 0 3603 0 1 6867
box 0 0 144 799
use nand2 g8046
timestamp 1386234792
transform 1 0 3747 0 1 6867
box 0 0 96 799
use nand2 g8123
timestamp 1386234792
transform 1 0 3843 0 1 6867
box 0 0 96 799
use nand2 g8222
timestamp 1386234792
transform 1 0 3939 0 1 6867
box 0 0 96 799
use nand2 g8102
timestamp 1386234792
transform 1 0 4035 0 1 6867
box 0 0 96 799
use nand2 g8098
timestamp 1386234792
transform 1 0 4131 0 1 6867
box 0 0 96 799
use nand2 g8012
timestamp 1386234792
transform 1 0 4227 0 1 6867
box 0 0 96 799
use and2 g8187
timestamp 1386234845
transform 1 0 4323 0 1 6867
box 0 0 120 799
use nand2 g7951
timestamp 1386234792
transform 1 0 4443 0 1 6867
box 0 0 96 799
use nand3 g8135
timestamp 1386234893
transform 1 0 4539 0 1 6867
box 0 0 120 799
use inv g8171
timestamp 1386238110
transform 1 0 4659 0 1 6867
box 0 0 120 799
use nand3 g8154
timestamp 1386234893
transform 1 0 4779 0 1 6867
box 0 0 120 799
use nor2 g8130
timestamp 1386235306
transform 1 0 4899 0 1 6867
box 0 0 120 799
use and2 g8027
timestamp 1386234845
transform 1 0 5019 0 1 6867
box 0 0 120 799
use nand3 g8082
timestamp 1386234893
transform 1 0 5139 0 1 6867
box 0 0 120 799
use nor2 g8035
timestamp 1386235306
transform 1 0 5259 0 1 6867
box 0 0 120 799
use rowcrosser MemEn
timestamp 1386086759
transform 1 0 5379 0 1 6867
box 0 0 48 799
use nand3 g8019
timestamp 1386234893
transform 1 0 5427 0 1 6867
box 0 0 120 799
use nand2 g8168
timestamp 1386234792
transform 1 0 5547 0 1 6867
box 0 0 96 799
use nand2 g8238
timestamp 1386234792
transform 1 0 5643 0 1 6867
box 0 0 96 799
use nand2 g7989
timestamp 1386234792
transform 1 0 5739 0 1 6867
box 0 0 96 799
use nand3 g8225
timestamp 1386234893
transform 1 0 5835 0 1 6867
box 0 0 120 799
use nand2 g8143
timestamp 1386234792
transform 1 0 5955 0 1 6867
box 0 0 96 799
use mux2 g2
timestamp 1386235218
transform 1 0 6051 0 1 6867
box 0 0 192 799
use nand3 g8042
timestamp 1386234893
transform 1 0 6243 0 1 6867
box 0 0 120 799
use nand2 g8069
timestamp 1386234792
transform 1 0 6363 0 1 6867
box 0 0 96 799
use nand3 g8149
timestamp 1386234893
transform 1 0 6459 0 1 6867
box 0 0 120 799
use nand2 g7926
timestamp 1386234792
transform 1 0 6579 0 1 6867
box 0 0 96 799
use nand2 g7985
timestamp 1386234792
transform 1 0 6675 0 1 6867
box 0 0 96 799
use nand3 g8249
timestamp 1386234893
transform 1 0 6771 0 1 6867
box 0 0 120 799
use inv g8064
timestamp 1386238110
transform 1 0 6891 0 1 6867
box 0 0 120 799
use nand2 g8235
timestamp 1386234792
transform 1 0 7011 0 1 6867
box 0 0 96 799
use nand2 g7948
timestamp 1386234792
transform 1 0 7107 0 1 6867
box 0 0 96 799
use nand2 g8058
timestamp 1386234792
transform 1 0 7203 0 1 6867
box 0 0 96 799
use nand2 g8009
timestamp 1386234792
transform 1 0 7299 0 1 6867
box 0 0 96 799
use and2 g7903
timestamp 1386234845
transform 1 0 7395 0 1 6867
box 0 0 120 799
use nand2 g7939
timestamp 1386234792
transform 1 0 7515 0 1 6867
box 0 0 96 799
use nor2 g8055
timestamp 1386235306
transform 1 0 7611 0 1 6867
box 0 0 120 799
use nand2 g8088
timestamp 1386234792
transform 1 0 7731 0 1 6867
box 0 0 96 799
use nand2 g7947
timestamp 1386234792
transform 1 0 7827 0 1 6867
box 0 0 96 799
use inv g8214
timestamp 1386238110
transform 1 0 7923 0 1 6867
box 0 0 120 799
use nor2 g8056
timestamp 1386235306
transform 1 0 8043 0 1 6867
box 0 0 120 799
use nand2 g8183
timestamp 1386234792
transform 1 0 8163 0 1 6867
box 0 0 96 799
use nand2 g8170
timestamp 1386234792
transform 1 0 8259 0 1 6867
box 0 0 96 799
use nand2 g8124
timestamp 1386234792
transform 1 0 8355 0 1 6867
box 0 0 96 799
use nand2 g8106
timestamp 1386234792
transform 1 0 8451 0 1 6867
box 0 0 96 799
use nand2 g8119
timestamp 1386234792
transform 1 0 8547 0 1 6867
box 0 0 96 799
use nor2 g8146
timestamp 1386235306
transform 1 0 8643 0 1 6867
box 0 0 120 799
use nand2 g8127
timestamp 1386234792
transform 1 0 8763 0 1 6867
box 0 0 96 799
use nand2 g8155
timestamp 1386234792
transform 1 0 8859 0 1 6867
box 0 0 96 799
use nand2 g7909
timestamp 1386234792
transform 1 0 8955 0 1 6867
box 0 0 96 799
use nand3 g7890
timestamp 1386234893
transform 1 0 9051 0 1 6867
box 0 0 120 799
use nand3 g8033
timestamp 1386234893
transform 1 0 9171 0 1 6867
box 0 0 120 799
use nand3 g7921
timestamp 1386234893
transform 1 0 9291 0 1 6867
box 0 0 120 799
use nand2 g8252
timestamp 1386234792
transform 1 0 9411 0 1 6867
box 0 0 96 799
use rowcrosser Flags_91_1_93_
timestamp 1386086759
transform 1 0 9507 0 1 6867
box 0 0 48 799
use inv g7978
timestamp 1386238110
transform 1 0 9555 0 1 6867
box 0 0 120 799
use inv g7930
timestamp 1386238110
transform 1 0 9675 0 1 6867
box 0 0 120 799
use nand4 g7972
timestamp 1386234936
transform 1 0 9795 0 1 6867
box 0 0 144 799
use nand2 g8240
timestamp 1386234792
transform 1 0 9939 0 1 6867
box 0 0 96 799
use nand2 g8054
timestamp 1386234792
transform 1 0 10035 0 1 6867
box 0 0 96 799
use inv g8139
timestamp 1386238110
transform 1 0 10131 0 1 6867
box 0 0 120 799
use nand2 g8023
timestamp 1386234792
transform 1 0 10251 0 1 6867
box 0 0 96 799
use rowcrosser ALE
timestamp 1386086759
transform 1 0 10347 0 1 6867
box 0 0 48 799
use nand2 g8118
timestamp 1386234792
transform 1 0 10395 0 1 6867
box 0 0 96 799
use nand2 g7981
timestamp 1386234792
transform 1 0 10491 0 1 6867
box 0 0 96 799
use nand2 g8111
timestamp 1386234792
transform 1 0 10587 0 1 6867
box 0 0 96 799
use nor2 g8120
timestamp 1386235306
transform 1 0 10683 0 1 6867
box 0 0 120 799
use and2 g8091
timestamp 1386234845
transform 1 0 10803 0 1 6867
box 0 0 120 799
use and2 g7918
timestamp 1386234845
transform 1 0 10923 0 1 6867
box 0 0 120 799
use nand4 g8134
timestamp 1386234936
transform 1 0 11043 0 1 6867
box 0 0 144 799
use nand2 g8050
timestamp 1386234792
transform 1 0 11187 0 1 6867
box 0 0 96 799
use nand3 g8218
timestamp 1386234893
transform 1 0 11283 0 1 6867
box 0 0 120 799
use inv g7945
timestamp 1386238110
transform 1 0 11403 0 1 6867
box 0 0 120 799
use and2 g7995
timestamp 1386234845
transform 1 0 11523 0 1 6867
box 0 0 120 799
use nand3 g7964
timestamp 1386234893
transform 1 0 11643 0 1 6867
box 0 0 120 799
use nand2 g8198
timestamp 1386234792
transform 1 0 11763 0 1 6867
box 0 0 96 799
use inv g7901
timestamp 1386238110
transform 1 0 11859 0 1 6867
box 0 0 120 799
use nand2 g8199
timestamp 1386234792
transform 1 0 11979 0 1 6867
box 0 0 96 799
use nand2 g8221
timestamp 1386234792
transform 1 0 12075 0 1 6867
box 0 0 96 799
use inv g8220
timestamp 1386238110
transform 1 0 12171 0 1 6867
box 0 0 120 799
use nand2 g8230
timestamp 1386234792
transform 1 0 12291 0 1 6867
box 0 0 96 799
use nand2 g8004
timestamp 1386234792
transform 1 0 12387 0 1 6867
box 0 0 96 799
use nand2 rm_assigns_buf_StatusReg_1
timestamp 1386234792
transform 1 0 12483 0 1 6867
box 0 0 96 799
use buffer g8074
timestamp 1386236986
transform 1 0 12579 0 1 6867
box 0 0 120 799
use nand4 g8209
timestamp 1386234936
transform 1 0 12699 0 1 6867
box 0 0 144 799
use inv g8103
timestamp 1386238110
transform 1 0 12843 0 1 6867
box 0 0 120 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 12963 0 1 6867
box 0 0 48 799
use inv g8180
timestamp 1386238110
transform 1 0 13011 0 1 6867
box 0 0 120 799
use nand2 g8005
timestamp 1386234792
transform 1 0 13131 0 1 6867
box 0 0 96 799
use nand3 g8052
timestamp 1386234893
transform 1 0 13227 0 1 6867
box 0 0 120 799
use nand2 g8136
timestamp 1386234792
transform 1 0 13347 0 1 6867
box 0 0 96 799
use nand2 g8110
timestamp 1386234792
transform 1 0 13443 0 1 6867
box 0 0 96 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 13539 0 1 6867
box 0 0 96 799
use scandtype g7922
timestamp 1386241841
transform 1 0 13635 0 1 6867
box 0 0 624 799
use nand2 stateSub_reg_91_2_93_
timestamp 1386234792
transform 1 0 14259 0 1 6867
box 0 0 96 799
use scandtype g7943
timestamp 1386241841
transform 1 0 14355 0 1 6867
box 0 0 624 799
use nand2 g8024
timestamp 1386234792
transform 1 0 14979 0 1 6867
box 0 0 96 799
use nand2 g8099
timestamp 1386234792
transform 1 0 15075 0 1 6867
box 0 0 96 799
use nand3 g7898
timestamp 1386234893
transform 1 0 15171 0 1 6867
box 0 0 120 799
use nand4 g8057
timestamp 1386234936
transform 1 0 15291 0 1 6867
box 0 0 144 799
use nand2 g8190
timestamp 1386234792
transform 1 0 15435 0 1 6867
box 0 0 96 799
use nand2 g8045
timestamp 1386234792
transform 1 0 15531 0 1 6867
box 0 0 96 799
use inv g7913
timestamp 1386238110
transform 1 0 15627 0 1 6867
box 0 0 120 799
use nand4 g8092
timestamp 1386234936
transform 1 0 15747 0 1 6867
box 0 0 144 799
use inv g8018
timestamp 1386238110
transform 1 0 15891 0 1 6867
box 0 0 120 799
use and2 g8081
timestamp 1386234845
transform 1 0 16011 0 1 6867
box 0 0 120 799
use nand2 g8234
timestamp 1386234792
transform 1 0 16131 0 1 6867
box 0 0 96 799
use nor2 StatusReg_reg_91_1_93_
timestamp 1386235306
transform 1 0 16227 0 1 6867
box 0 0 120 799
use scandtype g7933
timestamp 1386241841
transform 1 0 16347 0 1 6867
box 0 0 624 799
use nand2 g8028
timestamp 1386234792
transform 1 0 16971 0 1 6867
box 0 0 96 799
use nand3 g8213
timestamp 1386234893
transform 1 0 17067 0 1 6867
box 0 0 120 799
use and2 g7963
timestamp 1386234845
transform 1 0 17187 0 1 6867
box 0 0 120 799
use nand2 g8096
timestamp 1386234792
transform 1 0 17307 0 1 6867
box 0 0 96 799
use nand2 g8212
timestamp 1386234792
transform 1 0 17403 0 1 6867
box 0 0 96 799
use nand2 g7911
timestamp 1386234792
transform 1 0 17499 0 1 6867
box 0 0 96 799
use nand4 g8015
timestamp 1386234936
transform 1 0 17595 0 1 6867
box 0 0 144 799
use nand3 g8084
timestamp 1386234893
transform 1 0 17739 0 1 6867
box 0 0 120 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 17859 0 1 6867
box 0 0 48 799
use nor2 g8200
timestamp 1386235306
transform 1 0 17907 0 1 6867
box 0 0 120 799
use nand2 g7896
timestamp 1386234792
transform 1 0 18027 0 1 6867
box 0 0 96 799
use nor2 g8108
timestamp 1386235306
transform 1 0 18123 0 1 6867
box 0 0 120 799
use nand3 g8049
timestamp 1386234893
transform 1 0 18243 0 1 6867
box 0 0 120 799
use nand2 g8144
timestamp 1386234792
transform 1 0 18363 0 1 6867
box 0 0 96 799
use inv g8159
timestamp 1386238110
transform 1 0 18459 0 1 6867
box 0 0 120 799
use and2 g8177
timestamp 1386234845
transform 1 0 18579 0 1 6867
box 0 0 120 799
use nand2 g7996
timestamp 1386234792
transform 1 0 18699 0 1 6867
box 0 0 96 799
use nand2 g8036
timestamp 1386234792
transform 1 0 18795 0 1 6867
box 0 0 96 799
use nand2 g8226
timestamp 1386234792
transform 1 0 18891 0 1 6867
box 0 0 96 799
use nand2 g7929
timestamp 1386234792
transform 1 0 18987 0 1 6867
box 0 0 96 799
use nand2 g7979
timestamp 1386234792
transform 1 0 19083 0 1 6867
box 0 0 96 799
use nand2 g7893
timestamp 1386234792
transform 1 0 19179 0 1 6867
box 0 0 96 799
use nand3 g7924
timestamp 1386234893
transform 1 0 19275 0 1 6867
box 0 0 120 799
use nand3 g8089
timestamp 1386234893
transform 1 0 19395 0 1 6867
box 0 0 120 799
use nand2 g8206
timestamp 1386234792
transform 1 0 19515 0 1 6867
box 0 0 96 799
use nand2 g8237
timestamp 1386234792
transform 1 0 19611 0 1 6867
box 0 0 96 799
use inv g8016
timestamp 1386238110
transform 1 0 19707 0 1 6867
box 0 0 120 799
use and2 g8181
timestamp 1386234845
transform 1 0 19827 0 1 6867
box 0 0 120 799
use nor2 g8216
timestamp 1386235306
transform 1 0 19947 0 1 6867
box 0 0 120 799
use nor2 StatusReg_reg_91_0_93_
timestamp 1386235306
transform 1 0 20067 0 1 6867
box 0 0 120 799
use scandtype g8253
timestamp 1386241841
transform 1 0 20187 0 1 6867
box 0 0 624 799
use inv g8186
timestamp 1386238110
transform 1 0 20811 0 1 6867
box 0 0 120 799
use inv g7946
timestamp 1386238110
transform 1 0 20931 0 1 6867
box 0 0 120 799
use nand2 g8090
timestamp 1386234792
transform 1 0 21051 0 1 6867
box 0 0 96 799
use and2 g8195
timestamp 1386234845
transform 1 0 21147 0 1 6867
box 0 0 120 799
use inv g8223
timestamp 1386238110
transform 1 0 21267 0 1 6867
box 0 0 120 799
use nand2 g8077
timestamp 1386234792
transform 1 0 21387 0 1 6867
box 0 0 96 799
use inv g8133
timestamp 1386238110
transform 1 0 21483 0 1 6867
box 0 0 120 799
use nand2 g7971
timestamp 1386234792
transform 1 0 21603 0 1 6867
box 0 0 96 799
use nand2 g8041
timestamp 1386234792
transform 1 0 21699 0 1 6867
box 0 0 96 799
use and2 g8002
timestamp 1386234845
transform 1 0 21795 0 1 6867
box 0 0 120 799
use nand2 g8128
timestamp 1386234792
transform 1 0 21915 0 1 6867
box 0 0 96 799
use and2 g8029
timestamp 1386234845
transform 1 0 22011 0 1 6867
box 0 0 120 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 22131 0 1 6867
box 0 0 48 799
use nand3 g8100
timestamp 1386234893
transform 1 0 22179 0 1 6867
box 0 0 120 799
use nand2 g8117
timestamp 1386234792
transform 1 0 22299 0 1 6867
box 0 0 96 799
use nand2 g8167
timestamp 1386234792
transform 1 0 22395 0 1 6867
box 0 0 96 799
use nand2 g7982
timestamp 1386234792
transform 1 0 22491 0 1 6867
box 0 0 96 799
use nand2 g8227
timestamp 1386234792
transform 1 0 22587 0 1 6867
box 0 0 96 799
use inv g8191
timestamp 1386238110
transform 1 0 22683 0 1 6867
box 0 0 120 799
use nand3 g7975
timestamp 1386234893
transform 1 0 22803 0 1 6867
box 0 0 120 799
use nand2 g8073
timestamp 1386234792
transform 1 0 22923 0 1 6867
box 0 0 96 799
use nand3 g7967
timestamp 1386234893
transform 1 0 23019 0 1 6867
box 0 0 120 799
use nor2 g7925
timestamp 1386235306
transform 1 0 23139 0 1 6867
box 0 0 120 799
use nand3 g8163
timestamp 1386234893
transform 1 0 23259 0 1 6867
box 0 0 120 799
use and2 g7969
timestamp 1386234845
transform 1 0 23379 0 1 6867
box 0 0 120 799
use inv g8051
timestamp 1386238110
transform 1 0 23499 0 1 6867
box 0 0 120 799
use nand2 g8147
timestamp 1386234792
transform 1 0 23619 0 1 6867
box 0 0 96 799
use nand2 g7955
timestamp 1386234792
transform 1 0 23715 0 1 6867
box 0 0 96 799
use nand4 g7928
timestamp 1386234936
transform 1 0 23811 0 1 6867
box 0 0 144 799
use nand2 g8030
timestamp 1386234792
transform 1 0 23955 0 1 6867
box 0 0 96 799
use nor2 g8217
timestamp 1386235306
transform 1 0 24051 0 1 6867
box 0 0 120 799
use and2 g7899
timestamp 1386234845
transform 1 0 24171 0 1 6867
box 0 0 120 799
use nand4 g7900
timestamp 1386234936
transform 1 0 24291 0 1 6867
box 0 0 144 799
use nand2 g8114
timestamp 1386234792
transform 1 0 24435 0 1 6867
box 0 0 96 799
use nand3 g8174
timestamp 1386234893
transform 1 0 24531 0 1 6867
box 0 0 120 799
use nand2 g8241
timestamp 1386234792
transform 1 0 24651 0 1 6867
box 0 0 96 799
use nand2 g7894
timestamp 1386234792
transform 1 0 24747 0 1 6867
box 0 0 96 799
use nand3 g7888
timestamp 1386234893
transform 1 0 24843 0 1 6867
box 0 0 120 799
use nand4 g8067
timestamp 1386234936
transform 1 0 24963 0 1 6867
box 0 0 144 799
use nand2 g7990
timestamp 1386234792
transform 1 0 25107 0 1 6867
box 0 0 96 799
use inv g8158
timestamp 1386238110
transform 1 0 25203 0 1 6867
box 0 0 120 799
use and2 g8063
timestamp 1386234845
transform 1 0 25323 0 1 6867
box 0 0 120 799
use nand2 g8257
timestamp 1386234792
transform 1 0 25443 0 1 6867
box 0 0 96 799
use inv OpcodeCondIn_91_4_93_
timestamp 1386238110
transform 1 0 25539 0 1 6867
box 0 0 120 799
use rowcrosser StatusReg_91_2_93_
timestamp 1386086759
transform 1 0 25659 0 1 6867
box 0 0 48 799
use rowcrosser PcEn
timestamp 1386086759
transform 1 0 25707 0 1 6867
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 26091 0 1 6867
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 898
box 0 0 1464 799
use and2 stateSub_reg_91_0_93_
timestamp 1386234845
transform 1 0 1587 0 1 898
box 0 0 120 799
use rowcrosser SysBus_91_2_93_
timestamp 1386086759
transform 1 0 1707 0 1 898
box 0 0 48 799
use scandtype g7886
timestamp 1386241841
transform 1 0 1755 0 1 898
box 0 0 624 799
use nand3 g7892
timestamp 1386234893
transform 1 0 2379 0 1 898
box 0 0 120 799
use nand3 g8020
timestamp 1386234893
transform 1 0 2499 0 1 898
box 0 0 120 799
use nand2 g8150
timestamp 1386234792
transform 1 0 2619 0 1 898
box 0 0 96 799
use and2 g8178
timestamp 1386234845
transform 1 0 2715 0 1 898
box 0 0 120 799
use and2 state_reg_91_1_93_
timestamp 1386234845
transform 1 0 2835 0 1 898
box 0 0 120 799
use scandtype g8250
timestamp 1386241841
transform 1 0 2955 0 1 898
box 0 0 624 799
use inv g8148
timestamp 1386238110
transform 1 0 3579 0 1 898
box 0 0 120 799
use nand2 g7976
timestamp 1386234792
transform 1 0 3699 0 1 898
box 0 0 96 799
use nand3 g7993
timestamp 1386234893
transform 1 0 3795 0 1 898
box 0 0 120 799
use nor2 g8196
timestamp 1386235306
transform 1 0 3915 0 1 898
box 0 0 120 799
use nand2 g8211
timestamp 1386234792
transform 1 0 4035 0 1 898
box 0 0 96 799
use inv g8175
timestamp 1386238110
transform 1 0 4131 0 1 898
box 0 0 120 799
use nand2 g8078
timestamp 1386234792
transform 1 0 4251 0 1 898
box 0 0 96 799
use nor2 g8093
timestamp 1386235306
transform 1 0 4347 0 1 898
box 0 0 120 799
use nand2 g7974
timestamp 1386234792
transform 1 0 4467 0 1 898
box 0 0 96 799
use nand2 g8104
timestamp 1386234792
transform 1 0 4563 0 1 898
box 0 0 96 799
use nor2 g7940
timestamp 1386235306
transform 1 0 4659 0 1 898
box 0 0 120 799
use and2 g8160
timestamp 1386234845
transform 1 0 4779 0 1 898
box 0 0 120 799
use xor2 g8076
timestamp 1386237344
transform 1 0 4899 0 1 898
box 0 0 192 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 5091 0 1 898
box 0 0 96 799
use scandtype g8161
timestamp 1386241841
transform 1 0 5187 0 1 898
box 0 0 624 799
use nand2 g8224
timestamp 1386234792
transform 1 0 5811 0 1 898
box 0 0 96 799
use nand2 g8094
timestamp 1386234792
transform 1 0 5907 0 1 898
box 0 0 96 799
use and2 g7910
timestamp 1386234845
transform 1 0 6003 0 1 898
box 0 0 120 799
use nand4 g8121
timestamp 1386234936
transform 1 0 6123 0 1 898
box 0 0 144 799
use and2 g8037
timestamp 1386234845
transform 1 0 6267 0 1 898
box 0 0 120 799
use nand2 g8189
timestamp 1386234792
transform 1 0 6387 0 1 898
box 0 0 96 799
use nand2 g8125
timestamp 1386234792
transform 1 0 6483 0 1 898
box 0 0 96 799
use nand2 g7915
timestamp 1386234792
transform 1 0 6579 0 1 898
box 0 0 96 799
use nand4 g8232
timestamp 1386234936
transform 1 0 6675 0 1 898
box 0 0 144 799
use inv g8152
timestamp 1386238110
transform 1 0 6819 0 1 898
box 0 0 120 799
use nand3 g8080
timestamp 1386234893
transform 1 0 6939 0 1 898
box 0 0 120 799
use nand2 g7937
timestamp 1386234792
transform 1 0 7059 0 1 898
box 0 0 96 799
use nand2 g7997
timestamp 1386234792
transform 1 0 7155 0 1 898
box 0 0 96 799
use nand2 g8236
timestamp 1386234792
transform 1 0 7251 0 1 898
box 0 0 96 799
use nor2 g8101
timestamp 1386235306
transform 1 0 7347 0 1 898
box 0 0 120 799
use nand3 g8011
timestamp 1386234893
transform 1 0 7467 0 1 898
box 0 0 120 799
use nand2 g7919
timestamp 1386234792
transform 1 0 7587 0 1 898
box 0 0 96 799
use nor2 g8185
timestamp 1386235306
transform 1 0 7683 0 1 898
box 0 0 120 799
use nand2 g7927
timestamp 1386234792
transform 1 0 7803 0 1 898
box 0 0 96 799
use nand2 g8255
timestamp 1386234792
transform 1 0 7899 0 1 898
box 0 0 96 799
use inv g8086
timestamp 1386238110
transform 1 0 7995 0 1 898
box 0 0 120 799
use and2 g7962
timestamp 1386234845
transform 1 0 8115 0 1 898
box 0 0 120 799
use nand2 g8192
timestamp 1386234792
transform 1 0 8235 0 1 898
box 0 0 96 799
use nand2 g7988
timestamp 1386234792
transform 1 0 8331 0 1 898
box 0 0 96 799
use nand3 g8254
timestamp 1386234893
transform 1 0 8427 0 1 898
box 0 0 120 799
use inv g8116
timestamp 1386238110
transform 1 0 8547 0 1 898
box 0 0 120 799
use nor2 g8145
timestamp 1386235306
transform 1 0 8667 0 1 898
box 0 0 120 799
use nand2 g8166
timestamp 1386234792
transform 1 0 8787 0 1 898
box 0 0 96 799
use nand2 g7907
timestamp 1386234792
transform 1 0 8883 0 1 898
box 0 0 96 799
use nor2 g8014
timestamp 1386235306
transform 1 0 8979 0 1 898
box 0 0 120 799
use nand3 g7959
timestamp 1386234893
transform 1 0 9099 0 1 898
box 0 0 120 799
use nand4 g8001
timestamp 1386234936
transform 1 0 9219 0 1 898
box 0 0 144 799
use nand3 g7998
timestamp 1386234893
transform 1 0 9363 0 1 898
box 0 0 120 799
use nand3 g8228
timestamp 1386234893
transform 1 0 9483 0 1 898
box 0 0 120 799
use nand2 g7987
timestamp 1386234792
transform 1 0 9603 0 1 898
box 0 0 96 799
use nand3 g8072
timestamp 1386234893
transform 1 0 9699 0 1 898
box 0 0 120 799
use nand4 g7966
timestamp 1386234936
transform 1 0 9819 0 1 898
box 0 0 144 799
use inv g8105
timestamp 1386238110
transform 1 0 9963 0 1 898
box 0 0 120 799
use nand4 g7897
timestamp 1386234936
transform 1 0 10083 0 1 898
box 0 0 144 799
use nand4 g8129
timestamp 1386234936
transform 1 0 10227 0 1 898
box 0 0 144 799
use nand2 g8122
timestamp 1386234792
transform 1 0 10371 0 1 898
box 0 0 96 799
use and2 g8059
timestamp 1386234845
transform 1 0 10467 0 1 898
box 0 0 120 799
use nand2 g8097
timestamp 1386234792
transform 1 0 10587 0 1 898
box 0 0 96 799
use and2 g8062
timestamp 1386234845
transform 1 0 10683 0 1 898
box 0 0 120 799
use rowcrosser ENB
timestamp 1386086759
transform 1 0 10803 0 1 898
box 0 0 48 799
use nand3 g8025
timestamp 1386234893
transform 1 0 10851 0 1 898
box 0 0 120 799
use nand4 g8247
timestamp 1386234936
transform 1 0 10971 0 1 898
box 0 0 144 799
use inv IntStatus_reg
timestamp 1386238110
transform 1 0 11115 0 1 898
box 0 0 120 799
use scanreg g8131
timestamp 1386241447
transform 1 0 11235 0 1 898
box 0 0 720 799
use nand2 g8087
timestamp 1386234792
transform 1 0 11955 0 1 898
box 0 0 96 799
use inv g7970
timestamp 1386238110
transform 1 0 12051 0 1 898
box 0 0 120 799
use nand3 g7932
timestamp 1386234893
transform 1 0 12171 0 1 898
box 0 0 120 799
use nand4 g7991
timestamp 1386234936
transform 1 0 12291 0 1 898
box 0 0 144 799
use nand4 g8137
timestamp 1386234936
transform 1 0 12435 0 1 898
box 0 0 144 799
use nand3 g8201
timestamp 1386234893
transform 1 0 12579 0 1 898
box 0 0 120 799
use nand3 g7952
timestamp 1386234893
transform 1 0 12699 0 1 898
box 0 0 120 799
use nand3 g7936
timestamp 1386234893
transform 1 0 12819 0 1 898
box 0 0 120 799
use nand2 g8242
timestamp 1386234792
transform 1 0 12939 0 1 898
box 0 0 96 799
use nand2 g8207
timestamp 1386234792
transform 1 0 13035 0 1 898
box 0 0 96 799
use nand2 g7889
timestamp 1386234792
transform 1 0 13131 0 1 898
box 0 0 96 799
use nand4 g8044
timestamp 1386234936
transform 1 0 13227 0 1 898
box 0 0 144 799
use nand2 g8006
timestamp 1386234792
transform 1 0 13371 0 1 898
box 0 0 96 799
use and2 g8173
timestamp 1386234845
transform 1 0 13467 0 1 898
box 0 0 120 799
use nand2 g7983
timestamp 1386234792
transform 1 0 13587 0 1 898
box 0 0 96 799
use and2 g7956
timestamp 1386234845
transform 1 0 13683 0 1 898
box 0 0 120 799
use inv g8157
timestamp 1386238110
transform 1 0 13803 0 1 898
box 0 0 120 799
use nor2 g8068
timestamp 1386235306
transform 1 0 13923 0 1 898
box 0 0 120 799
use nand3 g8040
timestamp 1386234893
transform 1 0 14043 0 1 898
box 0 0 120 799
use nand2 g7880
timestamp 1386234792
transform 1 0 14163 0 1 898
box 0 0 96 799
use nand4 g8140
timestamp 1386234936
transform 1 0 14259 0 1 898
box 0 0 144 799
use nand3 g8141
timestamp 1386234893
transform 1 0 14403 0 1 898
box 0 0 120 799
use and2 g8210
timestamp 1386234845
transform 1 0 14523 0 1 898
box 0 0 120 799
use nor2 g8003
timestamp 1386235306
transform 1 0 14643 0 1 898
box 0 0 120 799
use nand2 g8203
timestamp 1386234792
transform 1 0 14763 0 1 898
box 0 0 96 799
use xor2 g8065
timestamp 1386237344
transform 1 0 14859 0 1 898
box 0 0 192 799
use nand2 g8113
timestamp 1386234792
transform 1 0 15051 0 1 898
box 0 0 96 799
use nor2 g7977
timestamp 1386235306
transform 1 0 15147 0 1 898
box 0 0 120 799
use nand2 g8070
timestamp 1386234792
transform 1 0 15267 0 1 898
box 0 0 96 799
use nand3 g8038
timestamp 1386234893
transform 1 0 15363 0 1 898
box 0 0 120 799
use inv IRQ2_reg
timestamp 1386238110
transform 1 0 15483 0 1 898
box 0 0 120 799
use scandtype g8233
timestamp 1386241841
transform 1 0 15603 0 1 898
box 0 0 624 799
use nand2 g7980
timestamp 1386234792
transform 1 0 16227 0 1 898
box 0 0 96 799
use nand2 g7954
timestamp 1386234792
transform 1 0 16323 0 1 898
box 0 0 96 799
use nand4 g7920
timestamp 1386234936
transform 1 0 16419 0 1 898
box 0 0 144 799
use nor2 g8151
timestamp 1386235306
transform 1 0 16563 0 1 898
box 0 0 120 799
use and2 g7968
timestamp 1386234845
transform 1 0 16683 0 1 898
box 0 0 120 799
use and2 g8138
timestamp 1386234845
transform 1 0 16803 0 1 898
box 0 0 120 799
use nand2 g8188
timestamp 1386234792
transform 1 0 16923 0 1 898
box 0 0 96 799
use rowcrosser g7914
timestamp 1386086759
transform 1 0 17019 0 1 898
box 0 0 48 799
use nand2 g8176
timestamp 1386234792
transform 1 0 17067 0 1 898
box 0 0 96 799
use and2 g8172
timestamp 1386234845
transform 1 0 17163 0 1 898
box 0 0 120 799
use nand2 g8026
timestamp 1386234792
transform 1 0 17283 0 1 898
box 0 0 96 799
use nand3 g8031
timestamp 1386234893
transform 1 0 17379 0 1 898
box 0 0 120 799
use nor2 g7935
timestamp 1386235306
transform 1 0 17499 0 1 898
box 0 0 120 799
use nor2 g8162
timestamp 1386235306
transform 1 0 17619 0 1 898
box 0 0 120 799
use nor2 g8095
timestamp 1386235306
transform 1 0 17739 0 1 898
box 0 0 120 799
use nand2 g7950
timestamp 1386234792
transform 1 0 17859 0 1 898
box 0 0 96 799
use inv g8008
timestamp 1386238110
transform 1 0 17955 0 1 898
box 0 0 120 799
use nand2 g8013
timestamp 1386234792
transform 1 0 18075 0 1 898
box 0 0 96 799
use nand2 g7984
timestamp 1386234792
transform 1 0 18171 0 1 898
box 0 0 96 799
use nand2 IRQ1_reg
timestamp 1386234792
transform 1 0 18267 0 1 898
box 0 0 96 799
use scandtype g7986
timestamp 1386241841
transform 1 0 18363 0 1 898
box 0 0 624 799
use nand3 g7904
timestamp 1386234893
transform 1 0 18987 0 1 898
box 0 0 120 799
use nand4 g8164
timestamp 1386234936
transform 1 0 19107 0 1 898
box 0 0 144 799
use nor2 g7949
timestamp 1386235306
transform 1 0 19251 0 1 898
box 0 0 120 799
use and2 g8017
timestamp 1386234845
transform 1 0 19371 0 1 898
box 0 0 120 799
use nand2 g8010
timestamp 1386234792
transform 1 0 19491 0 1 898
box 0 0 96 799
use nand2 g8165
timestamp 1386234792
transform 1 0 19587 0 1 898
box 0 0 96 799
use inv g8245
timestamp 1386238110
transform 1 0 19683 0 1 898
box 0 0 120 799
use inv g8034
timestamp 1386238110
transform 1 0 19803 0 1 898
box 0 0 120 799
use nand2 g8215
timestamp 1386234792
transform 1 0 19923 0 1 898
box 0 0 96 799
use and2 g8079
timestamp 1386234845
transform 1 0 20019 0 1 898
box 0 0 120 799
use and2 g7999
timestamp 1386234845
transform 1 0 20139 0 1 898
box 0 0 120 799
use nand4 g8239
timestamp 1386234936
transform 1 0 20259 0 1 898
box 0 0 144 799
use inv g8007
timestamp 1386238110
transform 1 0 20403 0 1 898
box 0 0 120 799
use nand2 g7965
timestamp 1386234792
transform 1 0 20523 0 1 898
box 0 0 96 799
use nand2 g8109
timestamp 1386234792
transform 1 0 20619 0 1 898
box 0 0 96 799
use nand2 g8085
timestamp 1386234792
transform 1 0 20715 0 1 898
box 0 0 96 799
use and2 g7944
timestamp 1386234845
transform 1 0 20811 0 1 898
box 0 0 120 799
use and2 g8021
timestamp 1386234845
transform 1 0 20931 0 1 898
box 0 0 120 799
use nand2 g7961
timestamp 1386234792
transform 1 0 21051 0 1 898
box 0 0 96 799
use nor2 g7931
timestamp 1386235306
transform 1 0 21147 0 1 898
box 0 0 120 799
use nand4 g7938
timestamp 1386234936
transform 1 0 21267 0 1 898
box 0 0 144 799
use inv g8184
timestamp 1386238110
transform 1 0 21411 0 1 898
box 0 0 120 799
use xor2 g8132
timestamp 1386237344
transform 1 0 21531 0 1 898
box 0 0 192 799
use inv g7902
timestamp 1386238110
transform 1 0 21723 0 1 898
box 0 0 120 799
use nand2 g8219
timestamp 1386234792
transform 1 0 21843 0 1 898
box 0 0 96 799
use nand2 g7916
timestamp 1386234792
transform 1 0 21939 0 1 898
box 0 0 96 799
use nor2 g8061
timestamp 1386235306
transform 1 0 22035 0 1 898
box 0 0 120 799
use and2 g8115
timestamp 1386234845
transform 1 0 22155 0 1 898
box 0 0 120 799
use nand2 g8202
timestamp 1386234792
transform 1 0 22275 0 1 898
box 0 0 96 799
use nand3 g7973
timestamp 1386234893
transform 1 0 22371 0 1 898
box 0 0 120 799
use nor2 g7908
timestamp 1386235306
transform 1 0 22491 0 1 898
box 0 0 120 799
use nand3 g8208
timestamp 1386234893
transform 1 0 22611 0 1 898
box 0 0 120 799
use nand2 g7958
timestamp 1386234792
transform 1 0 22731 0 1 898
box 0 0 96 799
use inv g8156
timestamp 1386238110
transform 1 0 22827 0 1 898
box 0 0 120 799
use nor2 g8231
timestamp 1386235306
transform 1 0 22947 0 1 898
box 0 0 120 799
use nor2 g8047
timestamp 1386235306
transform 1 0 23067 0 1 898
box 0 0 120 799
use nand2 g7992
timestamp 1386234792
transform 1 0 23187 0 1 898
box 0 0 96 799
use nand3 g7957
timestamp 1386234893
transform 1 0 23283 0 1 898
box 0 0 120 799
use nand4 g8179
timestamp 1386234936
transform 1 0 23403 0 1 898
box 0 0 144 799
use nand3 g8022
timestamp 1386234893
transform 1 0 23547 0 1 898
box 0 0 120 799
use and2 g8193
timestamp 1386234845
transform 1 0 23667 0 1 898
box 0 0 120 799
use nand2 g8071
timestamp 1386234792
transform 1 0 23787 0 1 898
box 0 0 96 799
use nand3 g7953
timestamp 1386234893
transform 1 0 23883 0 1 898
box 0 0 120 799
use nand4 g8083
timestamp 1386234936
transform 1 0 24003 0 1 898
box 0 0 144 799
use nand3 g8204
timestamp 1386234893
transform 1 0 24147 0 1 898
box 0 0 120 799
use nand2 g8053
timestamp 1386234792
transform 1 0 24267 0 1 898
box 0 0 96 799
use nand2 g8000
timestamp 1386234792
transform 1 0 24363 0 1 898
box 0 0 96 799
use nand2 state_reg_91_0_93_
timestamp 1386234792
transform 1 0 24459 0 1 898
box 0 0 96 799
use scandtype g8142
timestamp 1386241841
transform 1 0 24555 0 1 898
box 0 0 624 799
use nand2 g7891
timestamp 1386234792
transform 1 0 25179 0 1 898
box 0 0 96 799
use nand4 stateSub_reg_91_1_93_
timestamp 1386234936
transform 1 0 25275 0 1 898
box 0 0 144 799
use scandtype SysBus_91_1_93_
timestamp 1386241841
transform 1 0 25419 0 1 898
box 0 0 624 799
use rowcrosser nIRQ
timestamp 1386086759
transform 1 0 26043 0 1 898
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 26091 0 1 898
box 0 0 320 799
<< labels >>
rlabel m2contact 26121 4258 26121 4258 6 RwSel[0]
rlabel m2contact 26121 1738 26121 1738 6 RwSel[0]
rlabel m2contact 26097 4762 26097 4762 6 RwSel[1]
rlabel m2contact 26097 1714 26097 1714 6 RwSel[1]
rlabel m2contact 26073 3562 26073 3562 6 ENB
rlabel m2contact 25929 6466 25929 6466 6 stateSub[1]
rlabel m2contact 25881 5410 25881 5410 6 n_66
rlabel m2contact 25737 2146 25737 2146 6 Flags[1]
rlabel m2contact 25689 2506 25689 2506 6 StatusRegEn
rlabel m2contact 25617 5098 25617 5098 6 n_42
rlabel m2contact 25569 2002 25569 2002 6 OpcodeCondIn[6]
rlabel m2contact 25521 2962 25521 2962 6 n_196
rlabel m2contact 25497 4954 25497 4954 6 n_197
rlabel m2contact 25473 4138 25473 4138 6 n_254
rlabel m2contact 25449 6466 25449 6466 6 stateSub[1]
rlabel m2contact 25449 4282 25449 4282 6 stateSub[1]
rlabel m2contact 25425 6442 25425 6442 6 n_40
rlabel m2contact 25401 4258 25401 4258 6 RwSel[0]
rlabel m2contact 25377 4282 25377 4282 6 stateSub[1]
rlabel m2contact 25377 5098 25377 5098 6 n_42
rlabel m2contact 25353 2314 25353 2314 6 n_255
rlabel m2contact 25329 2626 25329 2626 6 n_339
rlabel m2contact 25305 6634 25305 6634 6 n_212
rlabel m2contact 25281 4930 25281 4930 6 n_293
rlabel m2contact 25257 5026 25257 5026 6 n_271
rlabel m2contact 25257 1714 25257 1714 6 n_271
rlabel m2contact 25233 5026 25233 5026 6 n_271
rlabel m2contact 25233 5002 25233 5002 6 n_59
rlabel m2contact 25209 3130 25209 3130 6 state[0]
rlabel m2contact 25185 3010 25185 3010 6 n_231
rlabel m2contact 25161 3538 25161 3538 6 n_192
rlabel m2contact 25137 4570 25137 4570 6 n_157
rlabel m2contact 25101 4282 25101 4282 6 n_339
rlabel m2contact 25101 2626 25101 2626 6 n_339
rlabel m2contact 25089 4306 25089 4306 6 Rs1Sel[0]
rlabel m2contact 25065 4282 25065 4282 6 n_339
rlabel m2contact 25065 3130 25065 3130 6 state[0]
rlabel m2contact 25041 2194 25041 2194 6 n_319
rlabel m2contact 25017 5458 25017 5458 6 n_229
rlabel m2contact 25017 3274 25017 3274 6 n_100
rlabel m2contact 24993 3826 24993 3826 6 n_326
rlabel m2contact 24945 5242 24945 5242 6 n_355
rlabel m2contact 24921 5674 24921 5674 6 n_287
rlabel m2contact 24897 6298 24897 6298 6 n_331
rlabel m2contact 24873 6778 24873 6778 6 n_299
rlabel m2contact 24825 2434 24825 2434 6 n_7
rlabel m2contact 24801 5866 24801 5866 6 OpcodeCondIn[0]
rlabel m2contact 24777 3034 24777 3034 6 OpcodeCondIn[7]
rlabel m2contact 24729 4210 24729 4210 6 n_55
rlabel m2contact 24705 2866 24705 2866 6 n_188
rlabel m2contact 24681 5050 24681 5050 6 n_90
rlabel m2contact 24657 6010 24657 6010 6 StatusReg[0]
rlabel m2contact 24657 4306 24657 4306 6 StatusReg[0]
rlabel m2contact 24633 4354 24633 4354 6 n_67
rlabel m2contact 24609 5122 24609 5122 6 n_65
rlabel m2contact 24585 3130 24585 3130 6 state[0]
rlabel m2contact 24561 5410 24561 5410 6 n_66
rlabel m2contact 24537 4114 24537 4114 6 n_242
rlabel m2contact 24537 3442 24537 3442 6 n_242
rlabel m2contact 24537 5962 24537 5962 6 n_151
rlabel m2contact 24537 4234 24537 4234 6 n_151
rlabel m2contact 24513 3442 24513 3442 6 n_242
rlabel m2contact 24513 3466 24513 3466 6 n_302
rlabel m2contact 24489 6010 24489 6010 6 StatusReg[0]
rlabel m2contact 24489 5986 24489 5986 6 n_120
rlabel m2contact 24465 2482 24465 2482 6 n_298
rlabel m2contact 24441 4546 24441 4546 6 n_266
rlabel m2contact 24441 2218 24441 2218 6 n_266
rlabel m2contact 24417 4690 24417 4690 6 n_201
rlabel m2contact 24393 5626 24393 5626 6 n_141
rlabel m2contact 24393 3754 24393 3754 6 n_198
rlabel m2contact 24369 5434 24369 5434 6 n_270
rlabel m2contact 24345 3874 24345 3874 6 n_303
rlabel m2contact 24321 5386 24321 5386 6 n_349
rlabel m2contact 24297 6562 24297 6562 6 OpcodeCondIn[6]
rlabel m2contact 24297 2002 24297 2002 6 OpcodeCondIn[6]
rlabel m2contact 24273 4282 24273 4282 6 n_31
rlabel m2contact 24249 3442 24249 3442 6 n_68
rlabel m2contact 24225 2002 24225 2002 6 OpcodeCondIn[6]
rlabel m2contact 24225 5818 24225 5818 6 OpcodeCondIn[1]
rlabel m2contact 24201 2698 24201 2698 6 n_37
rlabel m2contact 24201 4258 24201 4258 6 n_35
rlabel m2contact 24177 3730 24177 3730 6 OpcodeCondIn[4]
rlabel m2contact 24153 3946 24153 3946 6 n_263
rlabel m2contact 24129 4570 24129 4570 6 n_157
rlabel m2contact 24129 3922 24129 3922 6 n_157
rlabel m2contact 24105 4210 24105 4210 6 n_55
rlabel m2contact 24105 5746 24105 5746 6 OpcodeCondIn[2]
rlabel m2contact 24081 4234 24081 4234 6 n_151
rlabel m2contact 24081 4810 24081 4810 6 n_262
rlabel m2contact 24057 2098 24057 2098 6 n_80
rlabel m2contact 24033 4378 24033 4378 6 n_329
rlabel m2contact 24009 4330 24009 4330 6 n_318
rlabel m2contact 24009 1882 24009 1882 6 n_318
rlabel m2contact 23985 5074 23985 5074 6 n_166
rlabel m2contact 23985 6082 23985 6082 6 n_330
rlabel m2contact 23961 4234 23961 4234 6 n_214
rlabel m2contact 23937 4546 23937 4546 6 n_266
rlabel m2contact 23937 4522 23937 4522 6 n_248
rlabel m2contact 23913 6370 23913 6370 6 n_74
rlabel m2contact 23913 3130 23913 3130 6 state[0]
rlabel m2contact 23889 5698 23889 5698 6 n_138
rlabel m2contact 23865 3826 23865 3826 6 n_326
rlabel m2contact 23865 4474 23865 4474 6 n_187
rlabel m2contact 23841 4354 23841 4354 6 n_67
rlabel m2contact 23841 2746 23841 2746 6 stateSub[2]
rlabel m2contact 23817 3634 23817 3634 6 n_34
rlabel m2contact 23793 4210 23793 4210 6 n_38
rlabel m2contact 23769 6562 23769 6562 6 OpcodeCondIn[6]
rlabel m2contact 23769 6538 23769 6538 6 n_360
rlabel m2contact 23745 2698 23745 2698 6 n_37
rlabel m2contact 23721 4882 23721 4882 6 n_342
rlabel m2contact 23697 3994 23697 3994 6 n_243
rlabel m2contact 23697 3226 23697 3226 6 n_195
rlabel m2contact 23673 2170 23673 2170 6 n_125
rlabel m2contact 23649 6154 23649 6154 6 n_238
rlabel m2contact 23649 5002 23649 5002 6 n_59
rlabel m2contact 23625 2002 23625 2002 6 OpcodeCondIn[6]
rlabel m2contact 23601 6394 23601 6394 6 n_185
rlabel m2contact 23577 2818 23577 2818 6 OpcodeCondIn[3]
rlabel m2contact 23577 4714 23577 4714 6 n_309
rlabel m2contact 23553 5866 23553 5866 6 OpcodeCondIn[0]
rlabel m2contact 23553 4018 23553 4018 6 OpcodeCondIn[0]
rlabel m2contact 23529 6418 23529 6418 6 n_280
rlabel m2contact 23529 6082 23529 6082 6 n_330
rlabel m2contact 23493 4354 23493 4354 6 n_123
rlabel m2contact 23493 2290 23493 2290 6 n_123
rlabel m2contact 23481 4786 23481 4786 6 n_112
rlabel m2contact 23457 1786 23457 1786 6 n_189
rlabel m2contact 23433 4162 23433 4162 6 n_159
rlabel m2contact 23409 5050 23409 5050 6 n_90
rlabel m2contact 23385 6202 23385 6202 6 n_158
rlabel m2contact 23361 2986 23361 2986 6 n_230
rlabel m2contact 23337 3922 23337 3922 6 n_157
rlabel m2contact 23337 3970 23337 3970 6 n_219
rlabel m2contact 23313 5506 23313 5506 6 n_311
rlabel m2contact 23313 3538 23313 3538 6 n_192
rlabel m2contact 23289 6850 23289 6850 6 n_181
rlabel m2contact 23265 6010 23265 6010 6 n_272
rlabel m2contact 23265 1762 23265 1762 6 n_272
rlabel m2contact 23241 2578 23241 2578 6 n_332
rlabel m2contact 23241 2050 23241 2050 6 n_107
rlabel m2contact 23217 5890 23217 5890 6 n_97
rlabel m2contact 23193 2746 23193 2746 6 stateSub[2]
rlabel m2contact 23169 4330 23169 4330 6 n_318
rlabel m2contact 23169 2122 23169 2122 6 n_10
rlabel m2contact 23133 4330 23133 4330 6 OpcodeCondIn[7]
rlabel m2contact 23133 3034 23133 3034 6 OpcodeCondIn[7]
rlabel m2contact 23121 4354 23121 4354 6 n_123
rlabel m2contact 23121 2818 23121 2818 6 OpcodeCondIn[3]
rlabel m2contact 23097 4330 23097 4330 6 OpcodeCondIn[7]
rlabel m2contact 23097 3274 23097 3274 6 n_100
rlabel m2contact 23073 4546 23073 4546 6 n_111
rlabel m2contact 23049 4450 23049 4450 6 n_160
rlabel m2contact 23049 5938 23049 5938 6 n_96
rlabel m2contact 23025 5842 23025 5842 6 StatusReg[3]
rlabel m2contact 23025 3250 23025 3250 6 StatusReg[3]
rlabel m2contact 23001 4018 23001 4018 6 OpcodeCondIn[0]
rlabel m2contact 23001 4042 23001 4042 6 n_289
rlabel m2contact 22977 6010 22977 6010 6 n_272
rlabel m2contact 22977 5914 22977 5914 6 n_53
rlabel m2contact 22953 4066 22953 4066 6 n_133
rlabel m2contact 22929 4666 22929 4666 6 PcEn
rlabel m2contact 22929 3610 22929 3610 6 PcEn
rlabel m2contact 22905 4330 22905 4330 6 n_22
rlabel m2contact 22881 4738 22881 4738 6 OpcodeCondIn[5]
rlabel m2contact 22857 5098 22857 5098 6 n_42
rlabel m2contact 22833 2386 22833 2386 6 n_9
rlabel m2contact 22809 5818 22809 5818 6 OpcodeCondIn[1]
rlabel m2contact 22809 3154 22809 3154 6 OpcodeCondIn[1]
rlabel m2contact 22785 4306 22785 4306 6 StatusReg[0]
rlabel m2contact 22785 3202 22785 3202 6 StatusReg[0]
rlabel m2contact 22761 3250 22761 3250 6 StatusReg[3]
rlabel m2contact 22761 3298 22761 3298 6 n_249
rlabel m2contact 22737 5266 22737 5266 6 n_81
rlabel m2contact 22737 2026 22737 2026 6 n_81
rlabel m2contact 22713 3610 22713 3610 6 PcEn
rlabel m2contact 22713 3634 22713 3634 6 n_34
rlabel m2contact 22689 6346 22689 6346 6 n_87
rlabel m2contact 22665 3418 22665 3418 6 n_273
rlabel m2contact 22641 1762 22641 1762 6 n_272
rlabel m2contact 22617 4522 22617 4522 6 n_248
rlabel m2contact 22593 3658 22593 3658 6 ALE
rlabel m2contact 22569 3394 22569 3394 6 n_253
rlabel m2contact 22545 5410 22545 5410 6 n_66
rlabel m2contact 22545 3850 22545 3850 6 stateSub[0]
rlabel m2contact 22521 4090 22521 4090 6 n_73
rlabel m2contact 22497 5578 22497 5578 6 n_220
rlabel m2contact 22497 2794 22497 2794 6 n_220
rlabel m2contact 22473 3898 22473 3898 6 n_93
rlabel m2contact 22449 3154 22449 3154 6 OpcodeCondIn[1]
rlabel m2contact 22449 3178 22449 3178 6 n_41
rlabel m2contact 22425 3202 22425 3202 6 StatusReg[0]
rlabel m2contact 22425 3250 22425 3250 6 n_92
rlabel m2contact 22401 5866 22401 5866 6 OpcodeCondIn[0]
rlabel m2contact 22377 2890 22377 2890 6 n_108
rlabel m2contact 22353 2026 22353 2026 6 n_81
rlabel m2contact 22353 2050 22353 2050 6 n_107
rlabel m2contact 22329 6754 22329 6754 6 n_62
rlabel m2contact 22329 2674 22329 2674 6 n_227
rlabel m2contact 22305 2530 22305 2530 6 n_30
rlabel m2contact 22281 4426 22281 4426 6 n_215
rlabel m2contact 22257 2794 22257 2794 6 n_220
rlabel m2contact 22257 2818 22257 2818 6 OpcodeCondIn[3]
rlabel m2contact 22233 3754 22233 3754 6 n_198
rlabel m2contact 22209 4234 22209 4234 6 n_214
rlabel m2contact 22185 3754 22185 3754 6 n_198
rlabel m2contact 22161 2554 22161 2554 6 StatusReg[2]
rlabel m2contact 22137 5146 22137 5146 6 n_172
rlabel m2contact 22137 4498 22137 4498 6 n_172
rlabel m2contact 22113 4066 22113 4066 6 n_133
rlabel m2contact 22089 5026 22089 5026 6 n_118
rlabel m2contact 22065 6466 22065 6466 6 stateSub[1]
rlabel m2contact 22041 5986 22041 5986 6 n_120
rlabel m2contact 22017 6490 22017 6490 6 n_116
rlabel m2contact 21993 4186 21993 4186 6 n_226
rlabel m2contact 21993 3274 21993 3274 6 n_100
rlabel m2contact 21969 5146 21969 5146 6 n_172
rlabel m2contact 21969 5050 21969 5050 6 n_90
rlabel m2contact 21945 4018 21945 4018 6 n_225
rlabel m2contact 21921 6058 21921 6058 6 n_295
rlabel m2contact 21897 2554 21897 2554 6 StatusReg[2]
rlabel m2contact 21873 2482 21873 2482 6 n_298
rlabel m2contact 21849 5770 21849 5770 6 n_176
rlabel m2contact 21825 5650 21825 5650 6 n_177
rlabel m2contact 21801 4642 21801 4642 6 n_162
rlabel m2contact 21777 2410 21777 2410 6 n_277
rlabel m2contact 21753 5266 21753 5266 6 n_81
rlabel m2contact 21753 5218 21753 5218 6 n_126
rlabel m2contact 21729 6178 21729 6178 6 n_275
rlabel m2contact 21681 3922 21681 3922 6 n_19
rlabel m2contact 21681 5218 21681 5218 6 n_126
rlabel m2contact 21657 2818 21657 2818 6 OpcodeCondIn[3]
rlabel m2contact 21633 2050 21633 2050 6 n_107
rlabel m2contact 21585 5818 21585 5818 6 OpcodeCondIn[1]
rlabel m2contact 21561 6802 21561 6802 6 n_164
rlabel m2contact 21561 5866 21561 5866 6 OpcodeCondIn[0]
rlabel m2contact 21537 4594 21537 4594 6 OpcodeCondIn[6]
rlabel m2contact 21537 2002 21537 2002 6 OpcodeCondIn[6]
rlabel m2contact 21513 2794 21513 2794 6 n_246
rlabel m2contact 21489 6010 21489 6010 6 n_325
rlabel m2contact 21465 3802 21465 3802 6 n_15
rlabel m2contact 21441 4594 21441 4594 6 OpcodeCondIn[6]
rlabel m2contact 21441 4402 21441 4402 6 Op1Sel
rlabel m2contact 21417 6394 21417 6394 6 n_185
rlabel m2contact 21393 4354 21393 4354 6 n_327
rlabel m2contact 21369 3826 21369 3826 6 n_326
rlabel m2contact 21345 3898 21345 3898 6 n_93
rlabel m2contact 21345 5986 21345 5986 6 n_120
rlabel m2contact 21297 2914 21297 2914 6 n_70
rlabel m2contact 21249 3874 21249 3874 6 n_303
rlabel m2contact 21249 4570 21249 4570 6 n_157
rlabel m2contact 21225 5290 21225 5290 6 n_282
rlabel m2contact 21225 3898 21225 3898 6 n_282
rlabel m2contact 21201 3946 21201 3946 6 n_263
rlabel m2contact 21201 4786 21201 4786 6 n_112
rlabel m2contact 21177 3898 21177 3898 6 n_282
rlabel m2contact 21177 4138 21177 4138 6 n_254
rlabel m2contact 21153 6034 21153 6034 6 n_193
rlabel m2contact 21153 3946 21153 3946 6 n_193
rlabel m2contact 21129 4594 21129 4594 6 n_291
rlabel m2contact 21105 4978 21105 4978 6 n_88
rlabel m2contact 21105 4882 21105 4882 6 n_342
rlabel m2contact 21081 3946 21081 3946 6 n_193
rlabel m2contact 21081 5338 21081 5338 6 n_259
rlabel m2contact 21009 2338 21009 2338 6 n_102
rlabel m2contact 20985 4546 20985 4546 6 n_111
rlabel m2contact 20961 5314 20961 5314 6 n_94
rlabel m2contact 20913 3586 20913 3586 6 n_114
rlabel m2contact 20889 4834 20889 4834 6 n_1
rlabel m2contact 20841 3346 20841 3346 6 n_113
rlabel m2contact 20841 3826 20841 3826 6 nWait
rlabel m2contact 20793 3610 20793 3610 6 n_64
rlabel m2contact 20769 4858 20769 4858 6 n_17
rlabel m2contact 20745 6658 20745 6658 6 n_63
rlabel m2contact 20697 4306 20697 4306 6 StatusReg[0]
rlabel m2contact 20697 3370 20697 3370 6 n_284
rlabel m2contact 20649 3514 20649 3514 6 n_479
rlabel m2contact 20649 2938 20649 2938 6 n_286
rlabel m2contact 20577 3994 20577 3994 6 n_243
rlabel m2contact 20553 5170 20553 5170 6 n_210
rlabel m2contact 20481 3082 20481 3082 6 n_222
rlabel m2contact 20433 1906 20433 1906 6 n_12
rlabel m2contact 20385 5794 20385 5794 6 n_155
rlabel m2contact 20361 5770 20361 5770 6 n_176
rlabel m2contact 20337 4522 20337 4522 6 n_248
rlabel m2contact 20313 3130 20313 3130 6 state[0]
rlabel m2contact 20289 4234 20289 4234 6 n_214
rlabel m2contact 20289 4306 20289 4306 6 n_358
rlabel m2contact 20241 6586 20241 6586 6 IrWe
rlabel m2contact 20193 3274 20193 3274 6 n_100
rlabel m2contact 20169 4066 20169 4066 6 n_133
rlabel m2contact 20169 5722 20169 5722 6 n_29
rlabel m2contact 20121 5818 20121 5818 6 OpcodeCondIn[1]
rlabel m2contact 20121 5482 20121 5482 6 n_16
rlabel m2contact 20097 4258 20097 4258 6 n_35
rlabel m2contact 20073 3274 20073 3274 6 n_100
rlabel m2contact 20049 3178 20049 3178 6 n_41
rlabel m2contact 20049 4618 20049 4618 6 n_194
rlabel m2contact 20025 6826 20025 6826 6 n_182
rlabel m2contact 20025 4066 20025 4066 6 n_182
rlabel m2contact 20001 4066 20001 4066 6 n_182
rlabel m2contact 20001 4258 20001 4258 6 n_35
rlabel m2contact 19977 5914 19977 5914 6 n_53
rlabel m2contact 19977 5050 19977 5050 6 n_90
rlabel m2contact 19953 4570 19953 4570 6 n_143
rlabel m2contact 19929 4066 19929 4066 6 n_179
rlabel m2contact 19881 6706 19881 6706 6 n_135
rlabel m2contact 19881 2674 19881 2674 6 n_227
rlabel m2contact 19857 3058 19857 3058 6 n_233
rlabel m2contact 19833 2818 19833 2818 6 OpcodeCondIn[3]
rlabel m2contact 19785 1738 19785 1738 6 n_204
rlabel m2contact 19761 6250 19761 6250 6 n_109
rlabel m2contact 19737 5770 19737 5770 6 n_176
rlabel m2contact 19713 2026 19713 2026 6 n_56
rlabel m2contact 19689 4858 19689 4858 6 n_17
rlabel m2contact 19665 4834 19665 4834 6 n_1
rlabel m2contact 19665 1882 19665 1882 6 n_318
rlabel m2contact 19641 3178 19641 3178 6 n_41
rlabel m2contact 19617 4138 19617 4138 6 n_254
rlabel m2contact 19593 2770 19593 2770 6 n_163
rlabel m2contact 19569 4642 19569 4642 6 n_162
rlabel m2contact 19545 5530 19545 5530 6 n_153
rlabel m2contact 19497 4762 19497 4762 6 RwSel[1]
rlabel m2contact 19473 2266 19473 2266 6 n_333
rlabel m2contact 19449 6538 19449 6538 6 n_360
rlabel m2contact 19425 4426 19425 4426 6 n_215
rlabel m2contact 19377 5602 19377 5602 6 n_357
rlabel m2contact 19353 6106 19353 6106 6 n_32
rlabel m2contact 19353 6730 19353 6730 6 n_285
rlabel m2contact 19329 4378 19329 4378 6 n_329
rlabel m2contact 19305 6058 19305 6058 6 n_295
rlabel m2contact 19305 5746 19305 5746 6 OpcodeCondIn[2]
rlabel m2contact 19281 4282 19281 4282 6 n_31
rlabel m2contact 19257 6226 19257 6226 6 n_296
rlabel m2contact 19233 4858 19233 4858 6 n_103
rlabel m2contact 19209 6178 19209 6178 6 n_275
rlabel m2contact 19209 6130 19209 6130 6 n_21
rlabel m2contact 19185 6058 19185 6058 6 n_86
rlabel m2contact 19161 4426 19161 4426 6 n_328
rlabel m2contact 19137 5194 19137 5194 6 n_49
rlabel m2contact 19113 6082 19113 6082 6 n_330
rlabel m2contact 19065 1930 19065 1930 6 n_13
rlabel m2contact 19041 3058 19041 3058 6 n_233
rlabel m2contact 19041 4738 19041 4738 6 OpcodeCondIn[5]
rlabel m2contact 19017 6394 19017 6394 6 n_185
rlabel m2contact 19017 5554 19017 5554 6 n_264
rlabel m2contact 18969 2650 18969 2650 6 n_174
rlabel m2contact 18945 4378 18945 4378 6 n_39
rlabel m2contact 18921 3754 18921 3754 6 n_198
rlabel m2contact 18873 4474 18873 4474 6 n_187
rlabel m2contact 18849 6466 18849 6466 6 stateSub[1]
rlabel m2contact 18825 6562 18825 6562 6 n_147
rlabel m2contact 18777 4378 18777 4378 6 n_39
rlabel m2contact 18753 3154 18753 3154 6 n_281
rlabel m2contact 18729 5146 18729 5146 6 n_57
rlabel m2contact 18681 4762 18681 4762 6 n_79
rlabel m2contact 18633 3178 18633 3178 6 n_41
rlabel m2contact 18609 4546 18609 4546 6 n_111
rlabel m2contact 18585 4018 18585 4018 6 n_225
rlabel m2contact 18585 3946 18585 3946 6 n_225
rlabel m2contact 18561 4474 18561 4474 6 n_216
rlabel m2contact 18561 3202 18561 3202 6 n_216
rlabel m2contact 18537 3538 18537 3538 6 n_192
rlabel m2contact 18513 5266 18513 5266 6 n_9
rlabel m2contact 18513 2386 18513 2386 6 n_9
rlabel m2contact 18489 2170 18489 2170 6 n_125
rlabel m2contact 18465 6610 18465 6610 6 n_3
rlabel m2contact 18441 4906 18441 4906 6 n_203
rlabel m2contact 18417 4690 18417 4690 6 n_201
rlabel m2contact 18393 2602 18393 2602 6 n_202
rlabel m2contact 18357 4378 18357 4378 6 n_56
rlabel m2contact 18357 2026 18357 2026 6 n_56
rlabel m2contact 18345 4882 18345 4882 6 n_342
rlabel m2contact 18321 3946 18321 3946 6 n_225
rlabel m2contact 18321 3994 18321 3994 6 state[1]
rlabel m2contact 18297 3202 18297 3202 6 n_216
rlabel m2contact 18297 3250 18297 3250 6 n_92
rlabel m2contact 18273 2746 18273 2746 6 stateSub[2]
rlabel m2contact 18249 3970 18249 3970 6 n_219
rlabel m2contact 18225 3946 18225 3946 6 n_366
rlabel m2contact 18201 3682 18201 3682 6 n_223
rlabel m2contact 18177 2578 18177 2578 6 n_332
rlabel m2contact 18153 4834 18153 4834 6 n_345
rlabel m2contact 18129 4210 18129 4210 6 n_38
rlabel m2contact 18105 5194 18105 5194 6 n_49
rlabel m2contact 18105 3682 18105 3682 6 n_223
rlabel m2contact 18081 3130 18081 3130 6 state[0]
rlabel m2contact 18057 3634 18057 3634 6 n_34
rlabel m2contact 18033 5194 18033 5194 6 n_321
rlabel m2contact 18009 1834 18009 1834 6 n_115
rlabel m2contact 17985 5362 17985 5362 6 n_306
rlabel m2contact 17961 6106 17961 6106 6 n_32
rlabel m2contact 17937 4210 17937 4210 6 n_75
rlabel m2contact 17937 3778 17937 3778 6 n_161
rlabel m2contact 17913 3538 17913 3538 6 n_192
rlabel m2contact 17889 4666 17889 4666 6 PcEn
rlabel m2contact 17889 4450 17889 4450 6 n_160
rlabel m2contact 17865 6634 17865 6634 6 n_212
rlabel m2contact 17865 3322 17865 3322 6 n_212
rlabel m2contact 17841 3898 17841 3898 6 n_139
rlabel m2contact 17817 3394 17817 3394 6 n_253
rlabel m2contact 17793 3802 17793 3802 6 n_15
rlabel m2contact 17793 3874 17793 3874 6 n_99
rlabel m2contact 17769 4378 17769 4378 6 n_56
rlabel m2contact 17769 2746 17769 2746 6 stateSub[2]
rlabel m2contact 17745 5122 17745 5122 6 n_65
rlabel m2contact 17745 2458 17745 2458 6 n_65
rlabel m2contact 17721 4666 17721 4666 6 n_308
rlabel m2contact 17697 3490 17697 3490 6 n_368
rlabel m2contact 17673 4066 17673 4066 6 n_179
rlabel m2contact 17673 4378 17673 4378 6 n_235
rlabel m2contact 17649 1954 17649 1954 6 n_228
rlabel m2contact 17625 6538 17625 6538 6 n_360
rlabel m2contact 17601 3058 17601 3058 6 n_233
rlabel m2contact 17577 5122 17577 5122 6 n_65
rlabel m2contact 17553 5266 17553 5266 6 n_9
rlabel m2contact 17553 3730 17553 3730 6 OpcodeCondIn[4]
rlabel m2contact 17529 2722 17529 2722 6 n_130
rlabel m2contact 17529 3154 17529 3154 6 n_281
rlabel m2contact 17505 5266 17505 5266 6 n_26
rlabel m2contact 17505 3202 17505 3202 6 n_26
rlabel m2contact 17481 1762 17481 1762 6 n_272
rlabel m2contact 17481 1810 17481 1810 6 n_237
rlabel m2contact 17457 2842 17457 2842 6 n_142
rlabel m2contact 17457 4162 17457 4162 6 n_159
rlabel m2contact 17433 3130 17433 3130 6 state[0]
rlabel m2contact 17433 3538 17433 3538 6 n_192
rlabel m2contact 17409 1810 17409 1810 6 n_237
rlabel m2contact 17385 5674 17385 5674 6 n_287
rlabel m2contact 17361 3322 17361 3322 6 n_212
rlabel m2contact 17361 3706 17361 3706 6 SysBus[1]
rlabel m2contact 17337 2458 17337 2458 6 n_65
rlabel m2contact 17337 2938 17337 2938 6 n_286
rlabel m2contact 17313 3130 17313 3130 6 state[0]
rlabel m2contact 17289 4522 17289 4522 6 n_248
rlabel m2contact 17265 6658 17265 6658 6 n_63
rlabel m2contact 17241 3178 17241 3178 6 n_41
rlabel m2contact 17217 5050 17217 5050 6 n_90
rlabel m2contact 17193 6130 17193 6130 6 n_21
rlabel m2contact 17169 1978 17169 1978 6 n_250
rlabel m2contact 17145 2794 17145 2794 6 n_246
rlabel m2contact 17121 4522 17121 4522 6 n_248
rlabel m2contact 17121 3730 17121 3730 6 OpcodeCondIn[4]
rlabel m2contact 17097 3202 17097 3202 6 n_26
rlabel m2contact 17097 3298 17097 3298 6 n_249
rlabel m2contact 17049 5506 17049 5506 6 n_311
rlabel m2contact 17049 1762 17049 1762 6 SysBus[2]
rlabel m2contact 17025 3154 17025 3154 6 n_281
rlabel m2contact 17001 3322 17001 3322 6 n_77
rlabel m2contact 17001 4714 17001 4714 6 n_309
rlabel m2contact 16953 4618 16953 4618 6 n_194
rlabel m2contact 16857 3154 16857 3154 6 n_281
rlabel m2contact 16833 5290 16833 5290 6 n_282
rlabel m2contact 16785 4210 16785 4210 6 n_75
rlabel m2contact 16737 4162 16737 4162 6 n_159
rlabel m2contact 16617 5506 16617 5506 6 n_82
rlabel m2contact 16521 2362 16521 2362 6 n_244
rlabel m2contact 16497 3298 16497 3298 6 n_249
rlabel m2contact 16473 2626 16473 2626 6 n_339
rlabel m2contact 16449 5242 16449 5242 6 n_355
rlabel m2contact 16449 2746 16449 2746 6 stateSub[2]
rlabel m2contact 16377 2818 16377 2818 6 OpcodeCondIn[3]
rlabel m2contact 16329 4546 16329 4546 6 n_111
rlabel m2contact 16305 5266 16305 5266 6 n_26
rlabel m2contact 16281 2818 16281 2818 6 OpcodeCondIn[3]
rlabel m2contact 16281 3274 16281 3274 6 n_100
rlabel m2contact 16257 5410 16257 5410 6 n_66
rlabel m2contact 16257 3034 16257 3034 6 OpcodeCondIn[7]
rlabel m2contact 16209 5026 16209 5026 6 n_118
rlabel m2contact 16185 6490 16185 6490 6 n_116
rlabel m2contact 16161 2074 16161 2074 6 n_117
rlabel m2contact 16113 6682 16113 6682 6 n_124
rlabel m2contact 16065 3106 16065 3106 6 n_76
rlabel m2contact 16041 2290 16041 2290 6 n_123
rlabel m2contact 15969 3754 15969 3754 6 n_198
rlabel m2contact 15921 2722 15921 2722 6 n_130
rlabel m2contact 15873 4834 15873 4834 6 n_345
rlabel m2contact 15849 5674 15849 5674 6 n_247
rlabel m2contact 15825 4666 15825 4666 6 n_308
rlabel m2contact 15801 6106 15801 6106 6 n_294
rlabel m2contact 15777 2458 15777 2458 6 n_221
rlabel m2contact 15705 4498 15705 4498 6 n_172
rlabel m2contact 15681 5242 15681 5242 6 n_253
rlabel m2contact 15681 3394 15681 3394 6 n_253
rlabel m2contact 15657 5026 15657 5026 6 n_171
rlabel m2contact 15633 4666 15633 4666 6 n_227
rlabel m2contact 15633 2674 15633 2674 6 n_227
rlabel m2contact 15609 4210 15609 4210 6 n_51
rlabel m2contact 15585 5146 15585 5146 6 n_57
rlabel m2contact 15561 3202 15561 3202 6 n_245
rlabel m2contact 15561 4834 15561 4834 6 n_24
rlabel m2contact 15537 6466 15537 6466 6 stateSub[1]
rlabel m2contact 15537 4498 15537 4498 6 stateSub[1]
rlabel m2contact 15513 5962 15513 5962 6 n_151
rlabel m2contact 15513 4066 15513 4066 6 n_314
rlabel m2contact 15489 3034 15489 3034 6 OpcodeCondIn[7]
rlabel m2contact 15465 2242 15465 2242 6 n_129
rlabel m2contact 15441 3538 15441 3538 6 n_192
rlabel m2contact 15417 3754 15417 3754 6 n_198
rlabel m2contact 15417 3802 15417 3802 6 nOE
rlabel m2contact 15393 5242 15393 5242 6 n_253
rlabel m2contact 15393 4618 15393 4618 6 n_194
rlabel m2contact 15369 5194 15369 5194 6 n_321
rlabel m2contact 15345 5074 15345 5074 6 n_166
rlabel m2contact 15321 2314 15321 2314 6 n_255
rlabel m2contact 15321 5314 15321 5314 6 n_94
rlabel m2contact 15297 4186 15297 4186 6 n_226
rlabel m2contact 15273 3970 15273 3970 6 n_110
rlabel m2contact 15249 4666 15249 4666 6 n_227
rlabel m2contact 15249 4186 15249 4186 6 n_131
rlabel m2contact 15225 6250 15225 6250 6 n_109
rlabel m2contact 15201 4498 15201 4498 6 stateSub[1]
rlabel m2contact 15201 4690 15201 4690 6 n_201
rlabel m2contact 15177 5314 15177 5314 6 n_94
rlabel m2contact 15153 4474 15153 4474 6 n_216
rlabel m2contact 15129 5026 15129 5026 6 n_171
rlabel m2contact 15105 1810 15105 1810 6 n_237
rlabel m2contact 15105 2746 15105 2746 6 stateSub[2]
rlabel m2contact 15081 6154 15081 6154 6 n_238
rlabel m2contact 15057 6514 15057 6514 6 n_353
rlabel m2contact 15033 4450 15033 4450 6 n_160
rlabel m2contact 15009 2698 15009 2698 6 n_37
rlabel m2contact 15009 4474 15009 4474 6 n_322
rlabel m2contact 14913 2818 14913 2818 6 OpcodeCondIn[3]
rlabel m2contact 14889 4738 14889 4738 6 OpcodeCondIn[5]
rlabel m2contact 14865 2746 14865 2746 6 stateSub[2]
rlabel m2contact 14817 5050 14817 5050 6 n_90
rlabel m2contact 14817 3082 14817 3082 6 n_222
rlabel m2contact 14793 3058 14793 3058 6 n_233
rlabel m2contact 14745 4162 14745 4162 6 n_159
rlabel m2contact 14697 5866 14697 5866 6 OpcodeCondIn[0]
rlabel m2contact 14673 5818 14673 5818 6 OpcodeCondIn[1]
rlabel m2contact 14625 5170 14625 5170 6 n_210
rlabel m2contact 14577 3130 14577 3130 6 state[0]
rlabel m2contact 14553 6250 14553 6250 6 n_109
rlabel m2contact 14481 5746 14481 5746 6 OpcodeCondIn[2]
rlabel m2contact 14457 3514 14457 3514 6 n_479
rlabel m2contact 14457 4354 14457 4354 6 n_327
rlabel m2contact 14433 4282 14433 4282 6 n_31
rlabel m2contact 14385 6418 14385 6418 6 n_280
rlabel m2contact 14385 4282 14385 4282 6 n_280
rlabel m2contact 14361 4882 14361 4882 6 n_342
rlabel m2contact 14337 3946 14337 3946 6 n_366
rlabel m2contact 14313 4282 14313 4282 6 n_280
rlabel m2contact 14313 5386 14313 5386 6 n_349
rlabel m2contact 14289 4498 14289 4498 6 n_323
rlabel m2contact 14241 4282 14241 4282 6 n_208
rlabel m2contact 14217 1738 14217 1738 6 n_204
rlabel m2contact 14193 5650 14193 5650 6 n_177
rlabel m2contact 14157 4666 14157 4666 6 n_481
rlabel m2contact 14157 3514 14157 3514 6 n_481
rlabel m2contact 14145 5842 14145 5842 6 StatusReg[3]
rlabel m2contact 14121 3346 14121 3346 6 n_113
rlabel m2contact 14097 4666 14097 4666 6 n_481
rlabel m2contact 14097 4522 14097 4522 6 n_248
rlabel m2contact 14073 3298 14073 3298 6 n_249
rlabel m2contact 13977 6322 13977 6322 6 n_6
rlabel m2contact 13953 3946 13953 3946 6 n_258
rlabel m2contact 13833 6082 13833 6082 6 n_330
rlabel m2contact 13737 4354 13737 4354 6 n_137
rlabel m2contact 13737 4450 13737 4450 6 n_365
rlabel m2contact 13713 2890 13713 2890 6 n_108
rlabel m2contact 13641 2674 13641 2674 6 n_227
rlabel m2contact 13617 5242 13617 5242 6 n_95
rlabel m2contact 13617 4546 13617 4546 6 n_111
rlabel m2contact 13593 5194 13593 5194 4 n_8
rlabel m2contact 13569 4666 13569 4666 4 n_190
rlabel m2contact 13545 6274 13545 6274 4 n_240
rlabel m2contact 13545 2890 13545 2890 4 n_240
rlabel m2contact 13521 3394 13521 3394 4 n_253
rlabel m2contact 13521 5386 13521 5386 4 n_349
rlabel m2contact 13497 2890 13497 2890 4 n_240
rlabel m2contact 13497 3298 13497 3298 4 n_249
rlabel m2contact 13473 2338 13473 2338 4 n_102
rlabel m2contact 13449 5074 13449 5074 4 n_206
rlabel m2contact 13425 4114 13425 4114 4 n_242
rlabel m2contact 13425 1738 13425 1738 4 n_204
rlabel m2contact 13401 6802 13401 6802 4 n_164
rlabel m2contact 13401 5962 13401 5962 4 n_205
rlabel m2contact 13377 3130 13377 3130 4 state[0]
rlabel m2contact 13353 6802 13353 6802 4 n_188
rlabel m2contact 13353 2866 13353 2866 4 n_188
rlabel m2contact 13329 6850 13329 6850 4 n_181
rlabel m2contact 13329 6826 13329 6826 4 n_182
rlabel m2contact 13305 2890 13305 2890 4 n_180
rlabel m2contact 13281 2914 13281 2914 4 n_70
rlabel m2contact 13281 3754 13281 3754 4 n_198
rlabel m2contact 13257 6802 13257 6802 4 n_188
rlabel m2contact 13257 4114 13257 4114 4 n_69
rlabel m2contact 13209 6370 13209 6370 4 n_74
rlabel m2contact 13185 3514 13185 3514 4 n_481
rlabel m2contact 13185 4858 13185 4858 4 n_103
rlabel m2contact 13161 2554 13161 2554 4 StatusReg[2]
rlabel m2contact 13161 3850 13161 3850 4 stateSub[0]
rlabel m2contact 13089 6154 13089 6154 4 n_238
rlabel m2contact 13089 3850 13089 3850 4 stateSub[0]
rlabel m2contact 13065 2746 13065 2746 4 stateSub[2]
rlabel m2contact 13041 4954 13041 4954 4 n_197
rlabel m2contact 12993 3418 12993 3418 4 n_273
rlabel m2contact 12993 3514 12993 3514 4 MemEn
rlabel m2contact 12921 3514 12921 3514 4 MemEn
rlabel m2contact 12921 5194 12921 5194 4 n_8
rlabel m2contact 12897 4810 12897 4810 4 n_262
rlabel m2contact 12873 4162 12873 4162 4 n_159
rlabel m2contact 12873 4066 12873 4066 4 n_314
rlabel m2contact 12849 5194 12849 5194 4 n_230
rlabel m2contact 12849 2986 12849 2986 4 n_230
rlabel m2contact 12825 3418 12825 3418 4 n_121
rlabel m2contact 12801 1810 12801 1810 4 n_11
rlabel m2contact 12801 2818 12801 2818 4 OpcodeCondIn[3]
rlabel m2contact 12777 5986 12777 5986 4 n_120
rlabel m2contact 12777 3034 12777 3034 4 OpcodeCondIn[7]
rlabel m2contact 12753 3130 12753 3130 4 state[0]
rlabel m2contact 12729 5194 12729 5194 4 n_230
rlabel m2contact 12729 3730 12729 3730 4 OpcodeCondIn[4]
rlabel m2contact 12657 5722 12657 5722 4 n_29
rlabel m2contact 12609 6154 12609 6154 4 n_199
rlabel m2contact 12609 3394 12609 3394 4 n_199
rlabel m2contact 12585 6802 12585 6802 4 n_230
rlabel m2contact 12585 2986 12585 2986 4 n_230
rlabel m2contact 12561 1714 12561 1714 4 n_271
rlabel m2contact 12561 2698 12561 2698 4 n_183
rlabel m2contact 12537 6370 12537 6370 4 n_144
rlabel m2contact 12537 3514 12537 3514 4 n_173
rlabel m2contact 12513 6826 12513 6826 4 n_182
rlabel m2contact 12513 5194 12513 5194 4 n_156
rlabel m2contact 12489 5986 12489 5986 4 n_207
rlabel m2contact 12465 3394 12465 3394 4 n_199
rlabel m2contact 12465 4834 12465 4834 4 n_24
rlabel m2contact 12441 3034 12441 3034 4 OpcodeCondIn[7]
rlabel m2contact 12417 2674 12417 2674 4 n_227
rlabel m2contact 12393 4882 12393 4882 4 n_342
rlabel m2contact 12369 5914 12369 5914 4 n_53
rlabel m2contact 12345 5818 12345 5818 4 OpcodeCondIn[1]
rlabel m2contact 12321 6802 12321 6802 4 n_230
rlabel m2contact 12321 3010 12321 3010 4 n_231
rlabel m2contact 12297 6394 12297 6394 4 n_185
rlabel m2contact 12297 3394 12297 3394 4 n_185
rlabel m2contact 12273 6418 12273 6418 4 n_280
rlabel m2contact 12249 2674 12249 2674 4 n_227
rlabel m2contact 12249 2866 12249 2866 4 n_188
rlabel m2contact 12225 3682 12225 3682 4 n_223
rlabel m2contact 12201 3394 12201 3394 4 n_185
rlabel m2contact 12201 5146 12201 5146 4 n_57
rlabel m2contact 12165 3394 12165 3394 4 OpcodeCondIn[6]
rlabel m2contact 12165 2002 12165 2002 4 OpcodeCondIn[6]
rlabel m2contact 12153 6418 12153 6418 4 n_84
rlabel m2contact 12129 3394 12129 3394 4 OpcodeCondIn[6]
rlabel m2contact 12129 2602 12129 2602 4 n_202
rlabel m2contact 12105 2890 12105 2890 4 n_180
rlabel m2contact 12081 3394 12081 3394 4 n_140
rlabel m2contact 12057 6778 12057 6778 4 n_299
rlabel m2contact 12033 6754 12033 6754 4 n_62
rlabel m2contact 12009 1738 12009 1738 4 n_204
rlabel m2contact 12009 2482 12009 2482 4 n_298
rlabel m2contact 11985 4786 11985 4786 4 n_112
rlabel m2contact 11937 2050 11937 2050 4 n_107
rlabel m2contact 11889 6418 11889 6418 4 n_84
rlabel m2contact 11841 6730 11841 6730 4 n_285
rlabel m2contact 11817 1762 11817 1762 4 SysBus[2]
rlabel m2contact 11793 2938 11793 2938 4 n_286
rlabel m2contact 11745 1786 11745 1786 4 n_189
rlabel m2contact 11721 3154 11721 3154 4 n_281
rlabel m2contact 11697 3754 11697 3754 4 n_198
rlabel m2contact 11673 2866 11673 2866 4 n_188
rlabel m2contact 11625 5458 11625 5458 4 n_229
rlabel m2contact 11577 1810 11577 1810 4 n_11
rlabel m2contact 11553 5458 11553 5458 4 n_168
rlabel m2contact 11481 4090 11481 4090 4 n_73
rlabel m2contact 11433 6490 11433 6490 4 n_116
rlabel m2contact 11385 6706 11385 6706 4 n_135
rlabel m2contact 11361 3154 11361 3154 4 n_281
rlabel m2contact 11337 3322 11337 3322 4 n_77
rlabel m2contact 11313 5002 11313 5002 4 n_59
rlabel m2contact 11265 5002 11265 5002 4 n_104
rlabel m2contact 11241 2050 11241 2050 4 n_107
rlabel m2contact 11217 4858 11217 4858 4 n_103
rlabel m2contact 11193 6394 11193 6394 4 n_185
rlabel m2contact 11145 3034 11145 3034 4 OpcodeCondIn[7]
rlabel m2contact 11145 3850 11145 3850 4 stateSub[0]
rlabel m2contact 11121 6682 11121 6682 4 n_124
rlabel m2contact 11097 6658 11097 6658 4 n_63
rlabel m2contact 11097 3322 11097 3322 4 n_175
rlabel m2contact 11073 6634 11073 6634 4 n_212
rlabel m2contact 11049 1834 11049 1834 4 n_115
rlabel m2contact 11025 4570 11025 4570 4 n_143
rlabel m2contact 10977 3346 10977 3346 4 n_113
rlabel m2contact 10953 4546 10953 4546 4 n_111
rlabel m2contact 10929 4690 10929 4690 4 n_201
rlabel m2contact 10905 5554 10905 5554 4 n_264
rlabel m2contact 10905 5170 10905 5170 4 n_210
rlabel m2contact 10881 3946 10881 3946 4 n_258
rlabel m2contact 10857 2986 10857 2986 4 n_230
rlabel m2contact 10833 3706 10833 3706 4 SysBus[1]
rlabel m2contact 10833 3922 10833 3922 4 n_19
rlabel m2contact 10785 5506 10785 5506 4 n_82
rlabel m2contact 10737 5410 10737 5410 4 n_66
rlabel m2contact 10737 3850 10737 3850 4 stateSub[0]
rlabel m2contact 10713 5506 10713 5506 4 n_33
rlabel m2contact 10677 4234 10677 4234 4 n_214
rlabel m2contact 10677 1834 10677 1834 4 n_214
rlabel m2contact 10665 4378 10665 4378 4 n_235
rlabel m2contact 10641 4234 10641 4234 4 n_214
rlabel m2contact 10641 2866 10641 2866 4 n_188
rlabel m2contact 10617 4378 10617 4378 4 n_149
rlabel m2contact 10617 3754 10617 3754 4 n_198
rlabel m2contact 10593 6394 10593 6394 4 n_185
rlabel m2contact 10593 3922 10593 3922 4 n_185
rlabel m2contact 10569 1834 10569 1834 4 n_214
rlabel m2contact 10569 2842 10569 2842 4 n_142
rlabel m2contact 10545 5098 10545 5098 4 n_42
rlabel m2contact 10521 3922 10521 3922 4 n_185
rlabel m2contact 10521 4690 10521 4690 4 n_201
rlabel m2contact 10497 2050 10497 2050 4 n_107
rlabel m2contact 10473 4354 10473 4354 4 n_137
rlabel m2contact 10449 3034 10449 3034 4 OpcodeCondIn[7]
rlabel m2contact 10425 3274 10425 3274 4 n_100
rlabel m2contact 10425 4354 10425 4354 4 n_85
rlabel m2contact 10401 6250 10401 6250 4 n_109
rlabel m2contact 10377 3706 10377 3706 4 ImmSel
rlabel m2contact 10353 1858 10353 1858 4 Rs1Sel[1]
rlabel m2contact 10353 6538 10353 6538 4 n_360
rlabel m2contact 10353 3922 10353 3922 4 n_360
rlabel m2contact 10329 1882 10329 1882 4 n_318
rlabel m2contact 10329 4978 10329 4978 4 n_88
rlabel m2contact 10305 3994 10305 3994 4 state[1]
rlabel m2contact 10281 3922 10281 3922 4 n_360
rlabel m2contact 10281 6346 10281 6346 4 n_87
rlabel m2contact 10233 4978 10233 4978 4 n_145
rlabel m2contact 10233 1882 10233 1882 4 n_145
rlabel m2contact 10209 1882 10209 1882 4 n_145
rlabel m2contact 10209 3922 10209 3922 4 n_241
rlabel m2contact 10185 3730 10185 3730 4 OpcodeCondIn[4]
rlabel m2contact 10161 6274 10161 6274 4 n_240
rlabel m2contact 10161 3154 10161 3154 4 n_281
rlabel m2contact 10137 2002 10137 2002 4 OpcodeCondIn[6]
rlabel m2contact 10137 1882 10137 1882 4 OpcodeCondIn[6]
rlabel m2contact 10113 1882 10113 1882 4 OpcodeCondIn[6]
rlabel m2contact 10113 1906 10113 1906 4 n_12
rlabel m2contact 10089 4738 10089 4738 4 OpcodeCondIn[5]
rlabel m2contact 10065 2002 10065 2002 4 OpcodeCondIn[6]
rlabel m2contact 10041 2266 10041 2266 4 n_333
rlabel m2contact 10017 5458 10017 5458 4 n_168
rlabel m2contact 9993 2578 9993 2578 4 n_332
rlabel m2contact 9993 3154 9993 3154 4 n_281
rlabel m2contact 9969 2266 9969 2266 4 n_128
rlabel m2contact 9945 2578 9945 2578 4 n_122
rlabel m2contact 9921 1906 9921 1906 4 n_12
rlabel m2contact 9921 2002 9921 2002 4 n_363
rlabel m2contact 9897 5794 9897 5794 4 n_155
rlabel m2contact 9897 5458 9897 5458 4 n_25
rlabel m2contact 9873 6010 9873 6010 4 n_325
rlabel m2contact 9849 1930 9849 1930 4 n_13
rlabel m2contact 9849 5794 9849 5794 4 n_232
rlabel m2contact 9825 6010 9825 6010 4 n_211
rlabel m2contact 9777 4882 9777 4882 4 n_342
rlabel m2contact 9753 4474 9753 4474 4 n_322
rlabel m2contact 9705 6226 9705 6226 4 n_296
rlabel m2contact 9681 3634 9681 3634 4 n_34
rlabel m2contact 9657 6466 9657 6466 4 stateSub[1]
rlabel m2contact 9633 6610 9633 6610 4 n_3
rlabel m2contact 9633 3946 9633 3946 4 n_258
rlabel m2contact 9585 3634 9585 3634 4 nIRQ
rlabel m2contact 9561 6394 9561 6394 4 n_185
rlabel m2contact 9537 6586 9537 6586 4 IrWe
rlabel m2contact 9537 3754 9537 3754 4 n_198
rlabel m2contact 9513 5122 9513 5122 4 n_65
rlabel m2contact 9465 1954 9465 1954 4 n_228
rlabel m2contact 9465 5074 9465 5074 4 n_206
rlabel m2contact 9441 6514 9441 6514 4 n_353
rlabel m2contact 9441 2674 9441 2674 4 n_227
rlabel m2contact 9417 2602 9417 2602 4 n_202
rlabel m2contact 9393 6562 9393 6562 4 n_147
rlabel m2contact 9393 4690 9393 4690 4 n_201
rlabel m2contact 9369 5074 9369 5074 4 n_91
rlabel m2contact 9345 2074 9345 2074 4 n_117
rlabel m2contact 9321 1978 9321 1978 4 n_250
rlabel m2contact 9321 6490 9321 6490 4 n_116
rlabel m2contact 9297 2602 9297 2602 4 n_265
rlabel m2contact 9273 6490 9273 6490 4 n_105
rlabel m2contact 9249 3490 9249 3490 4 n_368
rlabel m2contact 9225 1978 9225 1978 4 n_367
rlabel m2contact 9201 6538 9201 6538 4 n_360
rlabel m2contact 9201 3490 9201 3490 4 n_368
rlabel m2contact 9177 5242 9177 5242 4 n_95
rlabel m2contact 9153 3754 9153 3754 4 n_198
rlabel m2contact 9129 5386 9129 5386 4 n_349
rlabel m2contact 9129 5242 9129 5242 4 n_200
rlabel m2contact 9105 6514 9105 6514 4 n_353
rlabel m2contact 9081 1978 9081 1978 4 n_367
rlabel m2contact 9081 6202 9081 6202 4 n_158
rlabel m2contact 9033 6202 9033 6202 4 n_36
rlabel m2contact 9033 4186 9033 4186 4 n_131
rlabel m2contact 9009 2002 9009 2002 4 n_363
rlabel m2contact 9009 4258 9009 4258 4 n_35
rlabel m2contact 8985 2314 8985 2314 4 n_255
rlabel m2contact 8961 2026 8961 2026 4 n_56
rlabel m2contact 8937 6490 8937 6490 4 n_105
rlabel m2contact 8937 5410 8937 5410 4 n_66
rlabel m2contact 8913 6466 8913 6466 4 stateSub[1]
rlabel m2contact 8913 4522 8913 4522 4 n_248
rlabel m2contact 8889 2338 8889 2338 4 n_102
rlabel m2contact 8865 2170 8865 2170 4 n_125
rlabel m2contact 8841 2338 8841 2338 4 n_83
rlabel m2contact 8817 2050 8817 2050 4 n_107
rlabel m2contact 8817 4738 8817 4738 4 OpcodeCondIn[5]
rlabel m2contact 8793 2170 8793 2170 4 n_52
rlabel m2contact 8769 2074 8769 2074 4 n_117
rlabel m2contact 8745 2098 8745 2098 4 n_80
rlabel m2contact 8697 2122 8697 2122 4 n_10
rlabel m2contact 8673 6442 8673 6442 4 n_40
rlabel m2contact 8625 2386 8625 2386 4 n_9
rlabel m2contact 8625 5890 8625 5890 4 n_97
rlabel m2contact 8601 2818 8601 2818 4 OpcodeCondIn[3]
rlabel m2contact 8577 5938 8577 5938 4 n_96
rlabel m2contact 8577 3730 8577 3730 4 OpcodeCondIn[4]
rlabel m2contact 8529 5890 8529 5890 4 n_89
rlabel m2contact 8505 6418 8505 6418 4 n_84
rlabel m2contact 8505 4666 8505 4666 4 n_190
rlabel m2contact 8481 5050 8481 5050 4 n_90
rlabel m2contact 8457 4978 8457 4978 4 n_145
rlabel m2contact 8433 4666 8433 4666 4 n_190
rlabel m2contact 8409 2890 8409 2890 4 n_180
rlabel m2contact 8385 6394 8385 6394 4 n_185
rlabel m2contact 8385 2890 8385 2890 4 n_180
rlabel m2contact 8361 5146 8361 5146 4 n_57
rlabel m2contact 8337 6346 8337 6346 4 n_87
rlabel m2contact 8313 3298 8313 3298 4 n_249
rlabel m2contact 8289 4090 8289 4090 4 n_73
rlabel m2contact 8265 2938 8265 2938 4 n_286
rlabel m2contact 8241 6370 8241 6370 4 n_144
rlabel m2contact 8241 6346 8241 6346 4 n_58
rlabel m2contact 8241 2386 8241 2386 4 n_58
rlabel m2contact 8217 6346 8217 6346 4 n_58
rlabel m2contact 8217 5962 8217 5962 4 n_205
rlabel m2contact 8193 4570 8193 4570 4 n_143
rlabel m2contact 8169 4234 8169 4234 4 n_214
rlabel m2contact 8145 6322 8145 6322 4 n_6
rlabel m2contact 8145 4570 8145 4570 4 n_209
rlabel m2contact 8097 5746 8097 5746 4 OpcodeCondIn[2]
rlabel m2contact 8073 2986 8073 2986 4 n_230
rlabel m2contact 8073 3034 8073 3034 4 OpcodeCondIn[7]
rlabel m2contact 8025 5746 8025 5746 4 OpcodeCondIn[2]
rlabel m2contact 7977 6298 7977 6298 4 n_331
rlabel m2contact 7953 2146 7953 2146 4 Flags[1]
rlabel m2contact 7953 4234 7953 4234 4 n_337
rlabel m2contact 7929 6082 7929 6082 4 n_330
rlabel m2contact 7905 3394 7905 3394 4 n_140
rlabel m2contact 7881 2170 7881 2170 4 n_52
rlabel m2contact 7881 3850 7881 3850 4 stateSub[0]
rlabel m2contact 7857 5170 7857 5170 4 n_210
rlabel m2contact 7857 5146 7857 5146 4 n_57
rlabel m2contact 7809 6274 7809 6274 4 n_240
rlabel m2contact 7785 2194 7785 2194 4 n_319
rlabel m2contact 7785 5242 7785 5242 4 n_200
rlabel m2contact 7761 6250 7761 6250 4 n_109
rlabel m2contact 7713 2218 7713 2218 4 n_266
rlabel m2contact 7713 4402 7713 4402 4 Op1Sel
rlabel m2contact 7665 2458 7665 2458 4 n_221
rlabel m2contact 7665 5554 7665 5554 4 n_264
rlabel m2contact 7641 6226 7641 6226 4 n_296
rlabel m2contact 7641 4738 7641 4738 4 OpcodeCondIn[5]
rlabel m2contact 7617 5578 7617 5578 4 n_220
rlabel m2contact 7593 4402 7593 4402 4 n_297
rlabel m2contact 7569 2242 7569 2242 4 n_129
rlabel m2contact 7569 5842 7569 5842 4 StatusReg[3]
rlabel m2contact 7545 2458 7545 2458 4 n_482
rlabel m2contact 7545 2482 7545 2482 4 n_298
rlabel m2contact 7521 6202 7521 6202 4 n_36
rlabel m2contact 7497 6178 7497 6178 4 n_275
rlabel m2contact 7497 5842 7497 5842 4 n_14
rlabel m2contact 7449 2314 7449 2314 4 n_255
rlabel m2contact 7449 3082 7449 3082 4 n_222
rlabel m2contact 7425 3682 7425 3682 4 n_223
rlabel m2contact 7401 3274 7401 3274 4 n_100
rlabel m2contact 7377 6154 7377 6154 4 n_199
rlabel m2contact 7377 5050 7377 5050 4 n_90
rlabel m2contact 7353 4954 7353 4954 4 n_197
rlabel m2contact 7329 2266 7329 2266 4 n_128
rlabel m2contact 7329 3754 7329 3754 4 n_198
rlabel m2contact 7281 2290 7281 2290 4 n_123
rlabel m2contact 7281 4234 7281 4234 4 n_337
rlabel m2contact 7257 4618 7257 4618 4 n_194
rlabel m2contact 7233 4474 7233 4474 4 n_322
rlabel m2contact 7185 2314 7185 2314 4 n_255
rlabel m2contact 7185 6130 7185 6130 4 n_21
rlabel m2contact 7161 3130 7161 3130 4 state[0]
rlabel m2contact 7137 3994 7137 3994 4 state[1]
rlabel m2contact 7089 2338 7089 2338 4 n_83
rlabel m2contact 7089 2362 7089 2362 4 n_244
rlabel m2contact 7065 3778 7065 3778 4 n_161
rlabel m2contact 7041 2386 7041 2386 4 n_58
rlabel m2contact 7041 3130 7041 3130 4 state[0]
rlabel m2contact 7017 3154 7017 3154 4 n_281
rlabel m2contact 6993 5146 6993 5146 4 n_57
rlabel m2contact 6969 4258 6969 4258 4 n_35
rlabel m2contact 6921 5866 6921 5866 4 OpcodeCondIn[0]
rlabel m2contact 6897 5266 6897 5266 4 n_26
rlabel m2contact 6897 3778 6897 3778 4 n_26
rlabel m2contact 6873 6106 6873 6106 4 n_294
rlabel m2contact 6873 4258 6873 4258 4 n_230
rlabel m2contact 6873 2986 6873 2986 4 n_230
rlabel m2contact 6849 3778 6849 3778 4 n_26
rlabel m2contact 6849 3826 6849 3826 4 nWait
rlabel m2contact 6825 3202 6825 3202 4 n_245
rlabel m2contact 6801 4258 6801 4258 4 n_230
rlabel m2contact 6801 3778 6801 3778 4 n_344
rlabel m2contact 6777 2962 6777 2962 4 n_196
rlabel m2contact 6753 3202 6753 3202 4 n_310
rlabel m2contact 6753 4258 6753 4258 4 n_334
rlabel m2contact 6705 2410 6705 2410 4 n_277
rlabel m2contact 6705 6082 6705 6082 4 n_330
rlabel m2contact 6681 4570 6681 4570 4 n_209
rlabel m2contact 6681 2962 6681 2962 4 n_209
rlabel m2contact 6657 6058 6657 6058 4 n_86
rlabel m2contact 6657 5626 6657 5626 4 n_141
rlabel m2contact 6633 4522 6633 4522 4 n_248
rlabel m2contact 6633 3850 6633 3850 4 stateSub[0]
rlabel m2contact 6609 2962 6609 2962 4 n_209
rlabel m2contact 6609 3250 6609 3250 4 n_92
rlabel m2contact 6561 6034 6561 6034 4 n_193
rlabel m2contact 6561 2962 6561 2962 4 n_72
rlabel m2contact 6537 2434 6537 2434 4 n_7
rlabel m2contact 6537 5554 6537 5554 4 n_264
rlabel m2contact 6513 2890 6513 2890 4 n_180
rlabel m2contact 6513 3754 6513 3754 4 n_198
rlabel m2contact 6489 3538 6489 3538 4 n_192
rlabel m2contact 6465 6010 6465 6010 4 n_211
rlabel m2contact 6441 5986 6441 5986 4 n_207
rlabel m2contact 6441 5242 6441 5242 4 n_200
rlabel m2contact 6417 5770 6417 5770 4 n_176
rlabel m2contact 6417 5170 6417 5170 4 n_210
rlabel m2contact 6393 5962 6393 5962 4 n_205
rlabel m2contact 6369 4138 6369 4138 4 n_254
rlabel m2contact 6345 2458 6345 2458 4 n_482
rlabel m2contact 6321 5866 6321 5866 4 OpcodeCondIn[0]
rlabel m2contact 6321 3946 6321 3946 4 n_258
rlabel m2contact 6297 5914 6297 5914 4 n_53
rlabel m2contact 6297 4762 6297 4762 4 n_79
rlabel m2contact 6273 3130 6273 3130 4 state[0]
rlabel m2contact 6249 2482 6249 2482 4 n_298
rlabel m2contact 6225 4666 6225 4666 4 n_190
rlabel m2contact 6201 5938 6201 5938 4 n_96
rlabel m2contact 6177 5914 6177 5914 4 n_53
rlabel m2contact 6177 4138 6177 4138 4 n_254
rlabel m2contact 6153 5890 6153 5890 4 n_89
rlabel m2contact 6129 5818 6129 5818 4 OpcodeCondIn[1]
rlabel m2contact 6105 2506 6105 2506 4 StatusRegEn
rlabel m2contact 6105 5866 6105 5866 4 OpcodeCondIn[0]
rlabel m2contact 6057 3538 6057 3538 4 n_192
rlabel m2contact 6033 5842 6033 5842 4 n_14
rlabel m2contact 6033 5530 6033 5530 4 n_153
rlabel m2contact 6009 5818 6009 5818 4 OpcodeCondIn[1]
rlabel m2contact 5985 5050 5985 5050 4 n_90
rlabel m2contact 5961 2818 5961 2818 4 OpcodeCondIn[3]
rlabel m2contact 5937 5794 5937 5794 4 n_232
rlabel m2contact 5937 5098 5937 5098 4 n_42
rlabel m2contact 5913 4738 5913 4738 4 OpcodeCondIn[5]
rlabel m2contact 5889 3058 5889 3058 4 n_233
rlabel m2contact 5865 2866 5865 2866 4 n_188
rlabel m2contact 5841 5098 5841 5098 4 n_42
rlabel m2contact 5817 5770 5817 5770 4 n_176
rlabel m2contact 5793 5746 5793 5746 4 OpcodeCondIn[2]
rlabel m2contact 5769 2818 5769 2818 4 OpcodeCondIn[3]
rlabel m2contact 5721 2530 5721 2530 4 n_30
rlabel m2contact 5697 2554 5697 2554 4 StatusReg[2]
rlabel m2contact 5697 2986 5697 2986 4 n_230
rlabel m2contact 5673 5722 5673 5722 4 n_29
rlabel m2contact 5625 5698 5625 5698 4 n_138
rlabel m2contact 5601 3130 5601 3130 4 state[0]
rlabel m2contact 5577 2578 5577 2578 4 n_122
rlabel m2contact 5529 5674 5529 5674 4 n_247
rlabel m2contact 5505 2794 5505 2794 4 n_246
rlabel m2contact 5481 4570 5481 4570 4 n_209
rlabel m2contact 5457 3850 5457 3850 4 stateSub[0]
rlabel m2contact 5409 3730 5409 3730 4 OpcodeCondIn[4]
rlabel m2contact 5361 5650 5361 5650 4 n_177
rlabel m2contact 5313 2842 5313 2842 4 n_142
rlabel m2contact 5289 5626 5289 5626 4 n_141
rlabel m2contact 5289 5602 5289 5602 4 n_357
rlabel m2contact 5241 2602 5241 2602 4 n_265
rlabel m2contact 5217 2890 5217 2890 4 n_180
rlabel m2contact 5193 5578 5193 5578 4 n_220
rlabel m2contact 5169 5554 5169 5554 4 n_264
rlabel m2contact 5145 3946 5145 3946 4 n_258
rlabel m2contact 5121 5530 5121 5530 4 n_153
rlabel m2contact 5121 4186 5121 4186 4 n_131
rlabel m2contact 5073 4618 5073 4618 4 n_194
rlabel m2contact 5049 2626 5049 2626 4 n_339
rlabel m2contact 5049 4570 5049 4570 4 n_209
rlabel m2contact 5001 5506 5001 5506 4 n_33
rlabel m2contact 4953 3274 4953 3274 4 n_100
rlabel m2contact 4953 3850 4953 3850 4 stateSub[0]
rlabel m2contact 4929 5482 4929 5482 4 n_16
rlabel m2contact 4929 3178 4929 3178 4 n_41
rlabel m2contact 4881 5458 4881 5458 4 n_25
rlabel m2contact 4881 5434 4881 5434 4 n_270
rlabel m2contact 4857 2674 4857 2674 4 n_227
rlabel m2contact 4833 2650 4833 2650 4 n_174
rlabel m2contact 4833 3946 4833 3946 4 n_258
rlabel m2contact 4809 5410 4809 5410 4 n_66
rlabel m2contact 4761 4954 4761 4954 4 n_197
rlabel m2contact 4713 2674 4713 2674 4 n_227
rlabel m2contact 4689 5386 4689 5386 4 n_349
rlabel m2contact 4689 2842 4689 2842 4 n_142
rlabel m2contact 4641 5362 4641 5362 4 n_306
rlabel m2contact 4641 5338 4641 5338 4 n_259
rlabel m2contact 4617 3970 4617 3970 4 n_110
rlabel m2contact 4617 3946 4617 3946 4 n_258
rlabel m2contact 4593 2698 4593 2698 4 n_183
rlabel m2contact 4593 2770 4593 2770 4 n_163
rlabel m2contact 4569 3970 4569 3970 4 n_269
rlabel m2contact 4545 2722 4545 2722 4 n_130
rlabel m2contact 4521 5314 4521 5314 4 n_94
rlabel m2contact 4521 2746 4521 2746 4 stateSub[2]
rlabel m2contact 4521 4138 4521 4138 4 n_254
rlabel m2contact 4521 2770 4521 2770 4 n_254
rlabel m2contact 4497 2770 4497 2770 4 n_254
rlabel m2contact 4497 3994 4497 3994 4 state[1]
rlabel m2contact 4473 4090 4473 4090 4 n_73
rlabel m2contact 4449 2794 4449 2794 4 n_246
rlabel m2contact 4425 5290 4425 5290 4 n_282
rlabel m2contact 4401 2818 4401 2818 4 OpcodeCondIn[3]
rlabel m2contact 4377 5266 4377 5266 4 n_26
rlabel m2contact 4377 2842 4377 2842 4 n_142
rlabel m2contact 4353 3682 4353 3682 4 n_223
rlabel m2contact 4305 5242 4305 5242 4 n_200
rlabel m2contact 4305 3154 4305 3154 4 n_281
rlabel m2contact 4281 2866 4281 2866 4 n_188
rlabel m2contact 4281 4666 4281 4666 4 n_190
rlabel m2contact 4257 5218 4257 5218 4 n_126
rlabel m2contact 4209 5194 4209 5194 4 n_156
rlabel m2contact 4209 2890 4209 2890 4 n_180
rlabel m2contact 4185 3538 4185 3538 4 n_192
rlabel m2contact 4161 5170 4161 5170 4 n_210
rlabel m2contact 4161 5122 4161 5122 4 n_65
rlabel m2contact 4113 5146 4113 5146 4 n_57
rlabel m2contact 4113 2914 4113 2914 4 n_70
rlabel m2contact 4113 5122 4113 5122 4 OpcodeCondIn[7]
rlabel m2contact 4113 3034 4113 3034 4 OpcodeCondIn[7]
rlabel m2contact 4089 5122 4089 5122 4 OpcodeCondIn[7]
rlabel m2contact 4089 3850 4089 3850 4 stateSub[0]
rlabel m2contact 4065 5098 4065 5098 4 n_42
rlabel m2contact 4065 4522 4065 4522 4 n_248
rlabel m2contact 4017 2938 4017 2938 4 n_286
rlabel m2contact 4017 5074 4017 5074 4 n_91
rlabel m2contact 3993 2962 3993 2962 4 n_72
rlabel m2contact 3969 5050 3969 5050 4 n_90
rlabel m2contact 3969 2986 3969 2986 4 n_230
rlabel m2contact 3945 3010 3945 3010 4 n_231
rlabel m2contact 3921 5026 3921 5026 4 n_171
rlabel m2contact 3897 5002 3897 5002 4 n_104
rlabel m2contact 3873 4978 3873 4978 4 n_145
rlabel m2contact 3873 3034 3873 3034 4 OpcodeCondIn[7]
rlabel m2contact 3849 3058 3849 3058 4 n_233
rlabel m2contact 3825 3082 3825 3082 4 n_222
rlabel m2contact 3825 4066 3825 4066 4 n_314
rlabel m2contact 3801 4954 3801 4954 4 n_197
rlabel m2contact 3777 3106 3777 3106 4 n_76
rlabel m2contact 3777 4570 3777 4570 4 n_209
rlabel m2contact 3753 4210 3753 4210 4 n_51
rlabel m2contact 3729 3130 3729 3130 4 state[0]
rlabel m2contact 3705 4210 3705 4210 4 n_106
rlabel m2contact 3681 4930 3681 4930 4 n_293
rlabel m2contact 3657 3154 3657 3154 4 n_281
rlabel m2contact 3657 4906 3657 4906 4 n_203
rlabel m2contact 3633 4882 3633 4882 4 n_342
rlabel m2contact 3609 4738 3609 4738 4 OpcodeCondIn[5]
rlabel m2contact 3561 4858 3561 4858 4 n_103
rlabel m2contact 3513 4834 3513 4834 4 n_24
rlabel m2contact 3465 4810 3465 4810 4 n_262
rlabel m2contact 3465 3994 3465 3994 4 state[1]
rlabel m2contact 3441 3538 3441 3538 4 n_192
rlabel m2contact 3417 4786 3417 4786 4 n_112
rlabel m2contact 3417 3178 3417 3178 4 n_41
rlabel m2contact 3393 4762 3393 4762 4 n_79
rlabel m2contact 3345 3202 3345 3202 4 n_310
rlabel m2contact 3321 4738 3321 4738 4 OpcodeCondIn[5]
rlabel m2contact 3297 4714 3297 4714 4 n_309
rlabel m2contact 3225 4690 3225 4690 4 n_201
rlabel m2contact 3177 4666 3177 4666 4 n_190
rlabel m2contact 3129 3226 3129 3226 4 n_195
rlabel m2contact 3105 4642 3105 4642 4 n_162
rlabel m2contact 3081 3754 3081 3754 4 n_198
rlabel m2contact 3057 4618 3057 4618 4 n_194
rlabel m2contact 3057 4594 3057 4594 4 n_291
rlabel m2contact 3009 4570 3009 4570 4 n_209
rlabel m2contact 2961 4546 2961 4546 4 n_111
rlabel m2contact 2937 4522 2937 4522 4 n_248
rlabel m2contact 2937 3250 2937 3250 4 n_92
rlabel m2contact 2889 3274 2889 3274 4 n_100
rlabel m2contact 2889 4498 2889 4498 4 n_323
rlabel m2contact 2865 3298 2865 3298 4 n_249
rlabel m2contact 2865 4474 2865 4474 4 n_322
rlabel m2contact 2841 3322 2841 3322 4 n_175
rlabel m2contact 2817 3346 2817 3346 4 n_113
rlabel m2contact 2793 4450 2793 4450 4 n_365
rlabel m2contact 2769 3370 2769 3370 4 n_284
rlabel m2contact 2745 4426 2745 4426 4 n_328
rlabel m2contact 2721 4402 2721 4402 4 n_297
rlabel m2contact 2697 4378 2697 4378 4 n_149
rlabel m2contact 2673 3394 2673 3394 4 n_140
rlabel m2contact 2673 4354 2673 4354 4 n_85
rlabel m2contact 2649 3418 2649 3418 4 n_121
rlabel m2contact 2649 4330 2649 4330 4 n_22
rlabel m2contact 2625 3442 2625 3442 4 n_68
rlabel m2contact 2601 4306 2601 4306 4 n_358
rlabel m2contact 2553 4282 2553 4282 4 n_208
rlabel m2contact 2553 4258 2553 4258 4 n_334
rlabel m2contact 2529 3466 2529 3466 4 n_302
rlabel m2contact 2529 4234 2529 4234 4 n_337
rlabel m2contact 2481 3706 2481 3706 4 ImmSel
rlabel m2contact 2457 3490 2457 3490 4 n_368
rlabel m2contact 2457 4210 2457 4210 4 n_106
rlabel m2contact 2433 3706 2433 3706 4 n_356
rlabel m2contact 2409 4186 2409 4186 4 n_131
rlabel m2contact 2361 3514 2361 3514 4 n_173
rlabel m2contact 2337 4162 2337 4162 4 n_159
rlabel m2contact 2313 4138 2313 4138 4 n_254
rlabel m2contact 2289 3538 2289 3538 4 n_192
rlabel m2contact 2265 3850 2265 3850 4 stateSub[0]
rlabel m2contact 2241 4114 2241 4114 4 n_69
rlabel m2contact 2241 3946 2241 3946 4 n_258
rlabel m2contact 2241 3538 2241 3538 4 n_258
rlabel m2contact 2217 3538 2217 3538 4 n_258
rlabel m2contact 2217 3850 2217 3850 4 stateSub[0]
rlabel m2contact 2193 4090 2193 4090 4 n_73
rlabel m2contact 2145 3562 2145 3562 4 ENB
rlabel m2contact 2121 4066 2121 4066 4 n_314
rlabel m2contact 2097 4042 2097 4042 4 n_289
rlabel m2contact 2049 4018 2049 4018 4 n_225
rlabel m2contact 2001 3586 2001 3586 4 n_114
rlabel m2contact 1977 3994 1977 3994 4 state[1]
rlabel m2contact 1929 3970 1929 3970 4 n_269
rlabel m2contact 1905 3946 1905 3946 4 n_258
rlabel m2contact 1881 3922 1881 3922 4 n_241
rlabel m2contact 1857 3898 1857 3898 4 n_139
rlabel m2contact 1833 3874 1833 3874 4 n_99
rlabel m2contact 1809 3850 1809 3850 4 stateSub[0]
rlabel m2contact 1785 3610 1785 3610 4 n_64
rlabel m2contact 1737 3634 1737 3634 4 nIRQ
rlabel m2contact 1737 3658 1737 3658 4 ALE
rlabel m2contact 1689 3682 1689 3682 4 n_223
rlabel m2contact 1665 3706 1665 3706 4 n_356
rlabel m2contact 1641 3730 1641 3730 4 OpcodeCondIn[4]
rlabel m2contact 1617 3754 1617 3754 4 n_198
rlabel m2contact 1617 3778 1617 3778 4 n_344
rlabel m2contact 26121 257 26121 257 8 AluOR[1]
rlabel m2contact 26121 41 26121 41 8 AluOR[1]
rlabel m2contact 26097 521 26097 521 8 RegWe
rlabel m2contact 26097 89 26097 89 8 RegWe
rlabel m2contact 26097 65 26097 65 8 AluOR[0]
rlabel m2contact 26097 41 26097 41 8 AluOR[0]
rlabel m2contact 26073 17 26073 17 8 ENB
rlabel metal2 26073 449 26073 449 8 ENB
rlabel m2contact 25521 809 25521 809 6 n_359
rlabel m2contact 25353 713 25353 713 8 n_304
rlabel m2contact 25257 617 25257 617 8 n_60
rlabel m2contact 24657 593 24657 593 8 n_312
rlabel m2contact 24537 665 24537 665 8 n_268
rlabel m2contact 24441 857 24441 857 6 n_170
rlabel m2contact 24345 785 24345 785 8 n_48
rlabel m2contact 24321 137 24321 137 8 n_46
rlabel m2contact 24297 737 24297 737 8 n_47
rlabel m2contact 24129 689 24129 689 8 n_252
rlabel m2contact 24033 89 24033 89 8 n_5
rlabel m2contact 23505 881 23505 881 6 n_224
rlabel m2contact 23481 569 23481 569 8 n_186
rlabel m2contact 23433 497 23433 497 8 n_184
rlabel m2contact 23265 473 23265 473 8 n_136
rlabel m2contact 22905 641 22905 641 8 n_336
rlabel m2contact 22857 545 22857 545 8 n_320
rlabel m2contact 22809 137 22809 137 8 n_46
rlabel m2contact 22785 281 22785 281 8 n_480
rlabel m2contact 22665 449 22665 449 8 n_305
rlabel m2contact 22641 641 22641 641 8 n_336
rlabel m2contact 22521 761 22521 761 8 n_300
rlabel m2contact 22473 641 22473 641 8 n_18
rlabel m2contact 22209 305 22209 305 8 n_169
rlabel m2contact 22137 713 22137 713 8 n_304
rlabel m2contact 22065 689 22065 689 8 n_252
rlabel m2contact 21321 377 21321 377 8 n_132
rlabel m2contact 21297 833 21297 833 6 n_276
rlabel m2contact 21129 713 21129 713 8 n_251
rlabel m2contact 21033 689 21033 689 8 n_292
rlabel m2contact 20961 401 20961 401 8 n_257
rlabel m2contact 20865 353 20865 353 8 n_71
rlabel metal2 20691 425 20691 425 8 SysBus[3]
rlabel m2contact 20673 425 20673 425 8 SysBus[3]
rlabel m2contact 20601 425 20601 425 8 n_267
rlabel m2contact 19641 113 19641 113 8 n_239
rlabel m2contact 19569 161 19569 161 8 n_218
rlabel m2contact 19545 857 19545 857 6 n_170
rlabel m2contact 19521 65 19521 65 8 n_217
rlabel m2contact 19473 209 19473 209 8 n_307
rlabel m2contact 19425 425 19425 425 8 n_267
rlabel m2contact 19401 857 19401 857 6 n_274
rlabel m2contact 19233 593 19233 593 8 n_312
rlabel m2contact 19161 425 19161 425 8 n_256
rlabel m2contact 19089 233 19089 233 8 n_234
rlabel m2contact 19065 305 19065 305 8 n_169
rlabel m2contact 18873 593 18873 593 8 IRQ1
rlabel m2contact 18345 401 18345 401 8 n_257
rlabel m2contact 18225 401 18225 401 8 n_119
rlabel m2contact 18153 881 18153 881 6 n_224
rlabel m2contact 17841 329 17841 329 8 n_45
rlabel m2contact 17649 881 17649 881 6 n_283
rlabel m2contact 17145 185 17145 185 8 n_27
rlabel metal2 17067 17 17067 17 8 SysBus[2]
rlabel m2contact 17049 17 17049 17 8 SysBus[2]
rlabel m2contact 16977 305 16977 305 8 n_169
rlabel m2contact 16905 881 16905 881 6 n_283
rlabel m2contact 16713 785 16713 785 8 n_48
rlabel m2contact 16665 785 16665 785 8 n_335
rlabel m2contact 16593 689 16593 689 8 n_292
rlabel m2contact 16545 689 16545 689 8 n_290
rlabel m2contact 16401 857 16401 857 6 n_274
rlabel m2contact 16353 161 16353 161 8 n_218
rlabel m2contact 16113 161 16113 161 8 IRQ2
rlabel m2contact 15705 593 15705 593 8 IRQ1
rlabel m2contact 15465 593 15465 593 8 n_260
rlabel m2contact 15345 833 15345 833 6 n_276
rlabel m2contact 15129 113 15129 113 8 n_239
rlabel m2contact 14841 497 14841 497 8 n_184
rlabel m2contact 14505 497 14505 497 8 n_44
rlabel m2contact 14385 521 14385 521 8 RegWe
rlabel m2contact 14289 521 14289 521 8 n_167
rlabel m2contact 14145 377 14145 377 8 n_132
rlabel m2contact 14025 113 14025 113 8 n_23
rlabel m2contact 13881 449 13881 449 8 n_305
rlabel m2contact 13785 377 13785 377 8 n_165
rlabel m2contact 13665 449 13665 449 8 n_28
rlabel m2contact 13569 761 13569 761 2 n_300
rlabel m2contact 13353 809 13353 809 4 n_359
rlabel m2contact 13305 785 13305 785 2 n_335
rlabel m2contact 13209 737 13209 737 2 n_47
rlabel m2contact 13113 89 13113 89 2 n_5
rlabel m2contact 13017 89 13017 89 2 nWE
rlabel m2contact 12969 761 12969 761 2 n_300
rlabel m2contact 12849 665 12849 665 2 n_268
rlabel m2contact 12681 665 12681 665 2 n_61
rlabel m2contact 12633 737 12633 737 2 n_47
rlabel m2contact 12609 137 12609 137 2 n_46
rlabel m2contact 12417 257 12417 257 2 AluOR[1]
rlabel m2contact 12369 257 12369 257 2 n_278
rlabel m2contact 12345 593 12345 593 2 n_260
rlabel m2contact 11841 137 11841 137 2 IntStatus
rlabel m2contact 11313 713 11313 713 2 n_251
rlabel m2contact 11265 689 11265 689 2 n_290
rlabel m2contact 11073 665 11073 665 2 n_61
rlabel m2contact 11025 641 11025 641 2 n_18
rlabel m2contact 11001 497 11001 497 2 n_44
rlabel m2contact 10953 65 10953 65 2 n_217
rlabel metal2 10851 497 10851 497 2 SysBus[1]
rlabel m2contact 10833 497 10833 497 2 SysBus[1]
rlabel m2contact 10785 497 10785 497 2 n_98
rlabel m2contact 10713 617 10713 617 2 n_60
rlabel m2contact 10665 521 10665 521 2 n_167
rlabel m2contact 10449 521 10449 521 2 n_101
rlabel m2contact 10305 209 10305 209 2 n_307
rlabel m2contact 10257 257 10257 257 2 n_278
rlabel m2contact 10137 305 10137 305 2 n_169
rlabel m2contact 9873 209 9873 209 2 n_54
rlabel m2contact 9801 41 9801 41 2 AluOR[0]
rlabel m2contact 9753 257 9753 257 2 n_278
rlabel m2contact 9729 593 9729 593 2 n_260
rlabel m2contact 9585 569 9585 569 2 n_186
rlabel m2contact 9345 545 9345 545 2 n_320
rlabel m2contact 9249 521 9249 521 2 n_101
rlabel m2contact 8841 305 8841 305 2 n_169
rlabel m2contact 8721 113 8721 113 2 n_23
rlabel m2contact 8697 329 8697 329 2 n_45
rlabel m2contact 8529 329 8529 329 2 n_191
rlabel m2contact 8481 473 8481 473 2 n_136
rlabel m2contact 8409 353 8409 353 2 n_71
rlabel m2contact 8313 113 8313 113 2 n_288
rlabel m2contact 8289 473 8289 473 2 SysBus[0]
rlabel m2contact 7833 353 7833 353 2 n_20
rlabel m2contact 7737 497 7737 497 2 n_98
rlabel m2contact 7701 473 7701 473 2 SysBus[0]
rlabel m2contact 7305 449 7305 449 2 n_28
rlabel m2contact 7233 425 7233 425 2 n_256
rlabel m2contact 7209 329 7209 329 2 n_191
rlabel m2contact 7137 401 7137 401 2 n_119
rlabel m2contact 7113 329 7113 329 2 n_43
rlabel m2contact 6969 185 6969 185 2 n_27
rlabel m2contact 6897 305 6897 305 2 n_169
rlabel m2contact 6729 185 6729 185 2 n_236
rlabel m2contact 6201 377 6201 377 2 n_165
rlabel m2contact 5985 353 5985 353 2 n_20
rlabel m2contact 5889 329 5889 329 2 n_43
rlabel m2contact 5865 305 5865 305 2 n_169
rlabel m2contact 5649 281 5649 281 2 n_480
rlabel m2contact 5169 257 5169 257 2 n_278
rlabel m2contact 4809 233 4809 233 2 n_234
rlabel m2contact 4329 209 4329 209 2 n_54
rlabel m2contact 3897 185 3897 185 2 n_236
rlabel m2contact 2769 161 2769 161 2 IRQ2
rlabel m2contact 2745 137 2745 137 2 IntStatus
rlabel m2contact 2577 113 2577 113 2 n_288
rlabel m2contact 2409 65 2409 65 2 n_217
rlabel m2contact 1737 65 1737 65 2 nIRQ
rlabel m2contact 25833 7827 25833 7827 6 Flags[2]
rlabel m2contact 25833 7731 25833 7731 6 Flags[2]
rlabel m2contact 25809 7755 25809 7755 6 Flags[3]
rlabel m2contact 25809 7731 25809 7731 6 Flags[3]
rlabel m2contact 25785 7803 25785 7803 6 CFlag
rlabel m2contact 25785 7779 25785 7779 6 CFlag
rlabel m2contact 25785 7755 25785 7755 6 Flags[1]
rlabel m2contact 25785 7707 25785 7707 6 Flags[1]
rlabel m2contact 25761 7779 25761 7779 6 Flags[0]
rlabel m2contact 25761 7683 25761 7683 6 Flags[0]
rlabel m2contact 25737 7755 25737 7755 6 Flags[1]
rlabel metal2 25707 7755 25707 7755 6 StatusRegEn
rlabel m2contact 25689 7755 25689 7755 6 StatusRegEn
rlabel m2contact 24489 7875 24489 7875 6 StatusReg[0]
rlabel m2contact 24417 7851 24417 7851 6 PcWe
rlabel m2contact 24285 7707 24285 7707 6 StatusReg[3]
rlabel m2contact 24009 7827 24009 7827 6 Flags[2]
rlabel m2contact 23481 7827 23481 7827 6 StatusReg[2]
rlabel m2contact 23361 7899 23361 7899 6 Op2Sel[0]
rlabel m2contact 22677 7755 22677 7755 6 StatusReg[1]
rlabel m2contact 22653 7875 22653 7875 6 StatusReg[0]
rlabel m2contact 22161 7827 22161 7827 6 StatusReg[2]
rlabel m2contact 21897 7875 21897 7875 6 WdSel
rlabel m2contact 21069 7923 21069 7923 6 AluEn
rlabel m2contact 20265 7683 20265 7683 6 AluWe
rlabel m2contact 19461 7827 19461 7827 6 Op2Sel[1]
rlabel m2contact 19437 7899 19437 7899 6 Op2Sel[0]
rlabel m2contact 19137 7731 19137 7731 6 Flags[3]
rlabel m2contact 17889 7899 17889 7899 6 PcEn
rlabel m2contact 17853 7731 17853 7731 6 Op1Sel
rlabel m2contact 17829 7899 17829 7899 6 PcEn
rlabel m2contact 17721 7683 17721 7683 6 AluWe
rlabel m2contact 17025 7875 17025 7875 6 WdSel
rlabel m2contact 16857 7803 16857 7803 6 CFlag
rlabel m2contact 16221 7851 16221 7851 6 PcWe
rlabel m2contact 14637 7851 14637 7851 6 PcSel[2]
rlabel m2contact 14337 7875 14337 7875 6 PcSel[0]
rlabel m2contact 14145 7707 14145 7707 6 StatusReg[3]
rlabel m2contact 13833 7899 13833 7899 6 PcSel[1]
rlabel m2contact 13809 7875 13809 7875 6 PcSel[0]
rlabel m2contact 12993 7683 12993 7683 4 MemEn
rlabel m2contact 12657 7755 12657 7755 4 StatusReg[1]
rlabel m2contact 12609 7803 12609 7803 4 CFlag
rlabel m2contact 12213 7947 12213 7947 4 LrEn
rlabel m2contact 12033 7803 12033 7803 4 CFlag
rlabel m2contact 11397 7803 11397 7803 4 LrWe
rlabel m2contact 11169 7755 11169 7755 4 nME
rlabel m2contact 10581 7707 10581 7707 4 LrSel
rlabel metal2 10395 7875 10395 7875 4 ImmSel
rlabel m2contact 10377 7875 10377 7875 4 ImmSel
rlabel m2contact 10065 7875 10065 7875 4 OpcodeCondIn[6]
rlabel metal2 9555 7971 9555 7971 4 IrWe
rlabel m2contact 9537 7971 9537 7971 4 IrWe
rlabel m2contact 9489 7947 9489 7947 4 LrEn
rlabel m2contact 9273 7923 9273 7923 4 AluEn
rlabel m2contact 9153 7899 9153 7899 4 PcSel[1]
rlabel m2contact 8913 7683 8913 7683 4 MemEn
rlabel metal2 8091 7683 8091 7683 4 OpcodeCondIn[7]
rlabel m2contact 8073 7683 8073 7683 4 OpcodeCondIn[7]
rlabel m2contact 8001 7707 8001 7707 4 LrSel
rlabel m2contact 7713 7731 7713 7731 4 Op1Sel
rlabel m2contact 7281 7875 7281 7875 4 OpcodeCondIn[6]
rlabel m2contact 6729 7779 6729 7779 4 Flags[0]
rlabel m2contact 6105 7779 6105 7779 4 OpcodeCondIn[0]
rlabel m2contact 6009 7731 6009 7731 4 OpcodeCondIn[1]
rlabel metal2 5931 7707 5931 7707 4 OpcodeCondIn[5]
rlabel m2contact 5913 7707 5913 7707 4 OpcodeCondIn[5]
rlabel m2contact 5793 7707 5793 7707 4 OpcodeCondIn[2]
rlabel m2contact 5769 7683 5769 7683 4 OpcodeCondIn[3]
rlabel metal2 5427 7875 5427 7875 4 OpcodeCondIn[4]
rlabel m2contact 5409 7875 5409 7875 4 OpcodeCondIn[4]
rlabel m2contact 4833 7683 4833 7683 4 OpcodeCondIn[3]
rlabel m2contact 4737 7851 4737 7851 4 PcSel[2]
rlabel m2contact 4017 7707 4017 7707 4 OpcodeCondIn[2]
rlabel m2contact 3729 7827 3729 7827 4 Op2Sel[1]
rlabel m2contact 3201 7731 3201 7731 4 OpcodeCondIn[1]
rlabel m2contact 2577 7803 2577 7803 4 LrWe
rlabel m2contact 2385 7779 2385 7779 4 OpcodeCondIn[0]
rlabel m2contact 1737 7779 1737 7779 4 ALE
rlabel metal2 25695 7988 25707 7988 6 StatusRegEn
rlabel metal2 24279 7988 24291 7988 6 StatusReg[3]
rlabel metal2 23475 7988 23487 7988 6 StatusReg[2]
rlabel metal2 22671 7988 22683 7988 6 StatusReg[1]
rlabel metal2 22647 7988 22659 7988 6 StatusReg[0]
rlabel metal2 21063 7988 21075 7988 6 AluEn
rlabel metal2 20259 7988 20271 7988 6 AluWe
rlabel metal2 19455 7988 19467 7988 6 Op2Sel[1]
rlabel metal2 19431 7988 19443 7988 6 Op2Sel[0]
rlabel metal2 17847 7988 17859 7988 6 Op1Sel
rlabel metal2 17823 7988 17835 7988 6 PcEn
rlabel metal2 17019 7988 17031 7988 6 WdSel
rlabel metal2 16215 7988 16227 7988 6 PcWe
rlabel metal2 14631 7988 14643 7988 6 PcSel[2]
rlabel metal2 13827 7988 13839 7988 6 PcSel[1]
rlabel metal2 13803 7988 13815 7988 6 PcSel[0]
rlabel metal2 12207 7988 12219 7988 4 LrEn
rlabel metal2 11391 7988 11403 7988 4 LrWe
rlabel metal2 10575 7988 10587 7988 4 LrSel
rlabel metal2 10383 7988 10395 7988 4 ImmSel
rlabel metal2 9543 7988 9555 7988 4 IrWe
rlabel metal2 8907 7988 8919 7988 4 MemEn
rlabel metal2 8079 7988 8091 7988 4 OpcodeCondIn[7]
rlabel metal2 7275 7988 7287 7988 4 OpcodeCondIn[6]
rlabel metal2 5919 7988 5931 7988 4 OpcodeCondIn[5]
rlabel metal2 5415 7988 5427 7988 4 OpcodeCondIn[4]
rlabel metal2 4827 7988 4839 7988 4 OpcodeCondIn[3]
rlabel metal2 4011 7988 4023 7988 4 OpcodeCondIn[2]
rlabel metal2 3195 7988 3207 7988 4 OpcodeCondIn[1]
rlabel metal2 2379 7988 2391 7988 4 OpcodeCondIn[0]
rlabel metal2 20679 0 20691 0 8 SysBus[3]
rlabel metal2 17055 0 17067 0 8 SysBus[2]
rlabel metal2 10839 0 10851 0 2 SysBus[1]
rlabel metal2 7695 0 7707 0 2 SysBus[0]
rlabel metal2 26535 83 26535 95 8 RegWe
rlabel metal2 26535 59 26535 71 8 AluOR[0]
rlabel metal2 26535 35 26535 47 8 AluOR[1]
rlabel metal2 26535 11 26535 23 8 ENB
rlabel metal2 26535 4300 26535 4312 6 Rs1Sel[0]
rlabel metal2 26535 1852 26535 1864 6 Rs1Sel[1]
rlabel metal2 26535 1732 26535 1744 6 RwSel[0]
rlabel metal2 26535 1708 26535 1720 6 RwSel[1]
rlabel metal2 26535 7773 26535 7785 6 CFlag
rlabel metal2 26535 7749 26535 7761 6 Flags[3]
rlabel metal2 26535 7725 26535 7737 6 Flags[2]
rlabel metal2 26535 7701 26535 7713 6 Flags[1]
rlabel metal2 26535 7677 26535 7689 6 Flags[0]
rlabel metal2 26211 7988 26412 7988 5 GND!
rlabel metal2 26211 0 26411 0 1 GND!
rlabel metal2 0 83 0 95 2 nWE
rlabel metal2 0 59 0 71 2 nIRQ
rlabel metal2 0 3820 0 3832 4 nWait
rlabel metal2 0 3796 0 3808 4 nOE
rlabel metal2 0 7773 0 7785 4 ALE
rlabel metal2 0 7749 0 7761 4 nME
rlabel metal2 123 7988 323 7988 5 Vdd!
rlabel metal2 339 7988 351 7988 5 SDO
rlabel metal2 363 7988 375 7988 5 Test
rlabel metal2 387 7988 399 7988 5 Clock
rlabel metal2 411 7988 423 7988 5 nReset
rlabel space 123 0 324 0 1 Vdd!
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 411 0 423 0 1 nReset
<< end >>
