../../../Design/Implementation/verilog/behavioural/io_timer.sv