magic
tech c035u
timestamp 1394494283
<< checkpaint >>
rect 21328 21911 24024 21914
rect -1300 21742 24208 21911
rect -1300 18343 25652 21742
rect -1300 18178 25048 18343
rect -1300 18003 24826 18178
rect -1300 17516 24441 18003
rect -1300 17515 24208 17516
rect -1300 17514 24207 17515
rect -1300 -1300 23897 17514
<< error_s >>
rect 19973 18816 19974 18828
rect 22397 18816 22401 18828
<< metal2 >>
rect 22565 18793 22577 18816
rect 22565 17617 22577 17751
rect 22565 16441 22577 16575
rect 22565 15265 22577 15399
rect 22565 14089 22577 14223
rect 22565 12913 22577 13047
rect 22565 11737 22577 11871
rect 22565 10561 22577 10695
rect 22565 9385 22577 9519
rect 22565 8209 22577 8343
rect 22565 7033 22577 7167
rect 22565 5857 22577 5991
rect 22565 4681 22577 4815
rect 22565 3505 22577 3639
rect 22565 2329 22577 2463
rect 22565 1153 22577 1287
rect 22565 0 22577 111
use slice17  slice17_0
timestamp 1394494283
transform 1 0 4334 0 1 18816
box -4329 0 19127 1795
use leftbuf_slice  leftbuf_slice_0
array 0 0 1469 0 15 1176
timestamp 1394489502
transform 1 0 0 0 1 6
box 0 -6 1469 1170
use IrAA  IrAA_0
array 0 0 1008 0 7 1176
timestamp 1394489502
transform 1 0 1469 0 1 9519
box 0 -111 1008 1065
use LLIcell_U  LLIcell_U_0
array 0 0 6 0 7 1176
timestamp 1393855556
transform 1 0 22517 0 1 9519
box 0 0 192 1042
use IrBA  IrBA_0
array 0 0 1008 0 2 1176
timestamp 1394489502
transform 1 0 1469 0 1 5991
box 0 -111 1008 1065
use IrBB  IrBB_0
array 0 0 1008 0 4 1176
timestamp 1394489502
transform 1 0 1469 0 1 112
box 0 -112 1008 1064
use LLIcell_L  LLIcell_L_0
array 0 0 1 0 7 1176
timestamp 1394447900
transform 1 0 22517 0 1 111
box 0 0 192 1042
use Datapath_slice  Datapath_slice_0
array 0 0 12364 0 15 1176
timestamp 1394491434
transform 1 0 2477 0 1 0
box 0 0 20768 1176
<< labels >>
rlabel metal2 22565 0 22577 0 1 LLI
rlabel metal2 22565 1176 22577 1176 1 LLI
rlabel metal2 22565 2352 22577 2352 1 LLI
rlabel metal2 22565 3528 22577 3528 1 LLI
rlabel metal2 22565 4704 22577 4704 1 LLI
rlabel metal2 22565 5880 22577 5880 1 LLI
rlabel metal2 22565 7056 22577 7056 1 LLI
rlabel metal2 22565 8232 22577 8232 1 LLI
rlabel metal2 22565 10584 22577 10584 1 LLI
rlabel metal2 22565 11760 22577 11760 1 LLI
rlabel metal2 22565 12936 22577 12936 1 LLI
rlabel metal2 22565 14112 22577 14112 1 LLI
rlabel metal2 22565 15288 22577 15288 1 LLI
rlabel metal2 22565 16464 22577 16464 1 LLI
rlabel metal2 22565 17640 22577 17640 1 LLI
rlabel space 22647 18816 22659 18816 1 LLI
<< end >>
