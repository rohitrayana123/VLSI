magic
tech c035u
timestamp 1395696754
<< nwell >>
rect 26115 1443 26427 1841
<< pwell >>
rect 26115 1042 26427 1443
<< pohmic >>
rect 26115 1118 26120 1128
rect 26420 1118 26427 1128
<< nohmic >>
rect 26115 1778 26121 1788
rect 26421 1778 26427 1788
<< psubstratetap >>
rect 26120 1118 26420 1134
<< nsubstratetap >>
rect 26121 1772 26421 1788
<< metal1 >>
rect 13264 7942 23798 7952
rect 10432 7916 10450 7930
rect 11320 7916 11338 7930
rect 12184 7918 22982 7928
rect 9088 7894 15638 7904
rect 20524 7894 20642 7904
rect 21340 7894 21842 7904
rect 3280 7868 3298 7882
rect 5248 7870 7394 7880
rect 8896 7870 12362 7880
rect 12880 7870 14822 7880
rect 17260 7870 17378 7880
rect 17992 7868 18010 7882
rect 19984 7870 26498 7880
rect 2872 7844 2890 7858
rect 3256 7846 4082 7856
rect 5104 7846 6566 7856
rect 6640 7846 11534 7856
rect 12040 7846 18086 7856
rect 19708 7846 23114 7856
rect 84 7822 7322 7832
rect 8632 7822 21350 7832
rect 84 7798 15626 7808
rect 17248 7798 26426 7808
rect 2338 7774 4418 7784
rect 4432 7774 12770 7784
rect 12784 7774 19274 7784
rect 19288 7774 25730 7784
rect 26416 7774 26450 7784
rect 5716 7750 6338 7760
rect 6544 7750 8954 7760
rect 9028 7750 25562 7760
rect 7144 7726 14138 7736
rect 14152 7726 20546 7736
rect 20560 7726 24614 7736
rect 26440 7726 26821 7736
rect 9856 7702 20882 7712
rect 21712 7702 22166 7712
rect 22624 7702 25430 7712
rect 26488 7702 26821 7712
rect 13096 7678 26426 7688
rect 26464 7678 26821 7688
rect 13996 7654 25010 7664
rect 26440 7654 26821 7664
rect 14812 7630 22418 7640
rect 23968 7630 26474 7640
rect 26512 7630 26821 7640
rect 21088 6797 22466 6807
rect 12016 6773 24650 6783
rect 11704 6749 12650 6759
rect 12664 6749 19298 6759
rect 19312 6749 20138 6759
rect 20152 6749 21170 6759
rect 21184 6749 25370 6759
rect 11656 6725 25010 6735
rect 11608 6701 16010 6711
rect 16120 6701 21074 6711
rect 21088 6701 25946 6711
rect 11320 6677 11330 6687
rect 11488 6677 16106 6687
rect 10264 6653 11690 6663
rect 11872 6653 23834 6663
rect 9808 6629 9866 6639
rect 10000 6629 23882 6639
rect 9736 6605 18938 6615
rect 9640 6581 15314 6591
rect 9280 6557 15554 6567
rect 9184 6533 10274 6543
rect 10696 6533 13586 6543
rect 13600 6533 14762 6543
rect 14776 6533 17954 6543
rect 17968 6533 18074 6543
rect 18088 6533 20378 6543
rect 20392 6533 21866 6543
rect 21880 6533 23786 6543
rect 23800 6533 24266 6543
rect 9064 6509 10562 6519
rect 10576 6509 16370 6519
rect 16384 6509 25562 6519
rect 8968 6485 10010 6495
rect 10024 6485 16034 6495
rect 16048 6485 16682 6495
rect 16696 6485 18026 6495
rect 18040 6485 19274 6495
rect 19288 6485 20474 6495
rect 8800 6461 8882 6471
rect 8944 6461 8954 6471
rect 9040 6461 12914 6471
rect 19912 6461 20018 6471
rect 8728 6437 15170 6447
rect 18832 6437 22658 6447
rect 8704 6413 23570 6423
rect 8464 6389 26138 6399
rect 8464 6365 24554 6375
rect 8368 6341 13634 6351
rect 18424 6341 25682 6351
rect 8248 6317 12410 6327
rect 12472 6317 26821 6327
rect 8104 6293 8354 6303
rect 8416 6293 24434 6303
rect 24448 6293 24914 6303
rect 8080 6269 13274 6279
rect 18160 6269 21914 6279
rect 21928 6269 23162 6279
rect 8032 6245 20354 6255
rect 25120 6245 25586 6255
rect 7936 6221 20210 6231
rect 24616 6221 25490 6231
rect 7696 6197 7922 6207
rect 7984 6197 10994 6207
rect 11008 6197 14618 6207
rect 14632 6197 15746 6207
rect 15760 6197 20354 6207
rect 20368 6197 22202 6207
rect 22216 6197 24602 6207
rect 24616 6197 25106 6207
rect 7624 6173 24962 6183
rect 7576 6149 13490 6159
rect 17944 6149 22922 6159
rect 7504 6125 7706 6135
rect 7792 6125 19898 6135
rect 7480 6101 15530 6111
rect 15544 6101 20426 6111
rect 20848 6101 21050 6111
rect 21064 6101 21194 6111
rect 23464 6101 23474 6111
rect 7288 6077 15122 6087
rect 16000 6077 16082 6087
rect 17824 6077 23618 6087
rect 7216 6053 7790 6063
rect 7804 6053 7898 6063
rect 7912 6053 8210 6063
rect 8224 6053 8666 6063
rect 8680 6053 9626 6063
rect 9640 6053 10946 6063
rect 10960 6053 11018 6063
rect 11032 6053 11138 6063
rect 11152 6053 16634 6063
rect 16648 6053 17882 6063
rect 17896 6053 20834 6063
rect 20848 6053 22970 6063
rect 22984 6053 23450 6063
rect 23464 6053 25634 6063
rect 7216 6029 21842 6039
rect 7168 6005 23258 6015
rect 7168 5981 12314 5991
rect 12400 5981 14762 5991
rect 15880 5981 20138 5991
rect 23056 5981 23138 5991
rect 7072 5957 26450 5967
rect 7048 5933 11066 5943
rect 11080 5933 11306 5943
rect 11320 5933 13874 5943
rect 15784 5933 23042 5943
rect 7024 5909 22154 5919
rect 7000 5885 17450 5895
rect 17464 5885 21794 5895
rect 6952 5861 13682 5871
rect 15736 5861 24530 5871
rect 6856 5837 15242 5847
rect 15712 5837 17618 5847
rect 17680 5837 18650 5847
rect 18664 5837 20306 5847
rect 25168 5837 25802 5847
rect 6784 5813 9410 5823
rect 9544 5813 10250 5823
rect 10432 5813 13658 5823
rect 15616 5813 25922 5823
rect 6568 5789 12434 5799
rect 12448 5789 21722 5799
rect 21736 5789 25154 5799
rect 6544 5765 9170 5775
rect 9184 5765 26162 5775
rect 6472 5741 20978 5751
rect 6352 5717 6362 5727
rect 6448 5717 21962 5727
rect 6232 5693 9362 5703
rect 9376 5693 10898 5703
rect 10912 5693 24338 5703
rect 24352 5693 25346 5703
rect 25360 5693 25418 5703
rect 6232 5669 26066 5679
rect 6064 5645 16922 5655
rect 16936 5645 18818 5655
rect 18832 5645 25730 5655
rect 5944 5621 9890 5631
rect 9952 5621 12482 5631
rect 15592 5621 18482 5631
rect 18544 5621 20714 5631
rect 20728 5621 21002 5631
rect 22408 5621 22418 5631
rect 5800 5597 8978 5607
rect 8992 5597 25922 5607
rect 5776 5573 17714 5583
rect 17776 5573 19802 5583
rect 19816 5573 20666 5583
rect 20680 5573 26378 5583
rect 5608 5549 8114 5559
rect 8248 5549 23210 5559
rect 5488 5525 6866 5535
rect 6880 5525 11498 5535
rect 11512 5525 12554 5535
rect 12568 5525 15890 5535
rect 15904 5525 15938 5535
rect 15952 5525 16874 5535
rect 16888 5525 19970 5535
rect 19984 5525 22394 5535
rect 5464 5501 6794 5511
rect 6808 5501 8858 5511
rect 8872 5501 9074 5511
rect 9088 5501 21914 5511
rect 5464 5477 8138 5487
rect 8200 5477 16346 5487
rect 17440 5477 23018 5487
rect 5440 5453 5978 5463
rect 5992 5453 8282 5463
rect 8296 5453 8522 5463
rect 8536 5453 10538 5463
rect 10552 5453 10922 5463
rect 10936 5453 13442 5463
rect 13456 5453 16418 5463
rect 16624 5453 17570 5463
rect 17584 5453 26114 5463
rect 5368 5429 19586 5439
rect 19600 5429 20282 5439
rect 4912 5405 8330 5415
rect 8344 5405 9146 5415
rect 9160 5405 11378 5415
rect 11392 5405 14330 5415
rect 14344 5405 16394 5415
rect 16408 5405 19658 5415
rect 19672 5405 23762 5415
rect 4888 5381 4898 5391
rect 5032 5381 13058 5391
rect 13072 5381 13286 5391
rect 13300 5381 20066 5391
rect 20080 5381 20906 5391
rect 20920 5381 21050 5391
rect 21064 5381 23114 5391
rect 25552 5381 26282 5391
rect 4816 5357 11042 5367
rect 11056 5357 25538 5367
rect 4792 5333 13178 5343
rect 15496 5333 21362 5343
rect 4768 5309 17906 5319
rect 17920 5309 23858 5319
rect 4744 5285 5498 5295
rect 5560 5285 6890 5295
rect 6904 5285 25202 5295
rect 25216 5285 25226 5295
rect 25240 5285 26210 5295
rect 4720 5261 20498 5271
rect 20608 5261 20762 5271
rect 21304 5261 21314 5271
rect 4696 5237 7274 5247
rect 7288 5237 7394 5247
rect 7408 5237 13346 5247
rect 13360 5237 18338 5247
rect 18352 5237 22010 5247
rect 4624 5213 10034 5223
rect 10216 5213 14882 5223
rect 15448 5213 25034 5223
rect 4600 5189 9722 5199
rect 9736 5189 10082 5199
rect 10144 5189 25778 5199
rect 4552 5165 22058 5175
rect 4528 5141 25874 5151
rect 4456 5117 7250 5127
rect 7264 5117 24362 5127
rect 4384 5093 5090 5103
rect 5104 5093 16658 5103
rect 16672 5093 17426 5103
rect 17440 5093 19826 5103
rect 19840 5093 20810 5103
rect 20824 5093 21290 5103
rect 21304 5093 21938 5103
rect 21952 5093 23186 5103
rect 23200 5093 24818 5103
rect 4264 5069 12242 5079
rect 12376 5069 12530 5079
rect 12808 5069 13418 5079
rect 15280 5069 24770 5079
rect 4240 5045 13010 5055
rect 15208 5045 22106 5055
rect 4216 5021 10442 5031
rect 10648 5021 10658 5031
rect 10984 5021 11090 5031
rect 11224 5021 13586 5031
rect 15160 5021 22994 5031
rect 4144 4997 5810 5007
rect 5920 4997 9506 5007
rect 9520 4997 10778 5007
rect 10792 4997 15794 5007
rect 15808 4997 19322 5007
rect 19336 4997 20618 5007
rect 20632 4997 25082 5007
rect 4072 4973 10826 4983
rect 10840 4973 21986 4983
rect 4024 4949 9938 4959
rect 9952 4949 11570 4959
rect 11584 4949 15818 4959
rect 15832 4949 19562 4959
rect 19576 4949 20594 4959
rect 20608 4949 21170 4959
rect 4000 4925 6434 4935
rect 6448 4925 10730 4935
rect 10744 4925 13538 4935
rect 13552 4925 14810 4935
rect 14824 4925 15770 4935
rect 15784 4925 18578 4935
rect 19504 4925 25754 4935
rect 3760 4901 10298 4911
rect 10312 4901 13610 4911
rect 14368 4901 14378 4911
rect 14968 4901 14978 4911
rect 15112 4901 23810 4911
rect 3712 4877 3866 4887
rect 3880 4877 20162 4887
rect 24592 4877 25130 4887
rect 3664 4853 3890 4863
rect 3904 4853 6818 4863
rect 6832 4853 6938 4863
rect 6952 4853 7658 4863
rect 7672 4853 9098 4863
rect 9112 4853 9674 4863
rect 9688 4853 11642 4863
rect 11656 4853 21146 4863
rect 21160 4853 24698 4863
rect 24712 4853 25826 4863
rect 3616 4829 25514 4839
rect 3592 4805 7250 4815
rect 7264 4805 9578 4815
rect 9592 4805 12434 4815
rect 12448 4805 24578 4815
rect 3568 4781 12674 4791
rect 12760 4781 17330 4791
rect 17344 4781 21698 4791
rect 3400 4757 10514 4767
rect 10624 4757 19466 4767
rect 3376 4733 5186 4743
rect 5200 4733 10010 4743
rect 10024 4733 11546 4743
rect 11560 4733 14858 4743
rect 14944 4733 24386 4743
rect 3352 4709 10034 4719
rect 10048 4709 10370 4719
rect 10384 4709 22826 4719
rect 22840 4709 25994 4719
rect 3280 4685 8018 4695
rect 8032 4685 12506 4695
rect 12520 4685 19514 4695
rect 19528 4685 19922 4695
rect 19936 4685 21626 4695
rect 21640 4685 25178 4695
rect 3208 4661 15290 4671
rect 15400 4661 18722 4671
rect 18808 4661 19130 4671
rect 19192 4661 19706 4671
rect 3184 4637 5882 4647
rect 5896 4637 7226 4647
rect 7240 4637 11066 4647
rect 11080 4637 12362 4647
rect 12376 4637 13370 4647
rect 13384 4637 14714 4647
rect 14728 4637 16538 4647
rect 16552 4637 16898 4647
rect 16912 4637 18794 4647
rect 18808 4637 20378 4647
rect 20392 4637 20858 4647
rect 20872 4637 21026 4647
rect 21040 4637 22658 4647
rect 22672 4637 24026 4647
rect 24040 4637 25274 4647
rect 25288 4637 25754 4647
rect 3160 4613 20186 4623
rect 23320 4613 26258 4623
rect 3112 4589 26042 4599
rect 3088 4565 6098 4575
rect 6112 4565 18362 4575
rect 18376 4565 22730 4575
rect 22744 4565 26330 4575
rect 3064 4541 10850 4551
rect 10864 4541 26306 4551
rect 3040 4517 8882 4527
rect 8896 4517 16250 4527
rect 16312 4517 20090 4527
rect 20968 4517 21218 4527
rect 22888 4517 23066 4527
rect 23296 4517 23978 4527
rect 3040 4493 20642 4503
rect 20800 4493 21098 4503
rect 22768 4493 26821 4503
rect 2992 4469 8930 4479
rect 8944 4469 12962 4479
rect 13744 4469 23330 4479
rect 23680 4469 24458 4479
rect 2944 4445 8210 4455
rect 8224 4445 18674 4455
rect 18688 4445 19778 4455
rect 19792 4445 22082 4455
rect 22312 4445 26426 4455
rect 2896 4421 6842 4431
rect 6856 4421 8762 4431
rect 8776 4421 16130 4431
rect 16288 4421 26174 4431
rect 2872 4397 12722 4407
rect 12736 4397 19250 4407
rect 19264 4397 21506 4407
rect 21520 4397 25706 4407
rect 2800 4373 15410 4383
rect 15472 4373 24938 4383
rect 2800 4349 17378 4359
rect 17608 4349 24506 4359
rect 25000 4349 25238 4359
rect 2752 4325 3794 4335
rect 3808 4325 4106 4335
rect 4120 4325 9122 4335
rect 9136 4325 10802 4335
rect 10816 4325 14834 4335
rect 14848 4325 17114 4335
rect 17128 4325 19334 4335
rect 19348 4325 20450 4335
rect 20464 4325 22778 4335
rect 22792 4325 24146 4335
rect 24160 4325 25514 4335
rect 26104 4325 26354 4335
rect 2728 4301 6386 4311
rect 6400 4301 17138 4311
rect 17896 4301 26282 4311
rect 2680 4277 7874 4287
rect 7888 4277 12626 4287
rect 12760 4277 16658 4287
rect 16672 4277 20762 4287
rect 21856 4277 21866 4287
rect 22144 4277 23090 4287
rect 23608 4277 26234 4287
rect 2632 4253 3914 4263
rect 3928 4253 9338 4263
rect 9520 4253 15674 4263
rect 16216 4253 20102 4263
rect 20116 4253 25802 4263
rect 2584 4229 8426 4239
rect 8512 4229 10754 4239
rect 10768 4229 11162 4239
rect 11176 4229 11426 4239
rect 11440 4229 14930 4239
rect 14944 4229 18314 4239
rect 18328 4229 22178 4239
rect 22192 4229 24722 4239
rect 24736 4229 25826 4239
rect 2560 4205 7538 4215
rect 7552 4205 9458 4215
rect 9472 4205 9914 4215
rect 9928 4205 11402 4215
rect 11416 4205 11522 4215
rect 11536 4205 20714 4215
rect 20728 4205 20954 4215
rect 20968 4205 23642 4215
rect 23776 4205 23786 4215
rect 25096 4205 25370 4215
rect 2560 4181 20042 4191
rect 20200 4181 26018 4191
rect 2488 4157 2954 4167
rect 2968 4157 10322 4167
rect 10336 4157 11906 4167
rect 11920 4157 12914 4167
rect 12976 4157 20978 4167
rect 20992 4157 24842 4167
rect 2368 4133 2834 4143
rect 2848 4133 5210 4143
rect 5224 4133 21482 4143
rect 22936 4133 23138 4143
rect 2272 4109 11162 4119
rect 11176 4109 12866 4119
rect 13216 4109 18242 4119
rect 18256 4109 22538 4119
rect 22552 4109 23714 4119
rect 23728 4109 24482 4119
rect 2224 4085 4634 4095
rect 4648 4085 15050 4095
rect 15112 4085 18158 4095
rect 18172 4085 19130 4095
rect 19144 4085 24074 4095
rect 2200 4061 9794 4071
rect 9808 4061 24290 4071
rect 2128 4037 7586 4047
rect 7600 4037 19850 4047
rect 19864 4037 21146 4047
rect 2080 4013 5162 4023
rect 5176 4013 18914 4023
rect 19576 4013 22226 4023
rect 2008 3989 10106 3999
rect 10384 3989 10514 3999
rect 10624 3989 24098 3999
rect 1864 3965 16490 3975
rect 16600 3965 19202 3975
rect 19864 3965 19922 3975
rect 20056 3965 20210 3975
rect 20536 3965 20882 3975
rect 1840 3941 4922 3951
rect 5152 3941 11810 3951
rect 11824 3941 14354 3951
rect 14368 3941 17738 3951
rect 17752 3941 21218 3951
rect 21232 3941 22850 3951
rect 22864 3941 25358 3951
rect 1792 3917 6194 3927
rect 6280 3917 19034 3927
rect 1744 3893 2450 3903
rect 2464 3893 3194 3903
rect 3208 3893 3242 3903
rect 3256 3893 7562 3903
rect 7576 3893 9578 3903
rect 9592 3893 11834 3903
rect 11848 3893 16058 3903
rect 16072 3893 16178 3903
rect 16192 3893 16466 3903
rect 16480 3893 16946 3903
rect 16960 3893 17786 3903
rect 17800 3893 18050 3903
rect 18064 3893 19178 3903
rect 19192 3893 21242 3903
rect 21256 3893 23546 3903
rect 23560 3893 24674 3903
rect 1720 3869 5642 3879
rect 5656 3869 19442 3879
rect 1720 3845 15338 3855
rect 16072 3845 16130 3855
rect 16360 3845 16370 3855
rect 16432 3845 16634 3855
rect 17800 3845 17906 3855
rect 18136 3845 25610 3855
rect 1672 3821 5042 3831
rect 5056 3821 9458 3831
rect 9472 3821 13322 3831
rect 13336 3821 17930 3831
rect 18928 3821 19298 3831
rect 1672 3797 1874 3807
rect 1960 3797 9410 3807
rect 9568 3797 19778 3807
rect 19792 3797 23522 3807
rect 1648 3773 2306 3783
rect 2320 3773 7754 3783
rect 7768 3773 14954 3783
rect 14968 3773 17498 3783
rect 17512 3773 25418 3783
rect 1648 3749 20738 3759
rect 1624 3725 5330 3735
rect 5344 3725 5402 3735
rect 5416 3725 9026 3735
rect 9040 3725 10706 3735
rect 10720 3725 10874 3735
rect 10888 3725 19154 3735
rect 19168 3725 23402 3735
rect 23416 3725 24338 3735
rect 24352 3725 25298 3735
rect 25312 3725 25610 3735
rect 25624 3725 25850 3735
rect 84 3701 7850 3711
rect 7864 3701 22466 3711
rect 25312 3701 25358 3711
rect 84 3677 10154 3687
rect 10696 3677 16274 3687
rect 16288 3677 22274 3687
rect 1624 3653 6410 3663
rect 6424 3653 8402 3663
rect 8416 3653 8570 3663
rect 8584 3653 15962 3663
rect 15976 3653 19634 3663
rect 20752 3653 20906 3663
rect 1768 3629 2642 3639
rect 2656 3629 11450 3639
rect 11464 3629 11618 3639
rect 11632 3629 17690 3639
rect 17704 3629 18698 3639
rect 18712 3629 18986 3639
rect 19000 3629 24722 3639
rect 1792 3605 2426 3615
rect 2440 3605 2762 3615
rect 2776 3605 4346 3615
rect 4360 3605 4970 3615
rect 4984 3605 5234 3615
rect 5248 3605 17762 3615
rect 17776 3605 19754 3615
rect 19768 3605 20258 3615
rect 20272 3605 21602 3615
rect 21616 3605 24818 3615
rect 24832 3605 25322 3615
rect 1840 3581 2522 3591
rect 2536 3581 18890 3591
rect 19168 3581 19334 3591
rect 1912 3557 7634 3567
rect 7696 3557 22706 3567
rect 2368 3533 4202 3543
rect 4216 3533 5306 3543
rect 5320 3533 9050 3543
rect 9064 3533 9386 3543
rect 9400 3533 12386 3543
rect 12400 3533 13154 3543
rect 13168 3533 13778 3543
rect 13792 3533 16802 3543
rect 16816 3533 19370 3543
rect 19384 3533 19610 3543
rect 19624 3533 21266 3543
rect 21280 3533 25442 3543
rect 25456 3533 25898 3543
rect 2536 3509 3386 3519
rect 3400 3509 4874 3519
rect 4888 3509 6338 3519
rect 6352 3509 17042 3519
rect 17056 3509 18098 3519
rect 18112 3509 19322 3519
rect 19336 3509 20162 3519
rect 20176 3509 20234 3519
rect 20248 3509 22802 3519
rect 22816 3509 23426 3519
rect 23440 3509 24866 3519
rect 25456 3509 25946 3519
rect 2608 3485 19730 3495
rect 19744 3485 24194 3495
rect 2632 3461 6314 3471
rect 6328 3461 16322 3471
rect 16336 3461 16706 3471
rect 19744 3461 19802 3471
rect 20248 3461 20282 3471
rect 22720 3461 23018 3471
rect 2680 3437 18866 3447
rect 18880 3437 24986 3447
rect 2728 3413 5690 3423
rect 5704 3413 17210 3423
rect 18880 3413 25130 3423
rect 2752 3389 3290 3399
rect 3304 3389 9818 3399
rect 9832 3389 18842 3399
rect 18856 3389 19610 3399
rect 22816 3389 23114 3399
rect 2968 3365 16154 3375
rect 16168 3365 19682 3375
rect 3016 3341 13394 3351
rect 13408 3341 24626 3351
rect 3088 3317 11738 3327
rect 11752 3317 24506 3327
rect 24520 3317 25394 3327
rect 25408 3317 25850 3327
rect 3112 3293 5090 3303
rect 5104 3293 7994 3303
rect 8008 3293 11042 3303
rect 11056 3293 13466 3303
rect 13480 3293 14210 3303
rect 14224 3293 22034 3303
rect 22048 3293 24242 3303
rect 3184 3269 3674 3279
rect 3688 3269 14402 3279
rect 14416 3269 19082 3279
rect 19096 3269 19418 3279
rect 22048 3269 22610 3279
rect 3232 3245 15050 3255
rect 15064 3245 20690 3255
rect 20704 3245 22274 3255
rect 3304 3221 6242 3231
rect 6256 3221 9602 3231
rect 9616 3221 10490 3231
rect 10504 3221 13034 3231
rect 13048 3221 15026 3231
rect 15040 3221 16562 3231
rect 16576 3221 19706 3231
rect 19720 3221 21122 3231
rect 21136 3221 23402 3231
rect 3448 3197 18002 3207
rect 19096 3197 19586 3207
rect 3472 3173 20306 3183
rect 3520 3149 16562 3159
rect 3952 3125 9818 3135
rect 9832 3125 10466 3135
rect 10480 3125 10970 3135
rect 10984 3125 15002 3135
rect 16168 3125 16250 3135
rect 16528 3125 23474 3135
rect 4096 3101 7106 3111
rect 7120 3101 13226 3111
rect 13240 3101 17306 3111
rect 17320 3101 22562 3111
rect 4120 3077 12122 3087
rect 12136 3077 17234 3087
rect 4168 3053 23690 3063
rect 4288 3029 4754 3039
rect 4816 3029 12842 3039
rect 13168 3029 13286 3039
rect 13336 3029 13418 3039
rect 13480 3029 13658 3039
rect 13720 3029 16826 3039
rect 4312 3005 6002 3015
rect 6016 3005 9770 3015
rect 9784 3005 15986 3015
rect 16000 3005 19538 3015
rect 19552 3005 20786 3015
rect 4336 2981 4514 2991
rect 4528 2981 9866 2991
rect 9880 2981 9914 2991
rect 9928 2981 11090 2991
rect 11104 2981 13130 2991
rect 13144 2981 17834 2991
rect 17848 2981 19394 2991
rect 19408 2981 21962 2991
rect 21976 2981 22442 2991
rect 4360 2957 5858 2967
rect 5872 2957 17234 2967
rect 17248 2957 19658 2967
rect 4432 2933 4898 2943
rect 4912 2933 9482 2943
rect 9496 2933 11546 2943
rect 11560 2933 19058 2943
rect 19072 2933 19226 2943
rect 19240 2933 19514 2943
rect 4864 2909 8138 2919
rect 8152 2909 8954 2919
rect 8968 2909 15842 2919
rect 5248 2885 12026 2895
rect 12280 2885 16226 2895
rect 5272 2861 17402 2871
rect 5296 2837 13106 2847
rect 13120 2837 18962 2847
rect 18976 2837 25634 2847
rect 5320 2813 6362 2823
rect 6376 2813 8090 2823
rect 8104 2813 10394 2823
rect 10408 2813 11930 2823
rect 11944 2813 21890 2823
rect 21904 2813 24170 2823
rect 24184 2813 24890 2823
rect 5344 2789 12530 2799
rect 12784 2789 25058 2799
rect 5584 2765 6002 2775
rect 6064 2765 9842 2775
rect 10072 2765 13178 2775
rect 13192 2765 17546 2775
rect 17560 2765 21098 2775
rect 21112 2765 22898 2775
rect 22912 2765 23498 2775
rect 5824 2741 20570 2751
rect 5872 2717 7442 2727
rect 7456 2717 13250 2727
rect 13360 2717 13490 2727
rect 13864 2717 19010 2727
rect 6112 2693 19106 2703
rect 6160 2669 16778 2679
rect 18976 2669 19466 2679
rect 6328 2645 9218 2655
rect 9232 2645 13898 2655
rect 14128 2645 20930 2655
rect 20944 2645 25970 2655
rect 6376 2621 14906 2631
rect 6496 2597 24794 2607
rect 6592 2573 10850 2583
rect 11224 2573 22418 2583
rect 22432 2573 25238 2583
rect 6640 2549 6650 2559
rect 6712 2549 20474 2559
rect 20488 2549 25466 2559
rect 6688 2525 23714 2535
rect 25480 2525 26174 2535
rect 6736 2501 16322 2511
rect 6928 2477 7058 2487
rect 7120 2477 8546 2487
rect 8560 2477 11594 2487
rect 11608 2477 22250 2487
rect 22264 2477 22682 2487
rect 6976 2453 7370 2463
rect 7384 2453 8306 2463
rect 8320 2453 10586 2463
rect 10600 2453 15002 2463
rect 15016 2453 16442 2463
rect 16456 2453 17858 2463
rect 22696 2453 22970 2463
rect 7000 2429 8426 2439
rect 8440 2429 9698 2439
rect 9712 2429 18266 2439
rect 18280 2429 24746 2439
rect 7192 2405 7418 2415
rect 7432 2405 10226 2415
rect 10240 2405 10634 2415
rect 11248 2405 17474 2415
rect 17872 2405 18158 2415
rect 7336 2381 7394 2391
rect 7480 2381 14090 2391
rect 14152 2381 25490 2391
rect 7384 2357 10658 2367
rect 11296 2357 25658 2367
rect 7528 2333 13754 2343
rect 14488 2333 19994 2343
rect 25672 2333 26378 2343
rect 7600 2309 17618 2319
rect 17632 2309 18218 2319
rect 20008 2309 22346 2319
rect 7768 2285 7790 2295
rect 7840 2285 22946 2295
rect 7816 2261 18434 2271
rect 7912 2237 7922 2247
rect 7984 2237 8810 2247
rect 8824 2237 15914 2247
rect 8008 2213 21650 2223
rect 8320 2189 12818 2199
rect 12832 2189 14042 2199
rect 14056 2189 19394 2199
rect 19408 2189 19946 2199
rect 19960 2189 23930 2199
rect 8344 2165 26402 2175
rect 8536 2141 12074 2151
rect 12568 2141 22514 2151
rect 8584 2117 8618 2127
rect 8680 2117 11330 2127
rect 11416 2117 11642 2127
rect 11968 2117 18050 2127
rect 19960 2117 20102 2127
rect 8752 2093 20018 2103
rect 20032 2093 22370 2103
rect 8848 2069 10754 2079
rect 10768 2069 13514 2079
rect 13528 2069 13562 2079
rect 13576 2069 18770 2079
rect 18784 2069 22490 2079
rect 22504 2069 24050 2079
rect 24064 2069 24890 2079
rect 9232 2045 20402 2055
rect 9280 2021 14378 2031
rect 14536 2021 21314 2031
rect 9496 1997 9626 2007
rect 9760 1997 17978 2007
rect 9616 1973 23378 1983
rect 10144 1949 25586 1959
rect 10504 1925 10562 1935
rect 11368 1925 21194 1935
rect 11656 1901 17522 1911
rect 12856 1877 13082 1887
rect 13456 1877 13634 1887
rect 14728 1877 14978 1887
rect 15928 1877 16010 1887
rect 26464 1877 26821 1887
rect 13528 1853 16082 1863
rect 16096 1853 19874 1863
rect 26440 1853 26821 1863
rect 26115 1824 26427 1834
rect 26115 1801 26427 1811
rect 26115 1772 26121 1788
rect 26421 1772 26427 1788
rect 26115 1763 26427 1772
rect 26115 1134 26427 1143
rect 26115 1118 26120 1134
rect 26420 1118 26427 1134
rect 13264 1020 16730 1030
rect 12880 996 13658 1006
rect 14512 996 25250 1006
rect 12664 972 16082 982
rect 16552 972 20906 982
rect 12616 948 15866 958
rect 15880 948 16706 958
rect 16720 948 21554 958
rect 9904 924 17666 934
rect 7792 900 7802 910
rect 8056 900 13274 910
rect 14464 900 17354 910
rect 7792 876 25226 886
rect 7504 852 12722 862
rect 12736 852 16682 862
rect 7360 828 16826 838
rect 7312 804 9386 814
rect 9688 804 10082 814
rect 12232 804 14186 814
rect 14272 804 15626 814
rect 16480 804 21746 814
rect 7144 780 8498 790
rect 8512 780 10322 790
rect 10336 780 13394 790
rect 14032 780 17162 790
rect 7024 756 9338 766
rect 9664 756 20090 766
rect 20272 756 21674 766
rect 6904 732 10154 742
rect 11344 732 14234 742
rect 14296 732 14594 742
rect 14704 732 16610 742
rect 19024 732 24626 742
rect 6736 708 9122 718
rect 9328 708 9962 718
rect 10216 708 13298 718
rect 13432 708 21410 718
rect 6640 684 17258 694
rect 17464 684 23786 694
rect 6544 660 22226 670
rect 22504 660 23642 670
rect 6280 636 16298 646
rect 16456 636 24290 646
rect 6160 612 22538 622
rect 6136 588 10802 598
rect 10912 588 19058 598
rect 19120 588 23930 598
rect 6088 564 6458 574
rect 6520 564 13802 574
rect 14008 564 22826 574
rect 23608 562 23626 576
rect 26104 564 26138 574
rect 4984 540 16010 550
rect 16384 540 26821 550
rect 4960 516 16970 526
rect 17080 516 23666 526
rect 26056 516 26114 526
rect 4912 492 7802 502
rect 7816 492 17498 502
rect 17512 492 20882 502
rect 20896 492 22754 502
rect 4672 468 22106 478
rect 4648 444 21098 454
rect 4576 420 6746 430
rect 6808 420 26090 430
rect 4552 396 22322 406
rect 22336 396 22418 406
rect 22432 396 24914 406
rect 4480 372 8954 382
rect 9376 372 11474 382
rect 12520 372 24842 382
rect 4456 348 25370 358
rect 4384 324 8762 334
rect 8992 324 17018 334
rect 4192 300 4994 310
rect 6016 300 14018 310
rect 15088 300 15818 310
rect 15832 300 21866 310
rect 4144 276 13634 286
rect 15232 276 18650 286
rect 3544 252 14642 262
rect 3424 228 13970 238
rect 3376 204 10538 214
rect 10552 204 14090 214
rect 14104 204 22874 214
rect 3328 180 9194 190
rect 9712 180 19442 190
rect 3280 156 11114 166
rect 11128 156 20066 166
rect 20080 156 24482 166
rect 3136 132 9242 142
rect 9856 132 14570 142
rect 2992 108 22586 118
rect 2512 84 21314 94
rect 84 60 1706 70
rect 1960 60 6554 70
rect 6616 60 8618 70
rect 8632 60 21194 70
rect 26152 60 26821 70
rect 84 36 2834 46
rect 2896 36 18242 46
rect 26128 36 26821 46
rect 7072 12 7814 22
rect 8272 12 13946 22
rect 26104 12 26821 22
<< m2contact >>
rect 13250 7940 13264 7954
rect 23798 7940 23812 7954
rect 10418 7916 10432 7930
rect 11306 7916 11320 7930
rect 12170 7916 12184 7930
rect 22982 7916 22996 7930
rect 9074 7892 9088 7906
rect 15638 7892 15652 7906
rect 20510 7892 20524 7906
rect 20642 7892 20656 7906
rect 21326 7892 21340 7906
rect 21842 7892 21856 7906
rect 3266 7868 3280 7882
rect 5234 7868 5248 7882
rect 7394 7868 7408 7882
rect 8882 7868 8896 7882
rect 12362 7868 12376 7882
rect 12866 7868 12880 7882
rect 14822 7868 14836 7882
rect 17246 7868 17260 7882
rect 17378 7868 17392 7882
rect 17978 7868 17992 7882
rect 19970 7868 19984 7882
rect 26498 7868 26512 7882
rect 2858 7844 2872 7858
rect 3242 7844 3256 7858
rect 4082 7844 4096 7858
rect 5090 7844 5104 7858
rect 6566 7844 6580 7858
rect 6626 7844 6640 7858
rect 11534 7844 11548 7858
rect 12026 7844 12040 7858
rect 18086 7844 18100 7858
rect 19694 7844 19708 7858
rect 23114 7844 23128 7858
rect 70 7820 84 7834
rect 7322 7820 7336 7834
rect 8618 7820 8632 7834
rect 21350 7820 21364 7834
rect 70 7796 84 7810
rect 15626 7796 15640 7810
rect 17234 7796 17248 7810
rect 26426 7796 26440 7810
rect 2306 7772 2338 7786
rect 4418 7772 4432 7786
rect 12770 7772 12784 7786
rect 19274 7772 19288 7786
rect 25730 7772 25744 7786
rect 26402 7772 26416 7786
rect 26450 7772 26464 7786
rect 5702 7748 5716 7762
rect 6338 7748 6352 7762
rect 6530 7748 6544 7762
rect 8954 7748 8968 7762
rect 9014 7748 9028 7762
rect 25562 7748 25576 7762
rect 7130 7724 7144 7738
rect 14138 7724 14152 7738
rect 20546 7724 20560 7738
rect 24614 7724 24628 7738
rect 26426 7724 26440 7738
rect 26821 7724 26835 7738
rect 9842 7700 9856 7714
rect 20882 7700 20896 7714
rect 21698 7700 21712 7714
rect 22166 7700 22180 7714
rect 22610 7700 22624 7714
rect 25430 7700 25444 7714
rect 26474 7700 26488 7714
rect 26821 7700 26835 7714
rect 13082 7676 13096 7690
rect 26426 7676 26440 7690
rect 26450 7676 26464 7690
rect 26821 7676 26835 7690
rect 13982 7652 13996 7666
rect 25010 7652 25024 7666
rect 26426 7652 26440 7666
rect 26821 7652 26835 7666
rect 14798 7628 14812 7642
rect 22418 7628 22432 7642
rect 23954 7628 23968 7642
rect 26474 7628 26488 7642
rect 26498 7628 26512 7642
rect 26821 7628 26835 7642
rect 21074 6795 21088 6809
rect 22466 6795 22480 6809
rect 12002 6771 12016 6785
rect 24650 6771 24664 6785
rect 11690 6747 11704 6761
rect 12650 6747 12664 6761
rect 19298 6747 19312 6761
rect 20138 6747 20152 6761
rect 21170 6747 21184 6761
rect 25370 6747 25384 6761
rect 11642 6723 11656 6737
rect 25010 6723 25024 6737
rect 11594 6699 11608 6713
rect 16010 6699 16024 6713
rect 16106 6699 16120 6713
rect 21074 6699 21088 6713
rect 25946 6699 25960 6713
rect 11306 6675 11320 6689
rect 11330 6675 11344 6689
rect 11474 6675 11488 6689
rect 16106 6675 16120 6689
rect 10250 6651 10264 6665
rect 11690 6651 11704 6665
rect 11858 6651 11872 6665
rect 23834 6651 23848 6665
rect 9794 6627 9808 6641
rect 9866 6627 9880 6641
rect 9986 6627 10000 6641
rect 23882 6627 23896 6641
rect 9722 6603 9736 6617
rect 18938 6603 18952 6617
rect 9626 6579 9640 6593
rect 15314 6579 15328 6593
rect 9266 6555 9280 6569
rect 15554 6555 15568 6569
rect 9170 6531 9184 6545
rect 10274 6531 10288 6545
rect 10682 6531 10696 6545
rect 13586 6531 13600 6545
rect 14762 6531 14776 6545
rect 17954 6531 17968 6545
rect 18074 6531 18088 6545
rect 20378 6531 20392 6545
rect 21866 6531 21880 6545
rect 23786 6531 23800 6545
rect 24266 6531 24280 6545
rect 9050 6507 9064 6521
rect 10562 6507 10576 6521
rect 16370 6507 16384 6521
rect 25562 6507 25576 6521
rect 8954 6483 8968 6497
rect 10010 6483 10024 6497
rect 16034 6483 16048 6497
rect 16682 6483 16696 6497
rect 18026 6483 18040 6497
rect 19274 6483 19288 6497
rect 20474 6483 20488 6497
rect 8786 6459 8800 6473
rect 8882 6459 8896 6473
rect 8930 6459 8944 6473
rect 8954 6459 8968 6473
rect 9026 6459 9040 6473
rect 12914 6459 12928 6473
rect 19898 6459 19912 6473
rect 20018 6459 20032 6473
rect 8714 6435 8728 6449
rect 15170 6435 15184 6449
rect 18818 6435 18832 6449
rect 22658 6435 22672 6449
rect 8690 6411 8704 6425
rect 23570 6411 23584 6425
rect 8450 6387 8464 6401
rect 26138 6387 26152 6401
rect 8450 6363 8464 6377
rect 24554 6363 24568 6377
rect 8354 6339 8368 6353
rect 13634 6339 13648 6353
rect 18410 6339 18424 6353
rect 25682 6339 25696 6353
rect 8234 6315 8248 6329
rect 12410 6315 12424 6329
rect 12458 6315 12472 6329
rect 26821 6315 26835 6329
rect 8090 6291 8104 6305
rect 8354 6291 8368 6305
rect 8402 6291 8416 6305
rect 24434 6291 24448 6305
rect 24914 6291 24928 6305
rect 8066 6267 8080 6281
rect 13274 6267 13288 6281
rect 18146 6267 18160 6281
rect 21914 6267 21928 6281
rect 23162 6267 23176 6281
rect 8018 6243 8032 6257
rect 20354 6243 20368 6257
rect 25106 6243 25120 6257
rect 25586 6243 25600 6257
rect 7922 6219 7936 6233
rect 20210 6219 20224 6233
rect 24602 6219 24616 6233
rect 25490 6219 25504 6233
rect 7682 6195 7696 6209
rect 7922 6195 7936 6209
rect 7970 6195 7984 6209
rect 10994 6195 11008 6209
rect 14618 6195 14632 6209
rect 15746 6195 15760 6209
rect 20354 6195 20368 6209
rect 22202 6195 22216 6209
rect 24602 6195 24616 6209
rect 25106 6195 25120 6209
rect 7610 6171 7624 6185
rect 24962 6171 24976 6185
rect 7562 6147 7576 6161
rect 13490 6147 13504 6161
rect 17930 6147 17944 6161
rect 22922 6147 22936 6161
rect 7490 6123 7504 6137
rect 7706 6123 7720 6137
rect 7778 6123 7792 6137
rect 19898 6123 19912 6137
rect 7466 6099 7480 6113
rect 15530 6099 15544 6113
rect 20426 6099 20440 6113
rect 20834 6099 20848 6113
rect 21050 6099 21064 6113
rect 21194 6099 21208 6113
rect 23450 6099 23464 6113
rect 23474 6099 23488 6113
rect 7274 6075 7288 6089
rect 15122 6075 15136 6089
rect 15986 6075 16000 6089
rect 16082 6075 16096 6089
rect 17810 6075 17824 6089
rect 23618 6075 23632 6089
rect 7202 6051 7216 6065
rect 7790 6051 7804 6065
rect 7898 6051 7912 6065
rect 8210 6051 8224 6065
rect 8666 6051 8680 6065
rect 9626 6051 9640 6065
rect 10946 6051 10960 6065
rect 11018 6051 11032 6065
rect 11138 6051 11152 6065
rect 16634 6051 16648 6065
rect 17882 6051 17896 6065
rect 20834 6051 20848 6065
rect 22970 6051 22984 6065
rect 23450 6051 23464 6065
rect 25634 6051 25648 6065
rect 7202 6027 7216 6041
rect 21842 6027 21856 6041
rect 7154 6003 7168 6017
rect 23258 6003 23272 6017
rect 7154 5979 7168 5993
rect 12314 5979 12328 5993
rect 12386 5979 12400 5993
rect 14762 5979 14776 5993
rect 15866 5979 15880 5993
rect 20138 5979 20152 5993
rect 23042 5979 23056 5993
rect 23138 5979 23152 5993
rect 7058 5955 7072 5969
rect 26450 5955 26464 5969
rect 7034 5931 7048 5945
rect 11066 5931 11080 5945
rect 11306 5931 11320 5945
rect 13874 5931 13888 5945
rect 15770 5931 15784 5945
rect 23042 5931 23056 5945
rect 7010 5907 7024 5921
rect 22154 5907 22168 5921
rect 6986 5883 7000 5897
rect 17450 5883 17464 5897
rect 21794 5883 21808 5897
rect 6938 5859 6952 5873
rect 13682 5859 13696 5873
rect 15722 5859 15736 5873
rect 24530 5859 24544 5873
rect 6842 5835 6856 5849
rect 15242 5835 15256 5849
rect 15698 5835 15712 5849
rect 17618 5835 17632 5849
rect 17666 5835 17680 5849
rect 18650 5835 18664 5849
rect 20306 5835 20320 5849
rect 25154 5835 25168 5849
rect 25802 5835 25816 5849
rect 6770 5811 6784 5825
rect 9410 5811 9424 5825
rect 9530 5811 9544 5825
rect 10250 5811 10264 5825
rect 10418 5811 10432 5825
rect 13658 5811 13672 5825
rect 15602 5811 15616 5825
rect 25922 5811 25936 5825
rect 6554 5787 6568 5801
rect 12434 5787 12448 5801
rect 21722 5787 21736 5801
rect 25154 5787 25168 5801
rect 6530 5763 6544 5777
rect 9170 5763 9184 5777
rect 26162 5763 26176 5777
rect 6458 5739 6472 5753
rect 20978 5739 20992 5753
rect 6338 5715 6352 5729
rect 6362 5715 6376 5729
rect 6434 5715 6448 5729
rect 21962 5715 21976 5729
rect 6218 5691 6232 5705
rect 9362 5691 9376 5705
rect 10898 5691 10912 5705
rect 24338 5691 24352 5705
rect 25346 5691 25360 5705
rect 25418 5691 25432 5705
rect 6218 5667 6232 5681
rect 26066 5667 26080 5681
rect 6050 5643 6064 5657
rect 16922 5643 16936 5657
rect 18818 5643 18832 5657
rect 25730 5643 25744 5657
rect 5930 5619 5944 5633
rect 9890 5619 9904 5633
rect 9938 5619 9952 5633
rect 12482 5619 12496 5633
rect 15578 5619 15592 5633
rect 18482 5619 18496 5633
rect 18530 5619 18544 5633
rect 20714 5619 20728 5633
rect 21002 5619 21016 5633
rect 22394 5619 22408 5633
rect 22418 5619 22432 5633
rect 5786 5595 5800 5609
rect 8978 5595 8992 5609
rect 25922 5595 25936 5609
rect 5762 5571 5776 5585
rect 17714 5571 17728 5585
rect 17762 5571 17776 5585
rect 19802 5571 19816 5585
rect 20666 5571 20680 5585
rect 26378 5571 26392 5585
rect 5594 5547 5608 5561
rect 8114 5547 8128 5561
rect 8234 5547 8248 5561
rect 23210 5547 23224 5561
rect 5474 5523 5488 5537
rect 6866 5523 6880 5537
rect 11498 5523 11512 5537
rect 12554 5523 12568 5537
rect 15890 5523 15904 5537
rect 15938 5523 15952 5537
rect 16874 5523 16888 5537
rect 19970 5523 19984 5537
rect 22394 5523 22408 5537
rect 5450 5499 5464 5513
rect 6794 5499 6808 5513
rect 8858 5499 8872 5513
rect 9074 5499 9088 5513
rect 21914 5499 21928 5513
rect 5450 5475 5464 5489
rect 8138 5475 8152 5489
rect 8186 5475 8200 5489
rect 16346 5475 16360 5489
rect 17426 5475 17440 5489
rect 23018 5475 23032 5489
rect 5426 5451 5440 5465
rect 5978 5451 5992 5465
rect 8282 5451 8296 5465
rect 8522 5451 8536 5465
rect 10538 5451 10552 5465
rect 10922 5451 10936 5465
rect 13442 5451 13456 5465
rect 16418 5451 16432 5465
rect 16610 5451 16624 5465
rect 17570 5451 17584 5465
rect 26114 5451 26128 5465
rect 5354 5427 5368 5441
rect 19586 5427 19600 5441
rect 20282 5427 20296 5441
rect 4898 5403 4912 5417
rect 8330 5403 8344 5417
rect 9146 5403 9160 5417
rect 11378 5403 11392 5417
rect 14330 5403 14344 5417
rect 16394 5403 16408 5417
rect 19658 5403 19672 5417
rect 23762 5403 23776 5417
rect 4874 5379 4888 5393
rect 4898 5379 4912 5393
rect 5018 5379 5032 5393
rect 13058 5379 13072 5393
rect 13286 5379 13300 5393
rect 20066 5379 20080 5393
rect 20906 5379 20920 5393
rect 21050 5379 21064 5393
rect 23114 5379 23128 5393
rect 25538 5379 25552 5393
rect 26282 5379 26296 5393
rect 4802 5355 4816 5369
rect 11042 5355 11056 5369
rect 25538 5355 25552 5369
rect 4778 5331 4792 5345
rect 13178 5331 13192 5345
rect 15482 5331 15496 5345
rect 21362 5331 21376 5345
rect 4754 5307 4768 5321
rect 17906 5307 17920 5321
rect 23858 5307 23872 5321
rect 4730 5283 4744 5297
rect 5498 5283 5512 5297
rect 5546 5283 5560 5297
rect 6890 5283 6904 5297
rect 25202 5283 25216 5297
rect 25226 5283 25240 5297
rect 26210 5283 26224 5297
rect 4706 5259 4720 5273
rect 20498 5259 20512 5273
rect 20594 5259 20608 5273
rect 20762 5259 20776 5273
rect 21290 5259 21304 5273
rect 21314 5259 21328 5273
rect 4682 5235 4696 5249
rect 7274 5235 7288 5249
rect 7394 5235 7408 5249
rect 13346 5235 13360 5249
rect 18338 5235 18352 5249
rect 22010 5235 22024 5249
rect 4610 5211 4624 5225
rect 10034 5211 10048 5225
rect 10202 5211 10216 5225
rect 14882 5211 14896 5225
rect 15434 5211 15448 5225
rect 25034 5211 25048 5225
rect 4586 5187 4600 5201
rect 9722 5187 9736 5201
rect 10082 5187 10096 5201
rect 10130 5187 10144 5201
rect 25778 5187 25792 5201
rect 4538 5163 4552 5177
rect 22058 5163 22072 5177
rect 4514 5139 4528 5153
rect 25874 5139 25888 5153
rect 4442 5115 4456 5129
rect 7250 5115 7264 5129
rect 24362 5115 24376 5129
rect 4370 5091 4384 5105
rect 5090 5091 5104 5105
rect 16658 5091 16672 5105
rect 17426 5091 17440 5105
rect 19826 5091 19840 5105
rect 20810 5091 20824 5105
rect 21290 5091 21304 5105
rect 21938 5091 21952 5105
rect 23186 5091 23200 5105
rect 24818 5091 24832 5105
rect 4250 5067 4264 5081
rect 12242 5067 12256 5081
rect 12362 5067 12376 5081
rect 12530 5067 12544 5081
rect 12794 5067 12808 5081
rect 13418 5067 13432 5081
rect 15266 5067 15280 5081
rect 24770 5067 24784 5081
rect 4226 5043 4240 5057
rect 13010 5043 13024 5057
rect 15194 5043 15208 5057
rect 22106 5043 22120 5057
rect 4202 5019 4216 5033
rect 10442 5019 10456 5033
rect 10634 5019 10648 5033
rect 10658 5019 10672 5033
rect 10970 5019 10984 5033
rect 11090 5019 11104 5033
rect 11210 5019 11224 5033
rect 13586 5019 13600 5033
rect 15146 5019 15160 5033
rect 22994 5019 23008 5033
rect 4130 4995 4144 5009
rect 5810 4995 5824 5009
rect 5906 4995 5920 5009
rect 9506 4995 9520 5009
rect 10778 4995 10792 5009
rect 15794 4995 15808 5009
rect 19322 4995 19336 5009
rect 20618 4995 20632 5009
rect 25082 4995 25096 5009
rect 4058 4971 4072 4985
rect 10826 4971 10840 4985
rect 21986 4971 22000 4985
rect 4010 4947 4024 4961
rect 9938 4947 9952 4961
rect 11570 4947 11584 4961
rect 15818 4947 15832 4961
rect 19562 4947 19576 4961
rect 20594 4947 20608 4961
rect 21170 4947 21184 4961
rect 3986 4923 4000 4937
rect 6434 4923 6448 4937
rect 10730 4923 10744 4937
rect 13538 4923 13552 4937
rect 14810 4923 14824 4937
rect 15770 4923 15784 4937
rect 18578 4923 18592 4937
rect 19490 4923 19504 4937
rect 25754 4923 25768 4937
rect 3746 4899 3760 4913
rect 10298 4899 10312 4913
rect 13610 4899 13624 4913
rect 14354 4899 14368 4913
rect 14378 4899 14392 4913
rect 14954 4899 14968 4913
rect 14978 4899 14992 4913
rect 15098 4899 15112 4913
rect 23810 4899 23824 4913
rect 3698 4875 3712 4889
rect 3866 4875 3880 4889
rect 20162 4875 20176 4889
rect 24578 4875 24592 4889
rect 25130 4875 25144 4889
rect 3650 4851 3664 4865
rect 3890 4851 3904 4865
rect 6818 4851 6832 4865
rect 6938 4851 6952 4865
rect 7658 4851 7672 4865
rect 9098 4851 9112 4865
rect 9674 4851 9688 4865
rect 11642 4851 11656 4865
rect 21146 4851 21160 4865
rect 24698 4851 24712 4865
rect 25826 4851 25840 4865
rect 3602 4827 3616 4841
rect 25514 4827 25528 4841
rect 3578 4803 3592 4817
rect 7250 4803 7264 4817
rect 9578 4803 9592 4817
rect 12434 4803 12448 4817
rect 24578 4803 24592 4817
rect 3554 4779 3568 4793
rect 12674 4779 12688 4793
rect 12746 4779 12760 4793
rect 17330 4779 17344 4793
rect 21698 4779 21712 4793
rect 3386 4755 3400 4769
rect 10514 4755 10528 4769
rect 10610 4755 10624 4769
rect 19466 4755 19480 4769
rect 3362 4731 3376 4745
rect 5186 4731 5200 4745
rect 10010 4731 10024 4745
rect 11546 4731 11560 4745
rect 14858 4731 14872 4745
rect 14930 4731 14944 4745
rect 24386 4731 24400 4745
rect 3338 4707 3352 4721
rect 10034 4707 10048 4721
rect 10370 4707 10384 4721
rect 22826 4707 22840 4721
rect 25994 4707 26008 4721
rect 3266 4683 3280 4697
rect 8018 4683 8032 4697
rect 12506 4683 12520 4697
rect 19514 4683 19528 4697
rect 19922 4683 19936 4697
rect 21626 4683 21640 4697
rect 25178 4683 25192 4697
rect 3194 4659 3208 4673
rect 15290 4659 15304 4673
rect 15386 4659 15400 4673
rect 18722 4659 18736 4673
rect 18794 4659 18808 4673
rect 19130 4659 19144 4673
rect 19178 4659 19192 4673
rect 19706 4659 19720 4673
rect 3170 4635 3184 4649
rect 5882 4635 5896 4649
rect 7226 4635 7240 4649
rect 11066 4635 11080 4649
rect 12362 4635 12376 4649
rect 13370 4635 13384 4649
rect 14714 4635 14728 4649
rect 16538 4635 16552 4649
rect 16898 4635 16912 4649
rect 18794 4635 18808 4649
rect 20378 4635 20392 4649
rect 20858 4635 20872 4649
rect 21026 4635 21040 4649
rect 22658 4635 22672 4649
rect 24026 4635 24040 4649
rect 25274 4635 25288 4649
rect 25754 4635 25768 4649
rect 3146 4611 3160 4625
rect 20186 4611 20200 4625
rect 23306 4611 23320 4625
rect 26258 4611 26272 4625
rect 3098 4587 3112 4601
rect 26042 4587 26056 4601
rect 3074 4563 3088 4577
rect 6098 4563 6112 4577
rect 18362 4563 18376 4577
rect 22730 4563 22744 4577
rect 26330 4563 26344 4577
rect 3050 4539 3064 4553
rect 10850 4539 10864 4553
rect 26306 4539 26320 4553
rect 3026 4515 3040 4529
rect 8882 4515 8896 4529
rect 16250 4515 16264 4529
rect 16298 4515 16312 4529
rect 20090 4515 20104 4529
rect 20954 4515 20968 4529
rect 21218 4515 21232 4529
rect 22874 4515 22888 4529
rect 23066 4515 23080 4529
rect 23282 4515 23296 4529
rect 23978 4515 23992 4529
rect 3026 4491 3040 4505
rect 20642 4491 20656 4505
rect 20786 4491 20800 4505
rect 21098 4491 21112 4505
rect 22754 4491 22768 4505
rect 26821 4491 26835 4505
rect 2978 4467 2992 4481
rect 8930 4467 8944 4481
rect 12962 4467 12976 4481
rect 13730 4467 13744 4481
rect 23330 4467 23344 4481
rect 23666 4467 23680 4481
rect 24458 4467 24472 4481
rect 2930 4443 2944 4457
rect 8210 4443 8224 4457
rect 18674 4443 18688 4457
rect 19778 4443 19792 4457
rect 22082 4443 22096 4457
rect 22298 4443 22312 4457
rect 26426 4443 26440 4457
rect 2882 4419 2896 4433
rect 6842 4419 6856 4433
rect 8762 4419 8776 4433
rect 16130 4419 16144 4433
rect 16274 4419 16288 4433
rect 26174 4419 26188 4433
rect 2858 4395 2872 4409
rect 12722 4395 12736 4409
rect 19250 4395 19264 4409
rect 21506 4395 21520 4409
rect 25706 4395 25720 4409
rect 2786 4371 2800 4385
rect 15410 4371 15424 4385
rect 15458 4371 15472 4385
rect 24938 4371 24952 4385
rect 2786 4347 2800 4361
rect 17378 4347 17392 4361
rect 17594 4347 17608 4361
rect 24506 4347 24520 4361
rect 24986 4347 25000 4361
rect 25238 4347 25252 4361
rect 2738 4323 2752 4337
rect 3794 4323 3808 4337
rect 4106 4323 4120 4337
rect 9122 4323 9136 4337
rect 10802 4323 10816 4337
rect 14834 4323 14848 4337
rect 17114 4323 17128 4337
rect 19334 4323 19348 4337
rect 20450 4323 20464 4337
rect 22778 4323 22792 4337
rect 24146 4323 24160 4337
rect 25514 4323 25528 4337
rect 26090 4323 26104 4337
rect 26354 4323 26368 4337
rect 2714 4299 2728 4313
rect 6386 4299 6400 4313
rect 17138 4299 17152 4313
rect 17882 4299 17896 4313
rect 26282 4299 26296 4313
rect 2666 4275 2680 4289
rect 7874 4275 7888 4289
rect 12626 4275 12640 4289
rect 12746 4275 12760 4289
rect 16658 4275 16672 4289
rect 20762 4275 20776 4289
rect 21842 4275 21856 4289
rect 21866 4275 21880 4289
rect 22130 4275 22144 4289
rect 23090 4275 23104 4289
rect 23594 4275 23608 4289
rect 26234 4275 26248 4289
rect 2618 4251 2632 4265
rect 3914 4251 3928 4265
rect 9338 4251 9352 4265
rect 9506 4251 9520 4265
rect 15674 4251 15688 4265
rect 16202 4251 16216 4265
rect 20102 4251 20116 4265
rect 25802 4251 25816 4265
rect 2570 4227 2584 4241
rect 8426 4227 8440 4241
rect 8498 4227 8512 4241
rect 10754 4227 10768 4241
rect 11162 4227 11176 4241
rect 11426 4227 11440 4241
rect 14930 4227 14944 4241
rect 18314 4227 18328 4241
rect 22178 4227 22192 4241
rect 24722 4227 24736 4241
rect 25826 4227 25840 4241
rect 2546 4203 2560 4217
rect 7538 4203 7552 4217
rect 9458 4203 9472 4217
rect 9914 4203 9928 4217
rect 11402 4203 11416 4217
rect 11522 4203 11536 4217
rect 20714 4203 20728 4217
rect 20954 4203 20968 4217
rect 23642 4203 23656 4217
rect 23762 4203 23776 4217
rect 23786 4203 23800 4217
rect 25082 4203 25096 4217
rect 25370 4203 25384 4217
rect 2546 4179 2560 4193
rect 20042 4179 20056 4193
rect 20186 4179 20200 4193
rect 26018 4179 26032 4193
rect 2474 4155 2488 4169
rect 2954 4155 2968 4169
rect 10322 4155 10336 4169
rect 11906 4155 11920 4169
rect 12914 4155 12928 4169
rect 12962 4155 12976 4169
rect 20978 4155 20992 4169
rect 24842 4155 24856 4169
rect 2354 4131 2368 4145
rect 2834 4131 2848 4145
rect 5210 4131 5224 4145
rect 21482 4131 21496 4145
rect 22922 4131 22936 4145
rect 23138 4131 23152 4145
rect 2258 4107 2272 4121
rect 11162 4107 11176 4121
rect 12866 4107 12880 4121
rect 13202 4107 13216 4121
rect 18242 4107 18256 4121
rect 22538 4107 22552 4121
rect 23714 4107 23728 4121
rect 24482 4107 24496 4121
rect 2210 4083 2224 4097
rect 4634 4083 4648 4097
rect 15050 4083 15064 4097
rect 15098 4083 15112 4097
rect 18158 4083 18172 4097
rect 19130 4083 19144 4097
rect 24074 4083 24088 4097
rect 2186 4059 2200 4073
rect 9794 4059 9808 4073
rect 24290 4059 24304 4073
rect 2114 4035 2128 4049
rect 7586 4035 7600 4049
rect 19850 4035 19864 4049
rect 21146 4035 21160 4049
rect 2066 4011 2080 4025
rect 5162 4011 5176 4025
rect 18914 4011 18928 4025
rect 19562 4011 19576 4025
rect 22226 4011 22240 4025
rect 1994 3987 2008 4001
rect 10106 3987 10120 4001
rect 10370 3987 10384 4001
rect 10514 3987 10528 4001
rect 10610 3987 10624 4001
rect 24098 3987 24112 4001
rect 1850 3963 1864 3977
rect 16490 3963 16504 3977
rect 16586 3963 16600 3977
rect 19202 3963 19216 3977
rect 19850 3963 19864 3977
rect 19922 3963 19936 3977
rect 20042 3963 20056 3977
rect 20210 3963 20224 3977
rect 20522 3963 20536 3977
rect 20882 3963 20896 3977
rect 1826 3939 1840 3953
rect 4922 3939 4936 3953
rect 5138 3939 5152 3953
rect 11810 3939 11824 3953
rect 14354 3939 14368 3953
rect 17738 3939 17752 3953
rect 21218 3939 21232 3953
rect 22850 3939 22864 3953
rect 25358 3939 25372 3953
rect 1778 3915 1792 3929
rect 6194 3915 6208 3929
rect 6266 3915 6280 3929
rect 19034 3915 19048 3929
rect 1730 3891 1744 3905
rect 2450 3891 2464 3905
rect 3194 3891 3208 3905
rect 3242 3891 3256 3905
rect 7562 3891 7576 3905
rect 9578 3891 9592 3905
rect 11834 3891 11848 3905
rect 16058 3891 16072 3905
rect 16178 3891 16192 3905
rect 16466 3891 16480 3905
rect 16946 3891 16960 3905
rect 17786 3891 17800 3905
rect 18050 3891 18064 3905
rect 19178 3891 19192 3905
rect 21242 3891 21256 3905
rect 23546 3891 23560 3905
rect 24674 3891 24688 3905
rect 1706 3867 1720 3881
rect 5642 3867 5656 3881
rect 19442 3867 19456 3881
rect 1706 3843 1720 3857
rect 15338 3843 15352 3857
rect 16058 3843 16072 3857
rect 16130 3843 16144 3857
rect 16346 3843 16360 3857
rect 16370 3843 16384 3857
rect 16418 3843 16432 3857
rect 16634 3843 16648 3857
rect 17786 3843 17800 3857
rect 17906 3843 17920 3857
rect 18122 3843 18136 3857
rect 25610 3843 25624 3857
rect 1658 3819 1672 3833
rect 5042 3819 5056 3833
rect 9458 3819 9472 3833
rect 13322 3819 13336 3833
rect 17930 3819 17944 3833
rect 18914 3819 18928 3833
rect 19298 3819 19312 3833
rect 1658 3795 1672 3809
rect 1874 3795 1888 3809
rect 1946 3795 1960 3809
rect 9410 3795 9424 3809
rect 9554 3795 9568 3809
rect 19778 3795 19792 3809
rect 23522 3795 23536 3809
rect 1634 3771 1648 3785
rect 2306 3771 2320 3785
rect 7754 3771 7768 3785
rect 14954 3771 14968 3785
rect 17498 3771 17512 3785
rect 25418 3771 25432 3785
rect 1634 3747 1648 3761
rect 20738 3747 20752 3761
rect 1610 3723 1624 3737
rect 5330 3723 5344 3737
rect 5402 3723 5416 3737
rect 9026 3723 9040 3737
rect 10706 3723 10720 3737
rect 10874 3723 10888 3737
rect 19154 3723 19168 3737
rect 23402 3723 23416 3737
rect 24338 3723 24352 3737
rect 25298 3723 25312 3737
rect 25610 3723 25624 3737
rect 25850 3723 25864 3737
rect 70 3699 84 3713
rect 7850 3699 7864 3713
rect 22466 3699 22480 3713
rect 25298 3699 25312 3713
rect 25358 3699 25372 3713
rect 70 3675 84 3689
rect 10154 3675 10168 3689
rect 10682 3675 10696 3689
rect 16274 3675 16288 3689
rect 22274 3675 22288 3689
rect 1610 3651 1624 3665
rect 6410 3651 6424 3665
rect 8402 3651 8416 3665
rect 8570 3651 8584 3665
rect 15962 3651 15976 3665
rect 19634 3651 19648 3665
rect 20738 3651 20752 3665
rect 20906 3651 20920 3665
rect 1754 3627 1768 3641
rect 2642 3627 2656 3641
rect 11450 3627 11464 3641
rect 11618 3627 11632 3641
rect 17690 3627 17704 3641
rect 18698 3627 18712 3641
rect 18986 3627 19000 3641
rect 24722 3627 24736 3641
rect 1778 3603 1792 3617
rect 2426 3603 2440 3617
rect 2762 3603 2776 3617
rect 4346 3603 4360 3617
rect 4970 3603 4984 3617
rect 5234 3603 5248 3617
rect 17762 3603 17776 3617
rect 19754 3603 19768 3617
rect 20258 3603 20272 3617
rect 21602 3603 21616 3617
rect 24818 3603 24832 3617
rect 25322 3603 25336 3617
rect 1826 3579 1840 3593
rect 2522 3579 2536 3593
rect 18890 3579 18904 3593
rect 19154 3579 19168 3593
rect 19334 3579 19348 3593
rect 1898 3555 1912 3569
rect 7634 3555 7648 3569
rect 7682 3555 7696 3569
rect 22706 3555 22720 3569
rect 2354 3531 2368 3545
rect 4202 3531 4216 3545
rect 5306 3531 5320 3545
rect 9050 3531 9064 3545
rect 9386 3531 9400 3545
rect 12386 3531 12400 3545
rect 13154 3531 13168 3545
rect 13778 3531 13792 3545
rect 16802 3531 16816 3545
rect 19370 3531 19384 3545
rect 19610 3531 19624 3545
rect 21266 3531 21280 3545
rect 25442 3531 25456 3545
rect 25898 3531 25912 3545
rect 2522 3507 2536 3521
rect 3386 3507 3400 3521
rect 4874 3507 4888 3521
rect 6338 3507 6352 3521
rect 17042 3507 17056 3521
rect 18098 3507 18112 3521
rect 19322 3507 19336 3521
rect 20162 3507 20176 3521
rect 20234 3507 20248 3521
rect 22802 3507 22816 3521
rect 23426 3507 23440 3521
rect 24866 3507 24880 3521
rect 25442 3507 25456 3521
rect 25946 3507 25960 3521
rect 2594 3483 2608 3497
rect 19730 3483 19744 3497
rect 24194 3483 24208 3497
rect 2618 3459 2632 3473
rect 6314 3459 6328 3473
rect 16322 3459 16336 3473
rect 16706 3459 16720 3473
rect 19730 3459 19744 3473
rect 19802 3459 19816 3473
rect 20234 3459 20248 3473
rect 20282 3459 20296 3473
rect 22706 3459 22720 3473
rect 23018 3459 23032 3473
rect 2666 3435 2680 3449
rect 18866 3435 18880 3449
rect 24986 3435 25000 3449
rect 2714 3411 2728 3425
rect 5690 3411 5704 3425
rect 17210 3411 17224 3425
rect 18866 3411 18880 3425
rect 25130 3411 25144 3425
rect 2738 3387 2752 3401
rect 3290 3387 3304 3401
rect 9818 3387 9832 3401
rect 18842 3387 18856 3401
rect 19610 3387 19624 3401
rect 22802 3387 22816 3401
rect 23114 3387 23128 3401
rect 2954 3363 2968 3377
rect 16154 3363 16168 3377
rect 19682 3363 19696 3377
rect 3002 3339 3016 3353
rect 13394 3339 13408 3353
rect 24626 3339 24640 3353
rect 3074 3315 3088 3329
rect 11738 3315 11752 3329
rect 24506 3315 24520 3329
rect 25394 3315 25408 3329
rect 25850 3315 25864 3329
rect 3098 3291 3112 3305
rect 5090 3291 5104 3305
rect 7994 3291 8008 3305
rect 11042 3291 11056 3305
rect 13466 3291 13480 3305
rect 14210 3291 14224 3305
rect 22034 3291 22048 3305
rect 24242 3291 24256 3305
rect 3170 3267 3184 3281
rect 3674 3267 3688 3281
rect 14402 3267 14416 3281
rect 19082 3267 19096 3281
rect 19418 3267 19432 3281
rect 22034 3267 22048 3281
rect 22610 3267 22624 3281
rect 3218 3243 3232 3257
rect 15050 3243 15064 3257
rect 20690 3243 20704 3257
rect 22274 3243 22288 3257
rect 3290 3219 3304 3233
rect 6242 3219 6256 3233
rect 9602 3219 9616 3233
rect 10490 3219 10504 3233
rect 13034 3219 13048 3233
rect 15026 3219 15040 3233
rect 16562 3219 16576 3233
rect 19706 3219 19720 3233
rect 21122 3219 21136 3233
rect 23402 3219 23416 3233
rect 3434 3195 3448 3209
rect 18002 3195 18016 3209
rect 19082 3195 19096 3209
rect 19586 3195 19600 3209
rect 3458 3171 3472 3185
rect 20306 3171 20320 3185
rect 3506 3147 3520 3161
rect 16562 3147 16576 3161
rect 3938 3123 3952 3137
rect 9818 3123 9832 3137
rect 10466 3123 10480 3137
rect 10970 3123 10984 3137
rect 15002 3123 15016 3137
rect 16154 3123 16168 3137
rect 16250 3123 16264 3137
rect 16514 3123 16528 3137
rect 23474 3123 23488 3137
rect 4082 3099 4096 3113
rect 7106 3099 7120 3113
rect 13226 3099 13240 3113
rect 17306 3099 17320 3113
rect 22562 3099 22576 3113
rect 4106 3075 4120 3089
rect 12122 3075 12136 3089
rect 17234 3075 17248 3089
rect 4154 3051 4168 3065
rect 23690 3051 23704 3065
rect 4274 3027 4288 3041
rect 4754 3027 4768 3041
rect 4802 3027 4816 3041
rect 12842 3027 12856 3041
rect 13154 3027 13168 3041
rect 13286 3027 13300 3041
rect 13322 3027 13336 3041
rect 13418 3027 13432 3041
rect 13466 3027 13480 3041
rect 13658 3027 13672 3041
rect 13706 3027 13720 3041
rect 16826 3027 16840 3041
rect 4298 3003 4312 3017
rect 6002 3003 6016 3017
rect 9770 3003 9784 3017
rect 15986 3003 16000 3017
rect 19538 3003 19552 3017
rect 20786 3003 20800 3017
rect 4322 2979 4336 2993
rect 4514 2979 4528 2993
rect 9866 2979 9880 2993
rect 9914 2979 9928 2993
rect 11090 2979 11104 2993
rect 13130 2979 13144 2993
rect 17834 2979 17848 2993
rect 19394 2979 19408 2993
rect 21962 2979 21976 2993
rect 22442 2979 22456 2993
rect 4346 2955 4360 2969
rect 5858 2955 5872 2969
rect 17234 2955 17248 2969
rect 19658 2955 19672 2969
rect 4418 2931 4432 2945
rect 4898 2931 4912 2945
rect 9482 2931 9496 2945
rect 11546 2931 11560 2945
rect 19058 2931 19072 2945
rect 19226 2931 19240 2945
rect 19514 2931 19528 2945
rect 4850 2907 4864 2921
rect 8138 2907 8152 2921
rect 8954 2907 8968 2921
rect 15842 2907 15856 2921
rect 5234 2883 5248 2897
rect 12026 2883 12040 2897
rect 12266 2883 12280 2897
rect 16226 2883 16240 2897
rect 5258 2859 5272 2873
rect 17402 2859 17416 2873
rect 5282 2835 5296 2849
rect 13106 2835 13120 2849
rect 18962 2835 18976 2849
rect 25634 2835 25648 2849
rect 5306 2811 5320 2825
rect 6362 2811 6376 2825
rect 8090 2811 8104 2825
rect 10394 2811 10408 2825
rect 11930 2811 11944 2825
rect 21890 2811 21904 2825
rect 24170 2811 24184 2825
rect 24890 2811 24904 2825
rect 5330 2787 5344 2801
rect 12530 2787 12544 2801
rect 12770 2787 12784 2801
rect 25058 2787 25072 2801
rect 5570 2763 5584 2777
rect 6002 2763 6016 2777
rect 6050 2763 6064 2777
rect 9842 2763 9856 2777
rect 10058 2763 10072 2777
rect 13178 2763 13192 2777
rect 17546 2763 17560 2777
rect 21098 2763 21112 2777
rect 22898 2763 22912 2777
rect 23498 2763 23512 2777
rect 5810 2739 5824 2753
rect 20570 2739 20584 2753
rect 5858 2715 5872 2729
rect 7442 2715 7456 2729
rect 13250 2715 13264 2729
rect 13346 2715 13360 2729
rect 13490 2715 13504 2729
rect 13850 2715 13864 2729
rect 19010 2715 19024 2729
rect 6098 2691 6112 2705
rect 19106 2691 19120 2705
rect 6146 2667 6160 2681
rect 16778 2667 16792 2681
rect 18962 2667 18976 2681
rect 19466 2667 19480 2681
rect 6314 2643 6328 2657
rect 9218 2643 9232 2657
rect 13898 2643 13912 2657
rect 14114 2643 14128 2657
rect 20930 2643 20944 2657
rect 25970 2643 25984 2657
rect 6362 2619 6376 2633
rect 14906 2619 14920 2633
rect 6482 2595 6496 2609
rect 24794 2595 24808 2609
rect 6578 2571 6592 2585
rect 10850 2571 10864 2585
rect 11210 2571 11224 2585
rect 22418 2571 22432 2585
rect 25238 2571 25252 2585
rect 6626 2547 6640 2561
rect 6650 2547 6664 2561
rect 6698 2547 6712 2561
rect 20474 2547 20488 2561
rect 25466 2547 25480 2561
rect 6674 2523 6688 2537
rect 23714 2523 23728 2537
rect 25466 2523 25480 2537
rect 26174 2523 26188 2537
rect 6722 2499 6736 2513
rect 16322 2499 16336 2513
rect 6914 2475 6928 2489
rect 7058 2475 7072 2489
rect 7106 2475 7120 2489
rect 8546 2475 8560 2489
rect 11594 2475 11608 2489
rect 22250 2475 22264 2489
rect 22682 2475 22696 2489
rect 6962 2451 6976 2465
rect 7370 2451 7384 2465
rect 8306 2451 8320 2465
rect 10586 2451 10600 2465
rect 15002 2451 15016 2465
rect 16442 2451 16456 2465
rect 17858 2451 17872 2465
rect 22682 2451 22696 2465
rect 22970 2451 22984 2465
rect 6986 2427 7000 2441
rect 8426 2427 8440 2441
rect 9698 2427 9712 2441
rect 18266 2427 18280 2441
rect 24746 2427 24760 2441
rect 7178 2403 7192 2417
rect 7418 2403 7432 2417
rect 10226 2403 10240 2417
rect 10634 2403 10648 2417
rect 11234 2403 11248 2417
rect 17474 2403 17488 2417
rect 17858 2403 17872 2417
rect 18158 2403 18172 2417
rect 7322 2379 7336 2393
rect 7394 2379 7408 2393
rect 7466 2379 7480 2393
rect 14090 2379 14104 2393
rect 14138 2379 14152 2393
rect 25490 2379 25504 2393
rect 7370 2355 7384 2369
rect 10658 2355 10672 2369
rect 11282 2355 11296 2369
rect 25658 2355 25672 2369
rect 7514 2331 7528 2345
rect 13754 2331 13768 2345
rect 14474 2331 14488 2345
rect 19994 2331 20008 2345
rect 25658 2331 25672 2345
rect 26378 2331 26392 2345
rect 7586 2307 7600 2321
rect 17618 2307 17632 2321
rect 18218 2307 18232 2321
rect 19994 2307 20008 2321
rect 22346 2307 22360 2321
rect 7754 2283 7768 2297
rect 7790 2283 7804 2297
rect 7826 2283 7840 2297
rect 22946 2283 22960 2297
rect 7802 2259 7816 2273
rect 18434 2259 18448 2273
rect 7898 2235 7912 2249
rect 7922 2235 7936 2249
rect 7970 2235 7984 2249
rect 8810 2235 8824 2249
rect 15914 2235 15928 2249
rect 7994 2211 8008 2225
rect 21650 2211 21664 2225
rect 8306 2187 8320 2201
rect 12818 2187 12832 2201
rect 14042 2187 14056 2201
rect 19394 2187 19408 2201
rect 19946 2187 19960 2201
rect 23930 2187 23944 2201
rect 8330 2163 8344 2177
rect 26402 2163 26416 2177
rect 8522 2139 8536 2153
rect 12074 2139 12088 2153
rect 12554 2139 12568 2153
rect 22514 2139 22528 2153
rect 8570 2115 8584 2129
rect 8618 2115 8632 2129
rect 8666 2115 8680 2129
rect 11330 2115 11344 2129
rect 11402 2115 11416 2129
rect 11642 2115 11656 2129
rect 11954 2115 11968 2129
rect 18050 2115 18064 2129
rect 19946 2115 19960 2129
rect 20102 2115 20116 2129
rect 8738 2091 8752 2105
rect 20018 2091 20032 2105
rect 22370 2091 22384 2105
rect 8834 2067 8848 2081
rect 10754 2067 10768 2081
rect 13514 2067 13528 2081
rect 13562 2067 13576 2081
rect 18770 2067 18784 2081
rect 22490 2067 22504 2081
rect 24050 2067 24064 2081
rect 24890 2067 24904 2081
rect 9218 2043 9232 2057
rect 20402 2043 20416 2057
rect 9266 2019 9280 2033
rect 14378 2019 14392 2033
rect 14522 2019 14536 2033
rect 21314 2019 21328 2033
rect 9482 1995 9496 2009
rect 9626 1995 9640 2009
rect 9746 1995 9760 2009
rect 17978 1995 17992 2009
rect 9602 1971 9616 1985
rect 23378 1971 23392 1985
rect 10130 1947 10144 1961
rect 25586 1947 25600 1961
rect 10490 1923 10504 1937
rect 10562 1923 10576 1937
rect 11354 1923 11368 1937
rect 21194 1923 21208 1937
rect 11642 1899 11656 1913
rect 17522 1899 17536 1913
rect 12842 1875 12856 1889
rect 13082 1875 13096 1889
rect 13442 1875 13456 1889
rect 13634 1875 13648 1889
rect 14714 1875 14728 1889
rect 14978 1875 14992 1889
rect 15914 1875 15928 1889
rect 16010 1875 16024 1889
rect 26450 1875 26464 1889
rect 26821 1875 26835 1889
rect 13514 1851 13528 1865
rect 16082 1851 16096 1865
rect 19874 1851 19888 1865
rect 26426 1851 26440 1865
rect 26821 1851 26835 1865
rect 13250 1018 13264 1032
rect 16730 1018 16744 1032
rect 12866 994 12880 1008
rect 13658 994 13672 1008
rect 14498 994 14512 1008
rect 25250 994 25264 1008
rect 12650 970 12664 984
rect 16082 970 16096 984
rect 16538 970 16552 984
rect 20906 970 20920 984
rect 12602 946 12616 960
rect 15866 946 15880 960
rect 16706 946 16720 960
rect 21554 946 21568 960
rect 9890 922 9904 936
rect 17666 922 17680 936
rect 7778 898 7792 912
rect 7802 898 7816 912
rect 8042 898 8056 912
rect 13274 898 13288 912
rect 14450 898 14464 912
rect 17354 898 17368 912
rect 7778 874 7792 888
rect 25226 874 25240 888
rect 7490 850 7504 864
rect 12722 850 12736 864
rect 16682 850 16696 864
rect 7346 826 7360 840
rect 16826 826 16840 840
rect 7298 802 7312 816
rect 9386 802 9400 816
rect 9674 802 9688 816
rect 10082 802 10096 816
rect 12218 802 12232 816
rect 14186 802 14200 816
rect 14258 802 14272 816
rect 15626 802 15640 816
rect 16466 802 16480 816
rect 21746 802 21760 816
rect 7130 778 7144 792
rect 8498 778 8512 792
rect 10322 778 10336 792
rect 13394 778 13408 792
rect 14018 778 14032 792
rect 17162 778 17176 792
rect 7010 754 7024 768
rect 9338 754 9352 768
rect 9650 754 9664 768
rect 20090 754 20104 768
rect 20258 754 20272 768
rect 21674 754 21688 768
rect 6890 730 6904 744
rect 10154 730 10168 744
rect 11330 730 11344 744
rect 14234 730 14248 744
rect 14282 730 14296 744
rect 14594 730 14608 744
rect 14690 730 14704 744
rect 16610 730 16624 744
rect 19010 730 19024 744
rect 24626 730 24640 744
rect 6722 706 6736 720
rect 9122 706 9136 720
rect 9314 706 9328 720
rect 9962 706 9976 720
rect 10202 706 10216 720
rect 13298 706 13312 720
rect 13418 706 13432 720
rect 21410 706 21424 720
rect 6626 682 6640 696
rect 17258 682 17272 696
rect 17450 682 17464 696
rect 23786 682 23800 696
rect 6530 658 6544 672
rect 22226 658 22240 672
rect 22490 658 22504 672
rect 23642 658 23656 672
rect 6266 634 6280 648
rect 16298 634 16312 648
rect 16442 634 16456 648
rect 24290 634 24304 648
rect 6146 610 6160 624
rect 22538 610 22552 624
rect 6122 586 6136 600
rect 10802 586 10816 600
rect 10898 586 10912 600
rect 19058 586 19072 600
rect 19106 586 19120 600
rect 23930 586 23944 600
rect 6074 562 6088 576
rect 6458 562 6472 576
rect 6506 562 6520 576
rect 13802 562 13816 576
rect 13994 562 14008 576
rect 22826 562 22840 576
rect 23594 562 23608 576
rect 26090 562 26104 576
rect 26138 562 26152 576
rect 4970 538 4984 552
rect 16010 538 16024 552
rect 16370 538 16384 552
rect 26821 538 26835 552
rect 4946 514 4960 528
rect 16970 514 16984 528
rect 17066 514 17080 528
rect 23666 514 23680 528
rect 26042 514 26056 528
rect 26114 514 26128 528
rect 4898 490 4912 504
rect 7802 490 7816 504
rect 17498 490 17512 504
rect 20882 490 20896 504
rect 22754 490 22768 504
rect 4658 466 4672 480
rect 22106 466 22120 480
rect 4634 442 4648 456
rect 21098 442 21112 456
rect 4562 418 4576 432
rect 6746 418 6760 432
rect 6794 418 6808 432
rect 26090 418 26104 432
rect 4538 394 4552 408
rect 22322 394 22336 408
rect 22418 394 22432 408
rect 24914 394 24928 408
rect 4466 370 4480 384
rect 8954 370 8968 384
rect 9362 370 9376 384
rect 11474 370 11488 384
rect 12506 370 12520 384
rect 24842 370 24856 384
rect 4442 346 4456 360
rect 25370 346 25384 360
rect 4370 322 4384 336
rect 8762 322 8776 336
rect 8978 322 8992 336
rect 17018 322 17032 336
rect 4178 298 4192 312
rect 4994 298 5008 312
rect 6002 298 6016 312
rect 14018 298 14032 312
rect 15074 298 15088 312
rect 15818 298 15832 312
rect 21866 298 21880 312
rect 4130 274 4144 288
rect 13634 274 13648 288
rect 15218 274 15232 288
rect 18650 274 18664 288
rect 3530 250 3544 264
rect 14642 250 14656 264
rect 3410 226 3424 240
rect 13970 226 13984 240
rect 3362 202 3376 216
rect 10538 202 10552 216
rect 14090 202 14104 216
rect 22874 202 22888 216
rect 3314 178 3328 192
rect 9194 178 9208 192
rect 9698 178 9712 192
rect 19442 178 19456 192
rect 3266 154 3280 168
rect 11114 154 11128 168
rect 20066 154 20080 168
rect 24482 154 24496 168
rect 3122 130 3136 144
rect 9242 130 9256 144
rect 9842 130 9856 144
rect 14570 130 14584 144
rect 2978 106 2992 120
rect 22586 106 22600 120
rect 2498 82 2512 96
rect 21314 82 21328 96
rect 70 58 84 72
rect 1706 58 1720 72
rect 1946 58 1960 72
rect 6554 58 6568 72
rect 6602 58 6616 72
rect 8618 58 8632 72
rect 21194 58 21208 72
rect 26138 58 26152 72
rect 26821 58 26835 72
rect 70 34 84 48
rect 2834 34 2848 48
rect 2882 34 2896 48
rect 18242 34 18256 48
rect 26114 34 26128 48
rect 26821 34 26835 48
rect 7058 10 7072 24
rect 7814 10 7828 24
rect 8258 10 8272 24
rect 13946 10 13960 24
rect 26090 10 26104 24
rect 26821 10 26835 24
<< metal2 >>
rect 0 7821 70 7833
rect 0 7797 70 7809
rect 123 7618 323 7964
rect 339 7618 351 7964
rect 363 7618 375 7964
rect 387 7618 399 7964
rect 411 7618 423 7964
rect 2319 7786 2331 7964
rect 2871 7858 2883 7964
rect 3279 7882 3291 7964
rect 3280 7868 3298 7882
rect 2872 7844 2890 7858
rect 2307 7618 2319 7772
rect 2859 7618 2871 7844
rect 3243 7618 3255 7844
rect 3267 7618 3279 7868
rect 4083 7858 4095 7964
rect 4419 7618 4431 7772
rect 5091 7618 5103 7844
rect 5235 7618 5247 7868
rect 5703 7762 5715 7964
rect 6531 7762 6543 7964
rect 6567 7858 6579 7964
rect 7395 7882 7407 7964
rect 6339 7618 6351 7748
rect 6627 7618 6639 7844
rect 7131 7618 7143 7724
rect 7323 7618 7335 7820
rect 8619 7618 8631 7820
rect 8883 7618 8895 7868
rect 9015 7762 9027 7964
rect 8955 7618 8967 7748
rect 9075 7618 9087 7892
rect 9843 7714 9855 7964
rect 10431 7930 10443 7964
rect 11319 7930 11331 7964
rect 10432 7916 10450 7930
rect 11320 7916 11338 7930
rect 10419 7618 10431 7916
rect 11307 7618 11319 7916
rect 11535 7858 11547 7964
rect 12027 7618 12039 7844
rect 12171 7618 12183 7916
rect 12363 7882 12375 7964
rect 12771 7618 12783 7772
rect 12867 7618 12879 7868
rect 13083 7618 13095 7676
rect 13251 7618 13263 7940
rect 13983 7666 13995 7964
rect 14139 7618 14151 7724
rect 14799 7642 14811 7964
rect 14823 7882 14835 7964
rect 15639 7906 15651 7964
rect 17247 7882 17259 7964
rect 17991 7882 18003 7964
rect 17992 7868 18010 7882
rect 15627 7618 15639 7796
rect 17235 7618 17247 7796
rect 17379 7618 17391 7868
rect 17979 7618 17991 7868
rect 18087 7858 18099 7964
rect 19695 7858 19707 7964
rect 20511 7906 20523 7964
rect 21327 7906 21339 7964
rect 19275 7618 19287 7772
rect 19971 7618 19983 7868
rect 20547 7618 20559 7724
rect 20643 7618 20655 7892
rect 21351 7834 21363 7964
rect 20883 7618 20895 7700
rect 21699 7618 21711 7700
rect 21843 7618 21855 7892
rect 22167 7714 22179 7964
rect 22983 7930 22995 7964
rect 23799 7954 23811 7964
rect 22419 7618 22431 7628
rect 22611 7618 22623 7700
rect 23115 7618 23127 7844
rect 24615 7738 24627 7964
rect 25431 7714 25443 7964
rect 23955 7618 23967 7628
rect 25011 7618 25023 7652
rect 25563 7618 25575 7748
rect 25731 7618 25743 7772
rect 26403 7618 26415 7772
rect 26427 7738 26439 7796
rect 26451 7690 26463 7772
rect 26427 7666 26439 7676
rect 26475 7642 26487 7700
rect 26499 7642 26511 7868
rect 26547 7618 26747 7964
rect 26835 7725 26905 7737
rect 26835 7701 26905 7713
rect 26835 7677 26905 7689
rect 26835 7653 26905 7665
rect 26835 7629 26905 7641
rect 0 3700 70 3712
rect 0 3676 70 3688
rect 123 1841 323 6819
rect 339 1841 351 6819
rect 363 1841 375 6819
rect 387 1841 399 6819
rect 411 1841 423 6819
rect 1611 3737 1623 6819
rect 1635 3785 1647 6819
rect 1659 3833 1671 6819
rect 1707 3881 1719 6819
rect 1731 3905 1743 6819
rect 1779 3929 1791 6819
rect 1827 3953 1839 6819
rect 1851 3977 1863 6819
rect 1611 1841 1623 3651
rect 1635 1841 1647 3747
rect 1659 1841 1671 3795
rect 1707 1841 1719 3843
rect 1875 3809 1887 6819
rect 1755 1841 1767 3627
rect 1779 1841 1791 3603
rect 1827 1841 1839 3579
rect 1899 3569 1911 6819
rect 1947 3809 1959 6819
rect 1995 4001 2007 6819
rect 2067 4025 2079 6819
rect 2115 4049 2127 6819
rect 2187 4073 2199 6819
rect 2211 4097 2223 6819
rect 2259 4121 2271 6819
rect 2355 4145 2367 6819
rect 2307 1841 2319 3771
rect 2427 3617 2439 6819
rect 2451 3905 2463 6819
rect 2475 4169 2487 6819
rect 2523 3593 2535 6819
rect 2547 4217 2559 6819
rect 2571 4241 2583 6819
rect 2619 4265 2631 6819
rect 2355 1841 2367 3531
rect 2523 1841 2535 3507
rect 2547 1841 2559 4179
rect 2643 3641 2655 6819
rect 2667 4289 2679 6819
rect 2715 4313 2727 6819
rect 2739 4337 2751 6819
rect 2763 3617 2775 6819
rect 2787 4385 2799 6819
rect 2595 1841 2607 3483
rect 2619 1841 2631 3459
rect 2667 1841 2679 3435
rect 2715 1841 2727 3411
rect 2739 1841 2751 3387
rect 2787 1841 2799 4347
rect 2835 4145 2847 6819
rect 2859 4409 2871 6819
rect 2883 4433 2895 6819
rect 2931 4457 2943 6819
rect 2955 4169 2967 6819
rect 2979 4481 2991 6819
rect 3027 4529 3039 6819
rect 3051 4553 3063 6819
rect 3075 4577 3087 6819
rect 3099 4601 3111 6819
rect 3147 4625 3159 6819
rect 3171 4649 3183 6819
rect 3195 4673 3207 6819
rect 2955 1841 2967 3363
rect 3003 1841 3015 3339
rect 3027 1841 3039 4491
rect 3243 3905 3255 6819
rect 3267 4697 3279 6819
rect 3075 1841 3087 3315
rect 3099 1841 3111 3291
rect 3171 1841 3183 3267
rect 3195 1841 3207 3891
rect 3291 3401 3303 6819
rect 3339 4721 3351 6819
rect 3363 4745 3375 6819
rect 3387 4769 3399 6819
rect 3219 1841 3231 3243
rect 3291 1841 3303 3219
rect 3387 1841 3399 3507
rect 3435 3209 3447 6819
rect 3459 3185 3471 6819
rect 3507 3161 3519 6819
rect 3555 4793 3567 6819
rect 3579 4817 3591 6819
rect 3603 4841 3615 6819
rect 3651 4865 3663 6819
rect 3675 3281 3687 6819
rect 3699 4889 3711 6819
rect 3747 4913 3759 6819
rect 3795 4337 3807 6819
rect 3867 4889 3879 6819
rect 3891 1841 3903 4851
rect 3915 4265 3927 6819
rect 3987 4937 3999 6819
rect 4011 4961 4023 6819
rect 4059 4985 4071 6819
rect 4107 4337 4119 6819
rect 4131 5009 4143 6819
rect 3939 1841 3951 3123
rect 4083 1841 4095 3099
rect 4107 1841 4119 3075
rect 4155 3065 4167 6819
rect 4203 5033 4215 6819
rect 4227 5057 4239 6819
rect 4203 1841 4215 3531
rect 4251 1841 4263 5067
rect 4275 3041 4287 6819
rect 4347 3617 4359 6819
rect 4371 5105 4383 6819
rect 4443 5129 4455 6819
rect 4515 5153 4527 6819
rect 4539 5177 4551 6819
rect 4587 5201 4599 6819
rect 4299 1841 4311 3003
rect 4323 1841 4335 2979
rect 4347 1841 4359 2955
rect 4419 1841 4431 2931
rect 4515 1841 4527 2979
rect 4611 1841 4623 5211
rect 4635 4097 4647 6819
rect 4683 5249 4695 6819
rect 4755 5321 4767 6819
rect 4803 5369 4815 6819
rect 4875 5393 4887 6819
rect 4899 5417 4911 6819
rect 4707 1841 4719 5259
rect 4731 1841 4743 5283
rect 4755 1841 4767 3027
rect 4779 1841 4791 5331
rect 4803 1841 4815 3027
rect 4851 1841 4863 2907
rect 4875 1841 4887 3507
rect 4899 2945 4911 5379
rect 4923 3953 4935 6819
rect 4971 3617 4983 6819
rect 5019 5393 5031 6819
rect 5091 5105 5103 6819
rect 5139 3953 5151 6819
rect 5043 1841 5055 3819
rect 5091 1841 5103 3291
rect 5163 1841 5175 4011
rect 5187 1841 5199 4731
rect 5211 4145 5223 6819
rect 5235 3617 5247 6819
rect 5235 1841 5247 2883
rect 5259 2873 5271 6819
rect 5307 3545 5319 6819
rect 5331 3737 5343 6819
rect 5355 5441 5367 6819
rect 5403 3737 5415 6819
rect 5427 5465 5439 6819
rect 5451 5513 5463 6819
rect 5475 5537 5487 6819
rect 5283 1841 5295 2835
rect 5307 1841 5319 2811
rect 5331 1841 5343 2787
rect 5451 1841 5463 5475
rect 5499 5297 5511 6819
rect 5547 5297 5559 6819
rect 5571 2777 5583 6819
rect 5595 5561 5607 6819
rect 5643 3881 5655 6819
rect 5691 3425 5703 6819
rect 5763 5585 5775 6819
rect 5787 5609 5799 6819
rect 5811 5009 5823 6819
rect 5859 2969 5871 6819
rect 5883 4649 5895 6819
rect 5907 5009 5919 6819
rect 5931 5633 5943 6819
rect 5979 5465 5991 6819
rect 6003 3017 6015 6819
rect 6051 5657 6063 6819
rect 6099 4577 6111 6819
rect 5811 1841 5823 2739
rect 5859 1841 5871 2715
rect 6003 1841 6015 2763
rect 6051 1841 6063 2763
rect 6099 1841 6111 2691
rect 6147 2681 6159 6819
rect 6219 5705 6231 6819
rect 6195 1841 6207 3915
rect 6219 1841 6231 5667
rect 6243 3233 6255 6819
rect 6267 3929 6279 6819
rect 6315 3473 6327 6819
rect 6339 5729 6351 6819
rect 6315 1841 6327 2643
rect 6339 1841 6351 3507
rect 6363 2825 6375 5715
rect 6387 4313 6399 6819
rect 6435 5729 6447 6819
rect 6459 5753 6471 6819
rect 6363 1841 6375 2619
rect 6411 1841 6423 3651
rect 6435 1841 6447 4923
rect 6483 2609 6495 6819
rect 6531 5777 6543 6819
rect 6555 5801 6567 6819
rect 6579 2585 6591 6819
rect 6627 2561 6639 6819
rect 6651 1841 6663 2547
rect 6675 2537 6687 6819
rect 6699 1841 6711 2547
rect 6723 2513 6735 6819
rect 6771 1841 6783 5811
rect 6795 5513 6807 6819
rect 6819 4865 6831 6819
rect 6843 5849 6855 6819
rect 6843 1841 6855 4419
rect 6867 1841 6879 5523
rect 6891 5297 6903 6819
rect 6915 2489 6927 6819
rect 6939 5873 6951 6819
rect 6987 5897 6999 6819
rect 7011 5921 7023 6819
rect 7035 5945 7047 6819
rect 7059 5969 7071 6819
rect 6939 1841 6951 4851
rect 7107 3113 7119 6819
rect 7155 6017 7167 6819
rect 7203 6065 7215 6819
rect 6963 1841 6975 2451
rect 6987 1841 6999 2427
rect 7059 1841 7071 2475
rect 7107 1841 7119 2475
rect 7155 1841 7167 5979
rect 7179 1841 7191 2403
rect 7203 1841 7215 6027
rect 7227 4649 7239 6819
rect 7251 5129 7263 6819
rect 7275 6089 7287 6819
rect 7251 1841 7263 4803
rect 7275 1841 7287 5235
rect 7323 2393 7335 6819
rect 7371 2465 7383 6819
rect 7395 5249 7407 6819
rect 7419 2417 7431 6819
rect 7467 6113 7479 6819
rect 7491 6137 7503 6819
rect 7371 1841 7383 2355
rect 7395 1841 7407 2379
rect 7443 1841 7455 2715
rect 7467 1841 7479 2379
rect 7515 2345 7527 6819
rect 7563 6161 7575 6819
rect 7539 1841 7551 4203
rect 7587 4049 7599 6819
rect 7611 6185 7623 6819
rect 7659 4865 7671 6819
rect 7683 6209 7695 6819
rect 7707 6137 7719 6819
rect 7563 1841 7575 3891
rect 7755 3785 7767 6819
rect 7779 6137 7791 6819
rect 7587 1841 7599 2307
rect 7635 1841 7647 3555
rect 7683 1841 7695 3555
rect 7791 2297 7803 6051
rect 7827 2297 7839 6819
rect 7875 4289 7887 6819
rect 7899 6065 7911 6819
rect 7923 6233 7935 6819
rect 7971 6209 7983 6819
rect 7755 1841 7767 2283
rect 7803 1841 7815 2259
rect 7851 1841 7863 3699
rect 7923 2249 7935 6195
rect 7995 3305 8007 6819
rect 8019 6257 8031 6819
rect 8067 6281 8079 6819
rect 8091 6305 8103 6819
rect 8115 5561 8127 6819
rect 8139 5489 8151 6819
rect 8187 5489 8199 6819
rect 8211 6065 8223 6819
rect 8235 6329 8247 6819
rect 7899 1841 7911 2235
rect 7971 1841 7983 2235
rect 7995 1841 8007 2211
rect 8019 1841 8031 4683
rect 8091 1841 8103 2811
rect 8139 1841 8151 2907
rect 8211 1841 8223 4443
rect 8235 1841 8247 5547
rect 8283 5465 8295 6819
rect 8307 2465 8319 6819
rect 8331 5417 8343 6819
rect 8355 6353 8367 6819
rect 8403 6305 8415 6819
rect 8307 1841 8319 2187
rect 8331 1841 8343 2163
rect 8355 1841 8367 6291
rect 8427 4241 8439 6819
rect 8451 6401 8463 6819
rect 8403 1841 8415 3651
rect 8427 1841 8439 2427
rect 8451 1841 8463 6363
rect 8499 4241 8511 6819
rect 8523 5465 8535 6819
rect 8571 3665 8583 6819
rect 8523 1841 8535 2139
rect 8547 1841 8559 2475
rect 8619 2129 8631 6819
rect 8667 6065 8679 6819
rect 8691 6425 8703 6819
rect 8715 6449 8727 6819
rect 8763 4433 8775 6819
rect 8571 1841 8583 2115
rect 8667 1841 8679 2115
rect 8739 1841 8751 2091
rect 8787 1841 8799 6459
rect 8811 2249 8823 6819
rect 8883 6473 8895 6819
rect 8931 6473 8943 6819
rect 8955 6497 8967 6819
rect 8835 1841 8847 2067
rect 8859 1841 8871 5499
rect 8883 1841 8895 4515
rect 8931 1841 8943 4467
rect 8955 2921 8967 6459
rect 8979 5609 8991 6819
rect 9027 6473 9039 6819
rect 9051 6521 9063 6819
rect 9027 1841 9039 3723
rect 9051 1841 9063 3531
rect 9075 1841 9087 5499
rect 9099 1841 9111 4851
rect 9123 4337 9135 6819
rect 9147 5417 9159 6819
rect 9171 6545 9183 6819
rect 9171 1841 9183 5763
rect 9219 2657 9231 6819
rect 9267 6569 9279 6819
rect 9339 4265 9351 6819
rect 9363 5705 9375 6819
rect 9387 3545 9399 6819
rect 9411 5825 9423 6819
rect 9459 4217 9471 6819
rect 9219 1841 9231 2043
rect 9267 1841 9279 2019
rect 9411 1841 9423 3795
rect 9459 1841 9471 3819
rect 9483 2945 9495 6819
rect 9507 5009 9519 6819
rect 9531 5825 9543 6819
rect 9579 4817 9591 6819
rect 9483 1841 9495 1995
rect 9507 1841 9519 4251
rect 9555 1841 9567 3795
rect 9579 1841 9591 3891
rect 9603 3233 9615 6819
rect 9627 6593 9639 6819
rect 9627 2009 9639 6051
rect 9675 4865 9687 6819
rect 9699 2441 9711 6819
rect 9723 6617 9735 6819
rect 9603 1841 9615 1971
rect 9723 1841 9735 5187
rect 9771 3017 9783 6819
rect 9795 6641 9807 6819
rect 9747 1841 9759 1995
rect 9795 1841 9807 4059
rect 9819 3401 9831 6819
rect 9819 1841 9831 3123
rect 9843 2777 9855 6819
rect 9867 2993 9879 6627
rect 9891 5633 9903 6819
rect 9915 4217 9927 6819
rect 9939 5633 9951 6819
rect 9987 6641 9999 6819
rect 10011 6497 10023 6819
rect 10035 5225 10047 6819
rect 10083 5201 10095 6819
rect 9915 1841 9927 2979
rect 9939 1841 9951 4947
rect 10011 1841 10023 4731
rect 10035 1841 10047 4707
rect 10107 4001 10119 6819
rect 10131 5201 10143 6819
rect 10155 3689 10167 6819
rect 10203 5225 10215 6819
rect 10059 1841 10071 2763
rect 10227 2417 10239 6819
rect 10251 6665 10263 6819
rect 10131 1841 10143 1947
rect 10251 1841 10263 5811
rect 10275 1841 10287 6531
rect 10299 4913 10311 6819
rect 10323 4169 10335 6819
rect 10371 4721 10383 6819
rect 10419 5825 10431 6819
rect 10371 1841 10383 3987
rect 10395 1841 10407 2811
rect 10443 1841 10455 5019
rect 10467 3137 10479 6819
rect 10491 3233 10503 6819
rect 10539 5465 10551 6819
rect 10515 4001 10527 4755
rect 10563 1937 10575 6507
rect 10587 2465 10599 6819
rect 10611 4769 10623 6819
rect 10635 5033 10647 6819
rect 10683 6545 10695 6819
rect 10491 1841 10503 1923
rect 10611 1841 10623 3987
rect 10635 1841 10647 2403
rect 10659 2369 10671 5019
rect 10707 3737 10719 6819
rect 10683 1841 10695 3675
rect 10731 1841 10743 4923
rect 10755 4241 10767 6819
rect 10755 1841 10767 2067
rect 10779 1841 10791 4995
rect 10803 4337 10815 6819
rect 10827 4985 10839 6819
rect 10851 4553 10863 6819
rect 10899 5705 10911 6819
rect 10923 5465 10935 6819
rect 10851 1841 10863 2571
rect 10875 1841 10887 3723
rect 10947 1841 10959 6051
rect 10971 5033 10983 6819
rect 10971 1841 10983 3123
rect 10995 1841 11007 6195
rect 11019 6065 11031 6819
rect 11043 5369 11055 6819
rect 11067 5945 11079 6819
rect 11139 6065 11151 6819
rect 11043 1841 11055 3291
rect 11067 1841 11079 4635
rect 11091 2993 11103 5019
rect 11163 4241 11175 6819
rect 11211 5033 11223 6819
rect 11163 1841 11175 4107
rect 11211 1841 11223 2571
rect 11235 2417 11247 6819
rect 11307 6689 11319 6819
rect 11283 1841 11295 2355
rect 11307 1841 11319 5931
rect 11331 2129 11343 6675
rect 11355 1937 11367 6819
rect 11379 1841 11391 5403
rect 11403 4217 11415 6819
rect 11475 6689 11487 6819
rect 11499 5537 11511 6819
rect 11547 4745 11559 6819
rect 11595 6713 11607 6819
rect 11403 1841 11415 2115
rect 11427 1841 11439 4227
rect 11451 1841 11463 3627
rect 11523 1841 11535 4203
rect 11547 1841 11559 2931
rect 11571 1841 11583 4947
rect 11619 3641 11631 6819
rect 11643 6737 11655 6819
rect 11691 6761 11703 6819
rect 11595 1841 11607 2475
rect 11643 2129 11655 4851
rect 11643 1841 11655 1899
rect 11691 1841 11703 6651
rect 11739 3329 11751 6819
rect 11811 3953 11823 6819
rect 11835 3905 11847 6819
rect 11859 6665 11871 6819
rect 11907 4169 11919 6819
rect 11931 2825 11943 6819
rect 11955 2129 11967 6819
rect 12003 6785 12015 6819
rect 12027 2897 12039 6819
rect 12075 2153 12087 6819
rect 12123 3089 12135 6819
rect 12243 5081 12255 6819
rect 12267 2897 12279 6819
rect 12315 5993 12327 6819
rect 12363 5081 12375 6819
rect 12387 5993 12399 6819
rect 12411 6329 12423 6819
rect 12435 5801 12447 6819
rect 12459 6329 12471 6819
rect 12363 1841 12375 4635
rect 12387 1841 12399 3531
rect 12435 1841 12447 4803
rect 12483 1841 12495 5619
rect 12507 4697 12519 6819
rect 12555 5537 12567 6819
rect 12531 2801 12543 5067
rect 12627 4289 12639 6819
rect 12651 6761 12663 6819
rect 12675 4793 12687 6819
rect 12723 4409 12735 6819
rect 12747 4793 12759 6819
rect 12795 5081 12807 6819
rect 12555 1841 12567 2139
rect 12747 1841 12759 4275
rect 12843 3041 12855 6819
rect 12867 4121 12879 6819
rect 12915 6473 12927 6819
rect 12963 4481 12975 6819
rect 13011 5057 13023 6819
rect 12771 1841 12783 2787
rect 12819 1841 12831 2187
rect 12843 1841 12855 1875
rect 12915 1841 12927 4155
rect 12963 1841 12975 4155
rect 13035 1841 13047 3219
rect 13059 1841 13071 5379
rect 13083 1889 13095 6819
rect 13131 2993 13143 6819
rect 13155 3545 13167 6819
rect 13179 5345 13191 6819
rect 13107 1841 13119 2835
rect 13155 1841 13167 3027
rect 13179 1841 13191 2763
rect 13203 1841 13215 4107
rect 13227 3113 13239 6819
rect 13251 2729 13263 6819
rect 13275 6281 13287 6819
rect 13287 3041 13299 5379
rect 13323 3833 13335 6819
rect 13347 5249 13359 6819
rect 13371 4649 13383 6819
rect 13395 3353 13407 6819
rect 13443 5465 13455 6819
rect 13419 3041 13431 5067
rect 13467 3305 13479 6819
rect 13323 1841 13335 3027
rect 13347 1841 13359 2715
rect 13443 1841 13455 1875
rect 13467 1841 13479 3027
rect 13491 2729 13503 6147
rect 13515 2081 13527 6819
rect 13515 1841 13527 1851
rect 13539 1841 13551 4923
rect 13563 2081 13575 6819
rect 13587 6545 13599 6819
rect 13587 1841 13599 5019
rect 13611 4913 13623 6819
rect 13635 1889 13647 6339
rect 13659 3041 13671 5811
rect 13683 1841 13695 5859
rect 13731 4481 13743 6819
rect 13707 1841 13719 3027
rect 13755 1841 13767 2331
rect 13779 1841 13791 3531
rect 13851 1841 13863 2715
rect 13875 1841 13887 5931
rect 13899 1841 13911 2643
rect 14091 2393 14103 6819
rect 14043 1841 14055 2187
rect 14115 1841 14127 2643
rect 14139 1841 14151 2379
rect 14211 1841 14223 3291
rect 14331 1841 14343 5403
rect 14355 4913 14367 6819
rect 14355 1841 14367 3939
rect 14379 2033 14391 4899
rect 14403 1841 14415 3267
rect 14475 1841 14487 2331
rect 14523 1841 14535 2019
rect 14619 1841 14631 6195
rect 14715 4649 14727 6819
rect 14763 6545 14775 6819
rect 14715 1841 14727 1875
rect 14763 1841 14775 5979
rect 14811 1841 14823 4923
rect 14835 1841 14847 4323
rect 14859 1841 14871 4731
rect 14883 1841 14895 5211
rect 14907 2633 14919 6819
rect 14931 4745 14943 6819
rect 14955 4913 14967 6819
rect 14931 1841 14943 4227
rect 14955 1841 14967 3771
rect 14979 1889 14991 4899
rect 15003 3137 15015 6819
rect 15027 3233 15039 6819
rect 15051 4097 15063 6819
rect 15099 4913 15111 6819
rect 15123 6089 15135 6819
rect 15147 5033 15159 6819
rect 15171 6449 15183 6819
rect 15195 5057 15207 6819
rect 15243 5849 15255 6819
rect 15267 5081 15279 6819
rect 15291 4673 15303 6819
rect 15315 6593 15327 6819
rect 15003 1841 15015 2451
rect 15051 1841 15063 3243
rect 15099 1841 15111 4083
rect 15339 3857 15351 6819
rect 15387 4673 15399 6819
rect 15411 4385 15423 6819
rect 15435 5225 15447 6819
rect 15459 4385 15471 6819
rect 15483 5345 15495 6819
rect 15531 6113 15543 6819
rect 15555 6569 15567 6819
rect 15579 5633 15591 6819
rect 15603 5825 15615 6819
rect 15675 4265 15687 6819
rect 15699 5849 15711 6819
rect 15723 5873 15735 6819
rect 15747 6209 15759 6819
rect 15771 5945 15783 6819
rect 15771 1841 15783 4923
rect 15795 1841 15807 4995
rect 15819 4961 15831 6819
rect 15843 2921 15855 6819
rect 15867 5993 15879 6819
rect 15891 1841 15903 5523
rect 15915 2249 15927 6819
rect 15939 5537 15951 6819
rect 15987 6089 15999 6819
rect 15915 1841 15927 1875
rect 15963 1841 15975 3651
rect 15987 1841 15999 3003
rect 16011 1889 16023 6699
rect 16035 6497 16047 6819
rect 16059 3905 16071 6819
rect 16107 6713 16119 6819
rect 16059 1841 16071 3843
rect 16083 1865 16095 6075
rect 16107 1841 16119 6675
rect 16131 3857 16143 4419
rect 16155 3377 16167 6819
rect 16179 3905 16191 6819
rect 16155 1841 16167 3123
rect 16203 1841 16215 4251
rect 16227 2897 16239 6819
rect 16251 3137 16263 4515
rect 16275 4433 16287 6819
rect 16299 4529 16311 6819
rect 16275 1841 16287 3675
rect 16323 3473 16335 6819
rect 16347 5489 16359 6819
rect 16371 3857 16383 6507
rect 16395 5417 16407 6819
rect 16419 5465 16431 6819
rect 16323 1841 16335 2499
rect 16347 1841 16359 3843
rect 16419 1841 16431 3843
rect 16443 2465 16455 6819
rect 16467 3905 16479 6819
rect 16491 3977 16503 6819
rect 16539 4649 16551 6819
rect 16563 3233 16575 6819
rect 16611 5465 16623 6819
rect 16515 1841 16527 3123
rect 16563 1841 16575 3147
rect 16587 1841 16599 3963
rect 16635 3857 16647 6051
rect 16659 5105 16671 6819
rect 16683 6497 16695 6819
rect 16659 1841 16671 4275
rect 16707 3473 16719 6819
rect 16779 1841 16791 2667
rect 16803 1841 16815 3531
rect 16827 3041 16839 6819
rect 16875 1841 16887 5523
rect 16899 1841 16911 4635
rect 16923 1841 16935 5643
rect 16947 1841 16959 3891
rect 17043 1841 17055 3507
rect 17115 1841 17127 4323
rect 17139 1841 17151 4299
rect 17211 1841 17223 3411
rect 17235 3089 17247 6819
rect 17235 1841 17247 2955
rect 17307 1841 17319 3099
rect 17331 1841 17343 4779
rect 17379 4361 17391 6819
rect 17427 5489 17439 6819
rect 17451 5897 17463 6819
rect 17403 1841 17415 2859
rect 17427 1841 17439 5091
rect 17475 2417 17487 6819
rect 17499 3785 17511 6819
rect 17523 1913 17535 6819
rect 17571 5465 17583 6819
rect 17595 4361 17607 6819
rect 17619 5849 17631 6819
rect 17667 5849 17679 6819
rect 17691 3641 17703 6819
rect 17715 5585 17727 6819
rect 17763 5585 17775 6819
rect 17547 1841 17559 2763
rect 17619 1841 17631 2307
rect 17739 1841 17751 3939
rect 17787 3905 17799 6819
rect 17811 6089 17823 6819
rect 17763 1841 17775 3603
rect 17787 1841 17799 3843
rect 17835 1841 17847 2979
rect 17859 2465 17871 6819
rect 17883 6065 17895 6819
rect 17931 6161 17943 6819
rect 17859 1841 17871 2403
rect 17883 1841 17895 4299
rect 17907 3857 17919 5307
rect 17931 1841 17943 3819
rect 17955 1841 17967 6531
rect 17979 2009 17991 6819
rect 18027 6497 18039 6819
rect 18051 3905 18063 6819
rect 18003 1841 18015 3195
rect 18051 1841 18063 2115
rect 18075 1841 18087 6531
rect 18147 6281 18159 6819
rect 18099 1841 18111 3507
rect 18123 1841 18135 3843
rect 18159 2417 18171 4083
rect 18219 2321 18231 6819
rect 18243 4121 18255 6819
rect 18267 2441 18279 6819
rect 18315 4241 18327 6819
rect 18339 5249 18351 6819
rect 18363 4577 18375 6819
rect 18411 6353 18423 6819
rect 18435 2273 18447 6819
rect 18483 5633 18495 6819
rect 18531 5633 18543 6819
rect 18579 4937 18591 6819
rect 18651 5849 18663 6819
rect 18675 4457 18687 6819
rect 18699 3641 18711 6819
rect 18723 4673 18735 6819
rect 18771 2081 18783 6819
rect 18795 4673 18807 6819
rect 18819 6449 18831 6819
rect 18795 1841 18807 4635
rect 18819 1841 18831 5643
rect 18867 3449 18879 6819
rect 18891 3593 18903 6819
rect 18915 4025 18927 6819
rect 18843 1841 18855 3387
rect 18867 1841 18879 3411
rect 18915 1841 18927 3819
rect 18939 1841 18951 6603
rect 18963 2849 18975 6819
rect 18987 3641 18999 6819
rect 19011 2729 19023 6819
rect 18963 1841 18975 2667
rect 19035 1841 19047 3915
rect 19059 2945 19071 6819
rect 19083 3281 19095 6819
rect 19083 1841 19095 3195
rect 19107 2705 19119 6819
rect 19131 4097 19143 4659
rect 19155 3737 19167 6819
rect 19179 4673 19191 6819
rect 19203 3977 19215 6819
rect 19251 4409 19263 6819
rect 19155 1841 19167 3579
rect 19179 1841 19191 3891
rect 19227 1841 19239 2931
rect 19275 1841 19287 6483
rect 19299 3833 19311 6747
rect 19323 5009 19335 6819
rect 19335 3593 19347 4323
rect 19371 3545 19383 6819
rect 19323 1841 19335 3507
rect 19395 2993 19407 6819
rect 19419 3281 19431 6819
rect 19443 3881 19455 6819
rect 19491 4937 19503 6819
rect 19467 2681 19479 4755
rect 19515 4697 19527 6819
rect 19563 4961 19575 6819
rect 19395 1841 19407 2187
rect 19515 1841 19527 2931
rect 19539 1841 19551 3003
rect 19563 1841 19575 4011
rect 19587 3209 19599 5427
rect 19611 3545 19623 6819
rect 19635 3665 19647 6819
rect 19659 5417 19671 6819
rect 19611 1841 19623 3387
rect 19683 3377 19695 6819
rect 19707 3233 19719 4659
rect 19731 3497 19743 6819
rect 19779 4457 19791 6819
rect 19659 1841 19671 2955
rect 19731 1841 19743 3459
rect 19755 1841 19767 3603
rect 19779 1841 19791 3795
rect 19803 3473 19815 5571
rect 19827 1841 19839 5091
rect 19851 4049 19863 6819
rect 19851 1841 19863 3963
rect 19875 1865 19887 6819
rect 19899 6473 19911 6819
rect 19899 1841 19911 6123
rect 19923 3977 19935 4683
rect 19947 2201 19959 6819
rect 19947 1841 19959 2115
rect 19971 1841 19983 5523
rect 19995 2345 20007 6819
rect 19995 1841 20007 2307
rect 20019 2105 20031 6459
rect 20043 4193 20055 6819
rect 20067 5393 20079 6819
rect 20091 4529 20103 6819
rect 20139 6761 20151 6819
rect 20043 1841 20055 3963
rect 20103 2129 20115 4251
rect 20139 1841 20151 5979
rect 20163 4889 20175 6819
rect 20187 4625 20199 6819
rect 20163 1841 20175 3507
rect 20187 1841 20199 4179
rect 20211 3977 20223 6219
rect 20235 3521 20247 6819
rect 20259 3617 20271 6819
rect 20307 5849 20319 6819
rect 20355 6257 20367 6819
rect 20379 6545 20391 6819
rect 20283 3473 20295 5427
rect 20235 1841 20247 3459
rect 20307 1841 20319 3171
rect 20355 1841 20367 6195
rect 20379 1841 20391 4635
rect 20403 2057 20415 6819
rect 20427 1841 20439 6099
rect 20451 4337 20463 6819
rect 20475 6497 20487 6819
rect 20499 5273 20511 6819
rect 20475 1841 20487 2547
rect 20523 1841 20535 3963
rect 20571 2753 20583 6819
rect 20595 5273 20607 6819
rect 20595 1841 20607 4947
rect 20619 1841 20631 4995
rect 20643 4505 20655 6819
rect 20667 1841 20679 5571
rect 20691 3257 20703 6819
rect 20715 5633 20727 6819
rect 20715 1841 20727 4203
rect 20739 3761 20751 6819
rect 20763 4289 20775 5259
rect 20787 4505 20799 6819
rect 20811 5105 20823 6819
rect 20835 6113 20847 6819
rect 20739 1841 20751 3651
rect 20787 1841 20799 3003
rect 20835 1841 20847 6051
rect 20859 1841 20871 4635
rect 20883 3977 20895 6819
rect 20907 3665 20919 5379
rect 20931 2657 20943 6819
rect 20955 4529 20967 6819
rect 20979 5753 20991 6819
rect 20955 1841 20967 4203
rect 20979 1841 20991 4155
rect 21003 1841 21015 5619
rect 21027 4649 21039 6819
rect 21051 6113 21063 6819
rect 21075 6809 21087 6819
rect 21051 1841 21063 5379
rect 21075 1841 21087 6699
rect 21099 2777 21111 4491
rect 21123 3233 21135 6819
rect 21147 4865 21159 6819
rect 21171 6761 21183 6819
rect 21147 1841 21159 4035
rect 21171 1841 21183 4947
rect 21195 1937 21207 6099
rect 21291 5273 21303 6819
rect 21219 3953 21231 4515
rect 21243 1841 21255 3891
rect 21267 1841 21279 3531
rect 21291 1841 21303 5091
rect 21315 2033 21327 5259
rect 21363 1841 21375 5331
rect 21483 1841 21495 4131
rect 21507 1841 21519 4395
rect 21603 1841 21615 3603
rect 21627 1841 21639 4683
rect 21651 2225 21663 6819
rect 21699 4793 21711 6819
rect 21843 6041 21855 6819
rect 21723 1841 21735 5787
rect 21795 1841 21807 5883
rect 21867 4289 21879 6531
rect 21843 1841 21855 4275
rect 21891 2825 21903 6819
rect 21915 6281 21927 6819
rect 21915 1841 21927 5499
rect 21939 5105 21951 6819
rect 21963 5729 21975 6819
rect 22011 5249 22023 6819
rect 21963 1841 21975 2979
rect 21987 1841 21999 4971
rect 22035 3305 22047 6819
rect 22059 5177 22071 6819
rect 22107 5057 22119 6819
rect 22155 5921 22167 6819
rect 22035 1841 22047 3267
rect 22083 1841 22095 4443
rect 22131 1841 22143 4275
rect 22179 1841 22191 4227
rect 22203 1841 22215 6195
rect 22227 4025 22239 6819
rect 22251 2489 22263 6819
rect 22275 3689 22287 6819
rect 22299 4457 22311 6819
rect 22275 1841 22287 3243
rect 22347 2321 22359 6819
rect 22371 2105 22383 6819
rect 22395 5633 22407 6819
rect 22467 6809 22479 6819
rect 22395 1841 22407 5523
rect 22419 2585 22431 5619
rect 22443 1841 22455 2979
rect 22467 1841 22479 3699
rect 22491 2081 22503 6819
rect 22515 2153 22527 6819
rect 22539 4121 22551 6819
rect 22563 3113 22575 6819
rect 22611 3281 22623 6819
rect 22659 6449 22671 6819
rect 22659 1841 22671 4635
rect 22683 2489 22695 6819
rect 22707 3569 22719 6819
rect 22731 4577 22743 6819
rect 22755 4505 22767 6819
rect 22683 1841 22695 2451
rect 22707 1841 22719 3459
rect 22779 1841 22791 4323
rect 22803 3521 22815 6819
rect 22827 4721 22839 6819
rect 22851 3953 22863 6819
rect 22875 4529 22887 6819
rect 22923 6161 22935 6819
rect 22803 1841 22815 3387
rect 22899 1841 22911 2763
rect 22923 1841 22935 4131
rect 22947 2297 22959 6819
rect 22971 2465 22983 6051
rect 22995 5033 23007 6819
rect 23043 5993 23055 6819
rect 23019 3473 23031 5475
rect 23043 1841 23055 5931
rect 23067 4529 23079 6819
rect 23091 4289 23103 6819
rect 23163 6281 23175 6819
rect 23115 3401 23127 5379
rect 23139 4145 23151 5979
rect 23187 5105 23199 6819
rect 23211 5561 23223 6819
rect 23259 6017 23271 6819
rect 23283 4529 23295 6819
rect 23307 4625 23319 6819
rect 23331 4481 23343 6819
rect 23379 1985 23391 6819
rect 23403 3737 23415 6819
rect 23427 3521 23439 6819
rect 23451 6113 23463 6819
rect 23403 1841 23415 3219
rect 23451 1841 23463 6051
rect 23475 3137 23487 6099
rect 23499 2777 23511 6819
rect 23523 3809 23535 6819
rect 23547 3905 23559 6819
rect 23571 6425 23583 6819
rect 23619 6089 23631 6819
rect 23595 1841 23607 4275
rect 23643 4217 23655 6819
rect 23667 4481 23679 6819
rect 23715 4121 23727 6819
rect 23763 5417 23775 6819
rect 23835 6665 23847 6819
rect 23787 4217 23799 6531
rect 23859 5321 23871 6819
rect 23883 6641 23895 6819
rect 23691 1841 23703 3051
rect 23715 1841 23727 2523
rect 23763 1841 23775 4203
rect 23811 1841 23823 4899
rect 23931 2201 23943 6819
rect 23979 4529 23991 6819
rect 24027 4649 24039 6819
rect 24051 2081 24063 6819
rect 24075 4097 24087 6819
rect 24099 4001 24111 6819
rect 24147 4337 24159 6819
rect 24171 2825 24183 6819
rect 24195 3497 24207 6819
rect 24243 3305 24255 6819
rect 24267 6545 24279 6819
rect 24291 4073 24303 6819
rect 24339 5705 24351 6819
rect 24363 5129 24375 6819
rect 24387 4745 24399 6819
rect 24435 6305 24447 6819
rect 24459 4481 24471 6819
rect 24483 4121 24495 6819
rect 24507 4361 24519 6819
rect 24555 6377 24567 6819
rect 24339 1841 24351 3723
rect 24507 1841 24519 3315
rect 24531 1841 24543 5859
rect 24579 4889 24591 6819
rect 24603 6233 24615 6819
rect 24579 1841 24591 4803
rect 24603 1841 24615 6195
rect 24627 3353 24639 6819
rect 24651 6785 24663 6819
rect 24699 4865 24711 6819
rect 24723 4241 24735 6819
rect 24675 1841 24687 3891
rect 24723 1841 24735 3627
rect 24747 2441 24759 6819
rect 24771 5081 24783 6819
rect 24819 5105 24831 6819
rect 24843 4169 24855 6819
rect 24795 1841 24807 2595
rect 24819 1841 24831 3603
rect 24867 3521 24879 6819
rect 24891 2825 24903 6819
rect 24915 6305 24927 6819
rect 24963 6185 24975 6819
rect 24891 1841 24903 2067
rect 24939 1841 24951 4371
rect 24987 4361 24999 6819
rect 24987 1841 24999 3435
rect 25011 1841 25023 6723
rect 25035 1841 25047 5211
rect 25059 2801 25071 6819
rect 25083 5009 25095 6819
rect 25107 6257 25119 6819
rect 25083 1841 25095 4203
rect 25107 1841 25119 6195
rect 25155 5849 25167 6819
rect 25131 3425 25143 4875
rect 25155 1841 25167 5787
rect 25179 4697 25191 6819
rect 25227 5297 25239 6819
rect 25203 1841 25215 5283
rect 25275 4649 25287 6819
rect 25239 2585 25251 4347
rect 25299 3737 25311 6819
rect 25347 5705 25359 6819
rect 25371 4217 25383 6747
rect 25359 3713 25371 3939
rect 25299 1841 25311 3699
rect 25323 1841 25335 3603
rect 25395 3329 25407 6819
rect 25419 5705 25431 6819
rect 25419 1841 25431 3771
rect 25443 3545 25455 6819
rect 25443 1841 25455 3507
rect 25467 2561 25479 6819
rect 25467 1841 25479 2523
rect 25491 2393 25503 6219
rect 25515 4841 25527 6819
rect 25539 5393 25551 6819
rect 25515 1841 25527 4323
rect 25539 1841 25551 5355
rect 25563 1841 25575 6507
rect 25587 1961 25599 6243
rect 25611 3857 25623 6819
rect 25635 6065 25647 6819
rect 25611 1841 25623 3723
rect 25635 1841 25647 2835
rect 25659 2369 25671 6819
rect 25659 1841 25671 2331
rect 25683 1841 25695 6339
rect 25707 4409 25719 6819
rect 25731 1841 25743 5643
rect 25755 4937 25767 6819
rect 25755 1841 25767 4635
rect 25779 1841 25791 5187
rect 25803 4265 25815 5835
rect 25827 4865 25839 6819
rect 25827 1841 25839 4227
rect 25851 3737 25863 6819
rect 25851 1841 25863 3315
rect 25875 1841 25887 5139
rect 25899 3545 25911 6819
rect 25923 5825 25935 6819
rect 25923 1841 25935 5595
rect 25947 3521 25959 6699
rect 25995 4721 26007 6819
rect 26019 4193 26031 6819
rect 26067 5681 26079 6819
rect 26115 5465 26127 6819
rect 26139 6401 26151 6819
rect 26163 5777 26175 6819
rect 26211 5297 26223 6819
rect 25971 1841 25983 2643
rect 26043 1841 26055 4587
rect 26091 1841 26103 4323
rect 26175 2537 26187 4419
rect 26235 4289 26247 6819
rect 26259 4625 26271 6819
rect 26283 4313 26295 5379
rect 26307 4553 26319 6819
rect 26331 4577 26343 6819
rect 26355 4337 26367 6819
rect 26379 2345 26391 5571
rect 26403 2177 26415 6819
rect 26427 1865 26439 4443
rect 26451 1889 26463 5955
rect 26547 1841 26747 6819
rect 26835 6316 26905 6328
rect 26835 4492 26905 4504
rect 26835 1876 26905 1888
rect 26835 1852 26905 1864
rect 0 59 70 71
rect 0 35 70 47
rect 123 0 323 1042
rect 339 0 351 1042
rect 363 0 375 1042
rect 387 0 399 1042
rect 411 0 423 1042
rect 1707 72 1719 1042
rect 1947 72 1959 1042
rect 2499 96 2511 1042
rect 2835 48 2847 1042
rect 2883 48 2895 1042
rect 2979 120 2991 1042
rect 3123 144 3135 1042
rect 3267 168 3279 1042
rect 3315 192 3327 1042
rect 3363 216 3375 1042
rect 3411 240 3423 1042
rect 3531 264 3543 1042
rect 4131 288 4143 1042
rect 4179 312 4191 1042
rect 4371 336 4383 1042
rect 4443 360 4455 1042
rect 4467 384 4479 1042
rect 4539 408 4551 1042
rect 4563 432 4575 1042
rect 4635 456 4647 1042
rect 4659 480 4671 1042
rect 4899 504 4911 1042
rect 4947 528 4959 1042
rect 4971 552 4983 1042
rect 4995 312 5007 1042
rect 6003 312 6015 1042
rect 6075 576 6087 1042
rect 6123 600 6135 1042
rect 6147 624 6159 1042
rect 6267 648 6279 1042
rect 6459 576 6471 1042
rect 6507 576 6519 1042
rect 6531 672 6543 1042
rect 6555 72 6567 1042
rect 6603 72 6615 1042
rect 6627 696 6639 1042
rect 6723 720 6735 1042
rect 6747 432 6759 1042
rect 6795 432 6807 1042
rect 6891 744 6903 1042
rect 7011 768 7023 1042
rect 7059 24 7071 1042
rect 7131 792 7143 1042
rect 7299 816 7311 1042
rect 7347 840 7359 1042
rect 7491 864 7503 1042
rect 7779 912 7791 1042
rect 8043 912 8055 1042
rect 7779 0 7791 874
rect 7803 504 7815 898
rect 8259 24 8271 1042
rect 8499 792 8511 1042
rect 8619 72 8631 1042
rect 8763 336 8775 1042
rect 8955 384 8967 1042
rect 8979 336 8991 1042
rect 9123 720 9135 1042
rect 9195 192 9207 1042
rect 9243 144 9255 1042
rect 9315 720 9327 1042
rect 9339 768 9351 1042
rect 9363 384 9375 1042
rect 9387 816 9399 1042
rect 9651 768 9663 1042
rect 9675 816 9687 1042
rect 9699 192 9711 1042
rect 9843 144 9855 1042
rect 9891 936 9903 1042
rect 9963 720 9975 1042
rect 10083 816 10095 1042
rect 10155 744 10167 1042
rect 10203 720 10215 1042
rect 10323 792 10335 1042
rect 10539 216 10551 1042
rect 10803 600 10815 1042
rect 10899 600 10911 1042
rect 11115 168 11127 1042
rect 11331 744 11343 1042
rect 11475 384 11487 1042
rect 12219 816 12231 1042
rect 12507 384 12519 1042
rect 12603 960 12615 1042
rect 12651 984 12663 1042
rect 12723 864 12735 1042
rect 12867 1008 12879 1042
rect 13251 1032 13263 1042
rect 13275 912 13287 1042
rect 13299 720 13311 1042
rect 13395 792 13407 1042
rect 13419 720 13431 1042
rect 13635 288 13647 1042
rect 13659 1008 13671 1042
rect 13803 576 13815 1042
rect 13947 24 13959 1042
rect 13971 240 13983 1042
rect 13995 576 14007 1042
rect 14019 792 14031 1042
rect 7815 0 7827 10
rect 14019 0 14031 298
rect 14091 216 14103 1042
rect 14187 816 14199 1042
rect 14235 744 14247 1042
rect 14259 816 14271 1042
rect 14283 744 14295 1042
rect 14451 912 14463 1042
rect 14499 1008 14511 1042
rect 14571 144 14583 1042
rect 14595 744 14607 1042
rect 14643 264 14655 1042
rect 14691 744 14703 1042
rect 15075 312 15087 1042
rect 15219 288 15231 1042
rect 15627 816 15639 1042
rect 15819 312 15831 1042
rect 15867 960 15879 1042
rect 16011 552 16023 1042
rect 16083 984 16095 1042
rect 16299 648 16311 1042
rect 16371 552 16383 1042
rect 16443 648 16455 1042
rect 16467 816 16479 1042
rect 16539 984 16551 1042
rect 16611 744 16623 1042
rect 16683 864 16695 1042
rect 16707 960 16719 1042
rect 16731 1032 16743 1042
rect 16827 840 16839 1042
rect 16971 528 16983 1042
rect 17019 336 17031 1042
rect 17067 528 17079 1042
rect 17163 792 17175 1042
rect 17259 696 17271 1042
rect 17355 912 17367 1042
rect 17451 696 17463 1042
rect 17499 504 17511 1042
rect 17667 936 17679 1042
rect 18243 48 18255 1042
rect 18651 288 18663 1042
rect 19011 744 19023 1042
rect 19059 600 19071 1042
rect 19107 600 19119 1042
rect 19443 192 19455 1042
rect 20067 168 20079 1042
rect 20091 768 20103 1042
rect 20259 768 20271 1042
rect 20883 504 20895 1042
rect 20907 984 20919 1042
rect 21099 456 21111 1042
rect 21195 72 21207 1042
rect 21315 96 21327 1042
rect 21411 720 21423 1042
rect 21555 960 21567 1042
rect 21675 768 21687 1042
rect 21747 816 21759 1042
rect 21867 312 21879 1042
rect 22107 480 22119 1042
rect 22227 672 22239 1042
rect 22323 408 22335 1042
rect 22419 408 22431 1042
rect 22491 672 22503 1042
rect 22539 624 22551 1042
rect 22587 120 22599 1042
rect 22755 504 22767 1042
rect 22827 576 22839 1042
rect 22875 216 22887 1042
rect 23595 576 23607 1042
rect 23643 672 23655 1042
rect 23608 562 23626 576
rect 23607 0 23619 562
rect 23667 528 23679 1042
rect 23787 696 23799 1042
rect 23931 600 23943 1042
rect 24291 648 24303 1042
rect 24483 168 24495 1042
rect 24627 744 24639 1042
rect 24843 384 24855 1042
rect 24915 408 24927 1042
rect 25227 888 25239 1042
rect 25251 1008 25263 1042
rect 25371 360 25383 1042
rect 26043 528 26055 1042
rect 26091 576 26103 1042
rect 26091 24 26103 418
rect 26115 48 26127 514
rect 26139 72 26151 562
rect 26547 0 26747 1042
rect 26835 539 26905 551
rect 26835 59 26905 71
rect 26835 35 26905 47
rect 26835 11 26905 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 123 0 1 6819
box 0 0 1464 799
use nand2 g8541
timestamp 1386234792
transform 1 0 1587 0 1 6819
box 0 0 96 799
use nor2 g8462
timestamp 1386235306
transform 1 0 1683 0 1 6819
box 0 0 120 799
use nand3 g8469
timestamp 1386234893
transform 1 0 1803 0 1 6819
box 0 0 120 799
use inv g8513
timestamp 1386238110
transform 1 0 1923 0 1 6819
box 0 0 120 799
use inv g8639
timestamp 1386238110
transform 1 0 2043 0 1 6819
box 0 0 120 799
use nor2 g8774
timestamp 1386235306
transform 1 0 2163 0 1 6819
box 0 0 120 799
use inv g8756
timestamp 1386238110
transform 1 0 2283 0 1 6819
box 0 0 120 799
use nand2 g8642
timestamp 1386234792
transform 1 0 2403 0 1 6819
box 0 0 96 799
use nand2 g8545
timestamp 1386234792
transform 1 0 2499 0 1 6819
box 0 0 96 799
use nand2 g8536
timestamp 1386234792
transform 1 0 2595 0 1 6819
box 0 0 96 799
use nand3 g8724
timestamp 1386234893
transform 1 0 2691 0 1 6819
box 0 0 120 799
use nand2 g8554
timestamp 1386234792
transform 1 0 2811 0 1 6819
box 0 0 96 799
use nand2 g8477
timestamp 1386234792
transform 1 0 2907 0 1 6819
box 0 0 96 799
use nand3 g8506
timestamp 1386234893
transform 1 0 3003 0 1 6819
box 0 0 120 799
use nand2 g8758
timestamp 1386234792
transform 1 0 3123 0 1 6819
box 0 0 96 799
use nand2 g8567
timestamp 1386234792
transform 1 0 3219 0 1 6819
box 0 0 96 799
use nand2 g8623
timestamp 1386234792
transform 1 0 3315 0 1 6819
box 0 0 96 799
use nor2 g8474
timestamp 1386235306
transform 1 0 3411 0 1 6819
box 0 0 120 799
use nand2 g8585
timestamp 1386234792
transform 1 0 3531 0 1 6819
box 0 0 96 799
use nand2 g8640
timestamp 1386234792
transform 1 0 3627 0 1 6819
box 0 0 96 799
use inv g8584
timestamp 1386238110
transform 1 0 3723 0 1 6819
box 0 0 120 799
use inv g8603
timestamp 1386238110
transform 1 0 3843 0 1 6819
box 0 0 120 799
use and2 g8597
timestamp 1386234845
transform 1 0 3963 0 1 6819
box 0 0 120 799
use nand2 g8472
timestamp 1386234792
transform 1 0 4083 0 1 6819
box 0 0 96 799
use nor2 g8712
timestamp 1386235306
transform 1 0 4179 0 1 6819
box 0 0 120 799
use mux2 g8655
timestamp 1386235218
transform 1 0 4299 0 1 6819
box 0 0 192 799
use and2 g8749
timestamp 1386234845
transform 1 0 4491 0 1 6819
box 0 0 120 799
use inv g8741
timestamp 1386238110
transform 1 0 4611 0 1 6819
box 0 0 120 799
use inv g8572
timestamp 1386238110
transform 1 0 4731 0 1 6819
box 0 0 120 799
use nand2 g8772
timestamp 1386234792
transform 1 0 4851 0 1 6819
box 0 0 96 799
use inv g8763
timestamp 1386238110
transform 1 0 4947 0 1 6819
box 0 0 120 799
use inv g8729
timestamp 1386238110
transform 1 0 5067 0 1 6819
box 0 0 120 799
use nand2 g8761
timestamp 1386234792
transform 1 0 5187 0 1 6819
box 0 0 96 799
use nand2 g8456
timestamp 1386234792
transform 1 0 5283 0 1 6819
box 0 0 96 799
use nand4 g8450
timestamp 1386234936
transform 1 0 5379 0 1 6819
box 0 0 144 799
use nand2 g8589
timestamp 1386234792
transform 1 0 5523 0 1 6819
box 0 0 96 799
use inv g8645
timestamp 1386238110
transform 1 0 5619 0 1 6819
box 0 0 120 799
use nand2 g8649
timestamp 1386234792
transform 1 0 5739 0 1 6819
box 0 0 96 799
use nand3 g8616
timestamp 1386234893
transform 1 0 5835 0 1 6819
box 0 0 120 799
use and2 g8690
timestamp 1386234845
transform 1 0 5955 0 1 6819
box 0 0 120 799
use inv g8683
timestamp 1386238110
transform 1 0 6075 0 1 6819
box 0 0 120 799
use nand2 g8667
timestamp 1386234792
transform 1 0 6195 0 1 6819
box 0 0 96 799
use nor2 g8547
timestamp 1386235306
transform 1 0 6291 0 1 6819
box 0 0 120 799
use nand2 g8493
timestamp 1386234792
transform 1 0 6411 0 1 6819
box 0 0 96 799
use nand2 g8440
timestamp 1386234792
transform 1 0 6507 0 1 6819
box 0 0 96 799
use rowcrosser AluWe
timestamp 1386086759
transform 1 0 6603 0 1 6819
box 0 0 48 799
use inv g8504
timestamp 1386238110
transform 1 0 6651 0 1 6819
box 0 0 120 799
use nand2 g8449
timestamp 1386234792
transform 1 0 6771 0 1 6819
box 0 0 96 799
use nand2 g8414
timestamp 1386234792
transform 1 0 6867 0 1 6819
box 0 0 96 799
use nand3 g8418
timestamp 1386234893
transform 1 0 6963 0 1 6819
box 0 0 120 799
use nand2 g8636
timestamp 1386234792
transform 1 0 7083 0 1 6819
box 0 0 96 799
use nand3 g8651
timestamp 1386234893
transform 1 0 7179 0 1 6819
box 0 0 120 799
use rowcrosser StatusRegEn
timestamp 1386086759
transform 1 0 7299 0 1 6819
box 0 0 48 799
use nand2 g8620
timestamp 1386234792
transform 1 0 7347 0 1 6819
box 0 0 96 799
use nand2 g8483
timestamp 1386234792
transform 1 0 7443 0 1 6819
box 0 0 96 799
use nand2 g8717
timestamp 1386234792
transform 1 0 7539 0 1 6819
box 0 0 96 799
use nand2 g8666
timestamp 1386234792
transform 1 0 7635 0 1 6819
box 0 0 96 799
use nor2 g8511
timestamp 1386235306
transform 1 0 7731 0 1 6819
box 0 0 120 799
use nand2 g8696
timestamp 1386234792
transform 1 0 7851 0 1 6819
box 0 0 96 799
use nand2 g8407
timestamp 1386234792
transform 1 0 7947 0 1 6819
box 0 0 96 799
use nand3 g8486
timestamp 1386234893
transform 1 0 8043 0 1 6819
box 0 0 120 799
use nand2 g8618
timestamp 1386234792
transform 1 0 8163 0 1 6819
box 0 0 96 799
use nand3 g8562
timestamp 1386234893
transform 1 0 8259 0 1 6819
box 0 0 120 799
use nand2 g8703
timestamp 1386234792
transform 1 0 8379 0 1 6819
box 0 0 96 799
use and2 g8489
timestamp 1386234845
transform 1 0 8475 0 1 6819
box 0 0 120 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 8595 0 1 6819
box 0 0 48 799
use nand2 g8723
timestamp 1386234792
transform 1 0 8643 0 1 6819
box 0 0 96 799
use inv g8735
timestamp 1386238110
transform 1 0 8739 0 1 6819
box 0 0 120 799
use rowcrosser ALE
timestamp 1386086759
transform 1 0 8859 0 1 6819
box 0 0 48 799
use nand2 g8403
timestamp 1386234792
transform 1 0 8907 0 1 6819
box 0 0 96 799
use nand2 g8612
timestamp 1386234792
transform 1 0 9003 0 1 6819
box 0 0 96 799
use nand2 g8631
timestamp 1386234792
transform 1 0 9099 0 1 6819
box 0 0 96 799
use inv g8532
timestamp 1386238110
transform 1 0 9195 0 1 6819
box 0 0 120 799
use nand3 g8529
timestamp 1386234893
transform 1 0 9315 0 1 6819
box 0 0 120 799
use nand3 g8676
timestamp 1386234893
transform 1 0 9435 0 1 6819
box 0 0 120 799
use nand2 g8538
timestamp 1386234792
transform 1 0 9555 0 1 6819
box 0 0 96 799
use nand2 g8580
timestamp 1386234792
transform 1 0 9651 0 1 6819
box 0 0 96 799
use nand3 g8594
timestamp 1386234893
transform 1 0 9747 0 1 6819
box 0 0 120 799
use nand2 g8648
timestamp 1386234792
transform 1 0 9867 0 1 6819
box 0 0 96 799
use nand2 g8425
timestamp 1386234792
transform 1 0 9963 0 1 6819
box 0 0 96 799
use nand3 g8524
timestamp 1386234893
transform 1 0 10059 0 1 6819
box 0 0 120 799
use nand2 g8609
timestamp 1386234792
transform 1 0 10179 0 1 6819
box 0 0 96 799
use nor2 g8743
timestamp 1386235306
transform 1 0 10275 0 1 6819
box 0 0 120 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 10395 0 1 6819
box 0 0 48 799
use nor2 g8479
timestamp 1386235306
transform 1 0 10443 0 1 6819
box 0 0 120 799
use nand2 g8728
timestamp 1386234792
transform 1 0 10563 0 1 6819
box 0 0 96 799
use nor2 g8564
timestamp 1386235306
transform 1 0 10659 0 1 6819
box 0 0 120 799
use nand2 g8699
timestamp 1386234792
transform 1 0 10779 0 1 6819
box 0 0 96 799
use and2 g8694
timestamp 1386234845
transform 1 0 10875 0 1 6819
box 0 0 120 799
use nand2 g8533
timestamp 1386234792
transform 1 0 10995 0 1 6819
box 0 0 96 799
use mux2 g8700
timestamp 1386235218
transform 1 0 11091 0 1 6819
box 0 0 192 799
use rowcrosser WdSel
timestamp 1386086759
transform 1 0 11283 0 1 6819
box 0 0 48 799
use inv g8627
timestamp 1386238110
transform 1 0 11331 0 1 6819
box 0 0 120 799
use and2 g8634
timestamp 1386234845
transform 1 0 11451 0 1 6819
box 0 0 120 799
use nand2 g8731
timestamp 1386234792
transform 1 0 11571 0 1 6819
box 0 0 96 799
use inv g8746
timestamp 1386238110
transform 1 0 11667 0 1 6819
box 0 0 120 799
use nand2 g8705
timestamp 1386234792
transform 1 0 11787 0 1 6819
box 0 0 96 799
use nand2 g8431
timestamp 1386234792
transform 1 0 11883 0 1 6819
box 0 0 96 799
use nor2 rm_assigns_buf_StatusReg_1
timestamp 1386235306
transform 1 0 11979 0 1 6819
box 0 0 120 799
use buffer g8421
timestamp 1386236986
transform 1 0 12099 0 1 6819
box 0 0 120 799
use nor2 g8399
timestamp 1386235306
transform 1 0 12219 0 1 6819
box 0 0 120 799
use nand4 g8778
timestamp 1386234936
transform 1 0 12339 0 1 6819
box 0 0 144 799
use inv g8507
timestamp 1386238110
transform 1 0 12483 0 1 6819
box 0 0 120 799
use nand2 g8688
timestamp 1386234792
transform 1 0 12603 0 1 6819
box 0 0 96 799
use nand3 g8411
timestamp 1386234893
transform 1 0 12699 0 1 6819
box 0 0 120 799
use nor2 g8553
timestamp 1386235306
transform 1 0 12819 0 1 6819
box 0 0 120 799
use inv g8646
timestamp 1386238110
transform 1 0 12939 0 1 6819
box 0 0 120 799
use rowcrosser PcEn
timestamp 1386086759
transform 1 0 13059 0 1 6819
box 0 0 48 799
use nand2 g8417
timestamp 1386234792
transform 1 0 13107 0 1 6819
box 0 0 96 799
use nand2 g8658
timestamp 1386234792
transform 1 0 13203 0 1 6819
box 0 0 96 799
use nand3 g8698
timestamp 1386234893
transform 1 0 13299 0 1 6819
box 0 0 120 799
use and2 g8641
timestamp 1386234845
transform 1 0 13419 0 1 6819
box 0 0 120 799
use nand2 StatusReg_reg_91_3_93_
timestamp 1386234792
transform 1 0 13539 0 1 6819
box 0 0 96 799
use scandtype stateSub_reg_91_2_93_
timestamp 1386241841
transform 1 0 13635 0 1 6819
box 0 0 624 799
use scandtype g8546
timestamp 1386241841
transform 1 0 14259 0 1 6819
box 0 0 624 799
use nand2 g8750
timestamp 1386234792
transform 1 0 14883 0 1 6819
box 0 0 96 799
use nand2 g8444
timestamp 1386234792
transform 1 0 14979 0 1 6819
box 0 0 96 799
use nand4 g8466
timestamp 1386234936
transform 1 0 15075 0 1 6819
box 0 0 144 799
use nand4 g8468
timestamp 1386234936
transform 1 0 15219 0 1 6819
box 0 0 144 799
use nand4 g8433
timestamp 1386234936
transform 1 0 15363 0 1 6819
box 0 0 144 799
use nand4 g8420
timestamp 1386234936
transform 1 0 15507 0 1 6819
box 0 0 144 799
use nand4 g8624
timestamp 1386234936
transform 1 0 15651 0 1 6819
box 0 0 144 799
use nand2 g8668
timestamp 1386234792
transform 1 0 15795 0 1 6819
box 0 0 96 799
use and2 g8733
timestamp 1386234845
transform 1 0 15891 0 1 6819
box 0 0 120 799
use nor2 g8537
timestamp 1386235306
transform 1 0 16011 0 1 6819
box 0 0 120 799
use nor2 g8531
timestamp 1386235306
transform 1 0 16131 0 1 6819
box 0 0 120 799
use nand3 g8542
timestamp 1386234893
transform 1 0 16251 0 1 6819
box 0 0 120 799
use nand4 g8754
timestamp 1386234936
transform 1 0 16371 0 1 6819
box 0 0 144 799
use nor2 g8760
timestamp 1386235306
transform 1 0 16515 0 1 6819
box 0 0 120 799
use nand2 StatusReg_reg_91_1_93_
timestamp 1386234792
transform 1 0 16635 0 1 6819
box 0 0 96 799
use scandtype g8435
timestamp 1386241841
transform 1 0 16731 0 1 6819
box 0 0 624 799
use rowcrosser LrWe
timestamp 1386086759
transform 1 0 17355 0 1 6819
box 0 0 48 799
use nand4 g8452
timestamp 1386234936
transform 1 0 17403 0 1 6819
box 0 0 144 799
use nand2 g8710
timestamp 1386234792
transform 1 0 17547 0 1 6819
box 0 0 96 799
use nand2 g8610
timestamp 1386234792
transform 1 0 17643 0 1 6819
box 0 0 96 799
use nand2 g8635
timestamp 1386234792
transform 1 0 17739 0 1 6819
box 0 0 96 799
use nor2 g8713
timestamp 1386235306
transform 1 0 17835 0 1 6819
box 0 0 120 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 17955 0 1 6819
box 0 0 48 799
use xor2 g8604
timestamp 1386237344
transform 1 0 18003 0 1 6819
box 0 0 192 799
use nand2 g8691
timestamp 1386234792
transform 1 0 18195 0 1 6819
box 0 0 96 799
use nand2 g8522
timestamp 1386234792
transform 1 0 18291 0 1 6819
box 0 0 96 799
use and2 g8656
timestamp 1386234845
transform 1 0 18387 0 1 6819
box 0 0 120 799
use inv g8535
timestamp 1386238110
transform 1 0 18507 0 1 6819
box 0 0 120 799
use nand3 g8516
timestamp 1386234893
transform 1 0 18627 0 1 6819
box 0 0 120 799
use nand2 g8514
timestamp 1386234792
transform 1 0 18747 0 1 6819
box 0 0 96 799
use nand2 g8673
timestamp 1386234792
transform 1 0 18843 0 1 6819
box 0 0 96 799
use nand2 g8559
timestamp 1386234792
transform 1 0 18939 0 1 6819
box 0 0 96 799
use nand2 g8748
timestamp 1386234792
transform 1 0 19035 0 1 6819
box 0 0 96 799
use nand2 g8718
timestamp 1386234792
transform 1 0 19131 0 1 6819
box 0 0 96 799
use nor2 g8590
timestamp 1386235306
transform 1 0 19227 0 1 6819
box 0 0 120 799
use nand3 g8670
timestamp 1386234893
transform 1 0 19347 0 1 6819
box 0 0 120 799
use nor2 g8619
timestamp 1386235306
transform 1 0 19467 0 1 6819
box 0 0 120 799
use nand3 g8599
timestamp 1386234893
transform 1 0 19587 0 1 6819
box 0 0 120 799
use inv g8480
timestamp 1386238110
transform 1 0 19707 0 1 6819
box 0 0 120 799
use nand2 g8436
timestamp 1386234792
transform 1 0 19827 0 1 6819
box 0 0 96 799
use nand2 g8586
timestamp 1386234792
transform 1 0 19923 0 1 6819
box 0 0 96 799
use nand2 g8548
timestamp 1386234792
transform 1 0 20019 0 1 6819
box 0 0 96 799
use nand2 g8740
timestamp 1386234792
transform 1 0 20115 0 1 6819
box 0 0 96 799
use nor2 g8653
timestamp 1386235306
transform 1 0 20211 0 1 6819
box 0 0 120 799
use nand2 g8595
timestamp 1386234792
transform 1 0 20331 0 1 6819
box 0 0 96 799
use nand2 g8720
timestamp 1386234792
transform 1 0 20427 0 1 6819
box 0 0 96 799
use nand2 g8573
timestamp 1386234792
transform 1 0 20523 0 1 6819
box 0 0 96 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 20619 0 1 6819
box 0 0 48 799
use nand2 g8701
timestamp 1386234792
transform 1 0 20667 0 1 6819
box 0 0 96 799
use nand2 g8674
timestamp 1386234792
transform 1 0 20763 0 1 6819
box 0 0 96 799
use rowcrosser Flags_91_1_93_
timestamp 1386086759
transform 1 0 20859 0 1 6819
box 0 0 48 799
use nand2 g8630
timestamp 1386234792
transform 1 0 20907 0 1 6819
box 0 0 96 799
use nand2 g8732
timestamp 1386234792
transform 1 0 21003 0 1 6819
box 0 0 96 799
use nand2 StatusReg_reg_91_0_93_
timestamp 1386234792
transform 1 0 21099 0 1 6819
box 0 0 96 799
use scandtype g8591
timestamp 1386241841
transform 1 0 21195 0 1 6819
box 0 0 624 799
use rowcrosser AluEn
timestamp 1386086759
transform 1 0 21819 0 1 6819
box 0 0 48 799
use nand3 g8702
timestamp 1386234893
transform 1 0 21867 0 1 6819
box 0 0 120 799
use nand2 g8443
timestamp 1386234792
transform 1 0 21987 0 1 6819
box 0 0 96 799
use inv g8427
timestamp 1386238110
transform 1 0 22083 0 1 6819
box 0 0 120 799
use nand3 g8432
timestamp 1386234893
transform 1 0 22203 0 1 6819
box 0 0 120 799
use nand3 g8424
timestamp 1386234893
transform 1 0 22323 0 1 6819
box 0 0 120 799
use nand4 g8410
timestamp 1386234936
transform 1 0 22443 0 1 6819
box 0 0 144 799
use rowcrosser Op2Sel_91_1_93_
timestamp 1386086759
transform 1 0 22587 0 1 6819
box 0 0 48 799
use nand4 g8503
timestamp 1386234936
transform 1 0 22635 0 1 6819
box 0 0 144 799
use nand3 g8588
timestamp 1386234893
transform 1 0 22779 0 1 6819
box 0 0 120 799
use nor2 g8495
timestamp 1386235306
transform 1 0 22899 0 1 6819
box 0 0 120 799
use nand3 g8659
timestamp 1386234893
transform 1 0 23019 0 1 6819
box 0 0 120 799
use nand2 g8406
timestamp 1386234792
transform 1 0 23139 0 1 6819
box 0 0 96 799
use nand3 g8487
timestamp 1386234893
transform 1 0 23235 0 1 6819
box 0 0 120 799
use nand3 g8508
timestamp 1386234893
transform 1 0 23355 0 1 6819
box 0 0 120 799
use nand3 g8563
timestamp 1386234893
transform 1 0 23475 0 1 6819
box 0 0 120 799
use nand2 g8677
timestamp 1386234792
transform 1 0 23595 0 1 6819
box 0 0 96 799
use inv g8706
timestamp 1386238110
transform 1 0 23691 0 1 6819
box 0 0 120 799
use nand2 g8439
timestamp 1386234792
transform 1 0 23811 0 1 6819
box 0 0 96 799
use nand2 g8473
timestamp 1386234792
transform 1 0 23907 0 1 6819
box 0 0 96 799
use nand3 g8600
timestamp 1386234893
transform 1 0 24003 0 1 6819
box 0 0 120 799
use nand2 g8695
timestamp 1386234792
transform 1 0 24123 0 1 6819
box 0 0 96 799
use nand2 g8637
timestamp 1386234792
transform 1 0 24219 0 1 6819
box 0 0 96 799
use nand2 g8494
timestamp 1386234792
transform 1 0 24315 0 1 6819
box 0 0 96 799
use nand3 g8465
timestamp 1386234893
transform 1 0 24411 0 1 6819
box 0 0 120 799
use nand4 g8523
timestamp 1386234936
transform 1 0 24531 0 1 6819
box 0 0 144 799
use nand3 g8615
timestamp 1386234893
transform 1 0 24675 0 1 6819
box 0 0 120 799
use nand4 g8455
timestamp 1386234936
transform 1 0 24795 0 1 6819
box 0 0 144 799
use nand2 g8650
timestamp 1386234792
transform 1 0 24939 0 1 6819
box 0 0 96 799
use nand2 g8478
timestamp 1386234792
transform 1 0 25035 0 1 6819
box 0 0 96 799
use and2 g8744
timestamp 1386234845
transform 1 0 25131 0 1 6819
box 0 0 120 799
use and2 g8663
timestamp 1386234845
transform 1 0 25251 0 1 6819
box 0 0 120 799
use nand3 g8447
timestamp 1386234893
transform 1 0 25371 0 1 6819
box 0 0 120 799
use nand2 g8575
timestamp 1386234792
transform 1 0 25491 0 1 6819
box 0 0 96 799
use nand2 g8759
timestamp 1386234792
transform 1 0 25587 0 1 6819
box 0 0 96 799
use nand2 g8714
timestamp 1386234792
transform 1 0 25683 0 1 6819
box 0 0 96 799
use mux2 g8540
timestamp 1386235218
transform 1 0 25779 0 1 6819
box 0 0 192 799
use and2 g8510
timestamp 1386234845
transform 1 0 25971 0 1 6819
box 0 0 120 799
use nand2 g8451
timestamp 1386234792
transform 1 0 26091 0 1 6819
box 0 0 96 799
use nand2 g8519
timestamp 1386234792
transform 1 0 26187 0 1 6819
box 0 0 96 799
use nand2 LrSel
timestamp 1386234792
transform 1 0 26283 0 1 6819
box 0 0 96 799
use rowcrosser LrEn
timestamp 1386086759
transform 1 0 26379 0 1 6819
box 0 0 48 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 26427 0 1 6819
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 123 0 1 1042
box 0 0 1464 799
use nand2 g8747
timestamp 1386234792
transform 1 0 1587 0 1 1042
box 0 0 96 799
use rowcrosser g8737
timestamp 1386086759
transform 1 0 1683 0 1 1042
box 0 0 48 799
use and2 stateSub_reg_91_0_93_
timestamp 1386234845
transform 1 0 1731 0 1 1042
box 0 0 120 799
use scandtype g8625
timestamp 1386241841
transform 1 0 1851 0 1 1042
box 0 0 624 799
use nand2 g8552
timestamp 1386234792
transform 1 0 2475 0 1 1042
box 0 0 96 799
use nor2 g8558
timestamp 1386235306
transform 1 0 2571 0 1 1042
box 0 0 120 799
use and2 g8777
timestamp 1386234845
transform 1 0 2691 0 1 1042
box 0 0 120 799
use inv g8430
timestamp 1386238110
transform 1 0 2811 0 1 1042
box 0 0 120 799
use nand3 g8697
timestamp 1386234893
transform 1 0 2931 0 1 1042
box 0 0 120 799
use nand2 g8614
timestamp 1386234792
transform 1 0 3051 0 1 1042
box 0 0 96 799
use nand2 g8629
timestamp 1386234792
transform 1 0 3147 0 1 1042
box 0 0 96 799
use nand2 g8543
timestamp 1386234792
transform 1 0 3243 0 1 1042
box 0 0 96 799
use nand2 state_reg_91_1_93_
timestamp 1386234792
transform 1 0 3339 0 1 1042
box 0 0 96 799
use scandtype g8416
timestamp 1386241841
transform 1 0 3435 0 1 1042
box 0 0 624 799
use nand2 g8434
timestamp 1386234792
transform 1 0 4059 0 1 1042
box 0 0 96 799
use and2 g8578
timestamp 1386234845
transform 1 0 4155 0 1 1042
box 0 0 120 799
use nand3 g8556
timestamp 1386234893
transform 1 0 4275 0 1 1042
box 0 0 120 799
use nand2 g8566
timestamp 1386234792
transform 1 0 4395 0 1 1042
box 0 0 96 799
use nand2 g8611
timestamp 1386234792
transform 1 0 4491 0 1 1042
box 0 0 96 799
use nand2 g8429
timestamp 1386234792
transform 1 0 4587 0 1 1042
box 0 0 96 799
use nand4 g8726
timestamp 1386234936
transform 1 0 4683 0 1 1042
box 0 0 144 799
use nand2 g8458
timestamp 1386234792
transform 1 0 4827 0 1 1042
box 0 0 96 799
use nand2 g8736
timestamp 1386234792
transform 1 0 4923 0 1 1042
box 0 0 96 799
use inv g8476
timestamp 1386238110
transform 1 0 5019 0 1 1042
box 0 0 120 799
use nor2 g8687
timestamp 1386235306
transform 1 0 5139 0 1 1042
box 0 0 120 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 5259 0 1 1042
box 0 0 96 799
use scandtype g8498
timestamp 1386241841
transform 1 0 5355 0 1 1042
box 0 0 624 799
use rowcrosser SysBus_91_3_93_
timestamp 1386086759
transform 1 0 5979 0 1 1042
box 0 0 48 799
use nand4 g8501
timestamp 1386234936
transform 1 0 6027 0 1 1042
box 0 0 144 799
use nor2 g8587
timestamp 1386235306
transform 1 0 6171 0 1 1042
box 0 0 120 799
use nand2 g8608
timestamp 1386234792
transform 1 0 6291 0 1 1042
box 0 0 96 799
use nand2 g8534
timestamp 1386234792
transform 1 0 6387 0 1 1042
box 0 0 96 799
use nand2 g8454
timestamp 1386234792
transform 1 0 6483 0 1 1042
box 0 0 96 799
use nand2 g8442
timestamp 1386234792
transform 1 0 6579 0 1 1042
box 0 0 96 799
use nand4 g8680
timestamp 1386234936
transform 1 0 6675 0 1 1042
box 0 0 144 799
use nand2 g8521
timestamp 1386234792
transform 1 0 6819 0 1 1042
box 0 0 96 799
use nand3 g8394
timestamp 1386234893
transform 1 0 6915 0 1 1042
box 0 0 120 799
use rowcrosser AluOR_91_1_93_
timestamp 1386086759
transform 1 0 7035 0 1 1042
box 0 0 48 799
use nand4 g8692
timestamp 1386234936
transform 1 0 7083 0 1 1042
box 0 0 144 799
use nand2 g8453
timestamp 1386234792
transform 1 0 7227 0 1 1042
box 0 0 96 799
use nand2 g8719
timestamp 1386234792
transform 1 0 7323 0 1 1042
box 0 0 96 799
use nand2 g8644
timestamp 1386234792
transform 1 0 7419 0 1 1042
box 0 0 96 799
use nand2 g8461
timestamp 1386234792
transform 1 0 7515 0 1 1042
box 0 0 96 799
use inv g8679
timestamp 1386238110
transform 1 0 7611 0 1 1042
box 0 0 120 799
use nand2 g8770
timestamp 1386234792
transform 1 0 7731 0 1 1042
box 0 0 96 799
use inv g8661
timestamp 1386238110
transform 1 0 7827 0 1 1042
box 0 0 120 799
use nand3 g8776
timestamp 1386234893
transform 1 0 7947 0 1 1042
box 0 0 120 799
use inv g8550
timestamp 1386238110
transform 1 0 8067 0 1 1042
box 0 0 120 799
use nand2 g8438
timestamp 1386234792
transform 1 0 8187 0 1 1042
box 0 0 96 799
use nand2 g8549
timestamp 1386234792
transform 1 0 8283 0 1 1042
box 0 0 96 799
use nand2 g8412
timestamp 1386234792
transform 1 0 8379 0 1 1042
box 0 0 96 799
use nand3 g8481
timestamp 1386234893
transform 1 0 8475 0 1 1042
box 0 0 120 799
use inv g8457
timestamp 1386238110
transform 1 0 8595 0 1 1042
box 0 0 120 799
use nand2 g8518
timestamp 1386234792
transform 1 0 8715 0 1 1042
box 0 0 96 799
use nand2 g8515
timestamp 1386234792
transform 1 0 8811 0 1 1042
box 0 0 96 799
use nand2 g8484
timestamp 1386234792
transform 1 0 8907 0 1 1042
box 0 0 96 799
use nand4 g8496
timestamp 1386234936
transform 1 0 9003 0 1 1042
box 0 0 144 799
use nand4 g8470
timestamp 1386234936
transform 1 0 9147 0 1 1042
box 0 0 144 799
use nand4 g8707
timestamp 1386234936
transform 1 0 9291 0 1 1042
box 0 0 144 799
use nand2 g8574
timestamp 1386234792
transform 1 0 9435 0 1 1042
box 0 0 96 799
use nand2 g8426
timestamp 1386234792
transform 1 0 9531 0 1 1042
box 0 0 96 799
use nand4 g8660
timestamp 1386234936
transform 1 0 9627 0 1 1042
box 0 0 144 799
use nand2 g8579
timestamp 1386234792
transform 1 0 9771 0 1 1042
box 0 0 96 799
use nand3 g8509
timestamp 1386234893
transform 1 0 9867 0 1 1042
box 0 0 120 799
use nand3 g8592
timestamp 1386234893
transform 1 0 9987 0 1 1042
box 0 0 120 799
use and2 g8490
timestamp 1386234845
transform 1 0 10107 0 1 1042
box 0 0 120 799
use and2 g8500
timestamp 1386234845
transform 1 0 10227 0 1 1042
box 0 0 120 799
use nor2 g8605
timestamp 1386235306
transform 1 0 10347 0 1 1042
box 0 0 120 799
use inv g8446
timestamp 1386238110
transform 1 0 10467 0 1 1042
box 0 0 120 799
use and2 g8560
timestamp 1386234845
transform 1 0 10587 0 1 1042
box 0 0 120 799
use nand3 g8459
timestamp 1386234893
transform 1 0 10707 0 1 1042
box 0 0 120 799
use nand2 g8753
timestamp 1386234792
transform 1 0 10827 0 1 1042
box 0 0 96 799
use nand2 g8684
timestamp 1386234792
transform 1 0 10923 0 1 1042
box 0 0 96 799
use and2 g8638
timestamp 1386234845
transform 1 0 11019 0 1 1042
box 0 0 120 799
use inv g8527
timestamp 1386238110
transform 1 0 11139 0 1 1042
box 0 0 120 799
use nand2 g8570
timestamp 1386234792
transform 1 0 11259 0 1 1042
box 0 0 96 799
use nand4 g8530
timestamp 1386234936
transform 1 0 11355 0 1 1042
box 0 0 144 799
use nand3 IntStatus_reg
timestamp 1386234893
transform 1 0 11499 0 1 1042
box 0 0 120 799
use scanreg g8745
timestamp 1386241447
transform 1 0 11619 0 1 1042
box 0 0 720 799
use and2 g8491
timestamp 1386234845
transform 1 0 12339 0 1 1042
box 0 0 120 799
use and2 g8721
timestamp 1386234845
transform 1 0 12459 0 1 1042
box 0 0 120 799
use inv g8715
timestamp 1386238110
transform 1 0 12579 0 1 1042
box 0 0 120 799
use nand2 g8437
timestamp 1386234792
transform 1 0 12699 0 1 1042
box 0 0 96 799
use nand2 g8755
timestamp 1386234792
transform 1 0 12795 0 1 1042
box 0 0 96 799
use inv g8752
timestamp 1386238110
transform 1 0 12891 0 1 1042
box 0 0 120 799
use nor2 g8678
timestamp 1386235306
transform 1 0 13011 0 1 1042
box 0 0 120 799
use nand2 g8526
timestamp 1386234792
transform 1 0 13131 0 1 1042
box 0 0 96 799
use nand4 g8423
timestamp 1386234936
transform 1 0 13227 0 1 1042
box 0 0 144 799
use nand3 g8601
timestamp 1386234893
transform 1 0 13371 0 1 1042
box 0 0 120 799
use and2 g8405
timestamp 1386234845
transform 1 0 13491 0 1 1042
box 0 0 120 799
use nand3 g8582
timestamp 1386234893
transform 1 0 13611 0 1 1042
box 0 0 120 799
use nand2 g8632
timestamp 1386234792
transform 1 0 13731 0 1 1042
box 0 0 96 799
use nand2 g8464
timestamp 1386234792
transform 1 0 13827 0 1 1042
box 0 0 96 799
use nand4 g8568
timestamp 1386234936
transform 1 0 13923 0 1 1042
box 0 0 144 799
use nand2 g8460
timestamp 1386234792
transform 1 0 14067 0 1 1042
box 0 0 96 799
use nand4 g8626
timestamp 1386234936
transform 1 0 14163 0 1 1042
box 0 0 144 799
use and2 g8404
timestamp 1386234845
transform 1 0 14307 0 1 1042
box 0 0 120 799
use nand3 g8428
timestamp 1386234893
transform 1 0 14427 0 1 1042
box 0 0 120 799
use nand3 g8413
timestamp 1386234893
transform 1 0 14547 0 1 1042
box 0 0 120 799
use nor2 g8577
timestamp 1386235306
transform 1 0 14667 0 1 1042
box 0 0 120 799
use nand3 g8682
timestamp 1386234893
transform 1 0 14787 0 1 1042
box 0 0 120 799
use and2 g8571
timestamp 1386234845
transform 1 0 14907 0 1 1042
box 0 0 120 799
use nand2 IRQ2_reg
timestamp 1386234792
transform 1 0 15027 0 1 1042
box 0 0 96 799
use scandtype g8602
timestamp 1386241841
transform 1 0 15123 0 1 1042
box 0 0 624 799
use nand2 g8669
timestamp 1386234792
transform 1 0 15747 0 1 1042
box 0 0 96 799
use nand2 g8593
timestamp 1386234792
transform 1 0 15843 0 1 1042
box 0 0 96 799
use nand2 g8686
timestamp 1386234792
transform 1 0 15939 0 1 1042
box 0 0 96 799
use nand2 g8517
timestamp 1386234792
transform 1 0 16035 0 1 1042
box 0 0 96 799
use inv g8402
timestamp 1386238110
transform 1 0 16131 0 1 1042
box 0 0 120 799
use nand4 g8738
timestamp 1386234936
transform 1 0 16251 0 1 1042
box 0 0 144 799
use nand2 g8422
timestamp 1386234792
transform 1 0 16395 0 1 1042
box 0 0 96 799
use nand4 g8622
timestamp 1386234936
transform 1 0 16491 0 1 1042
box 0 0 144 799
use nand3 g8633
timestamp 1386234893
transform 1 0 16635 0 1 1042
box 0 0 120 799
use nand2 g8488
timestamp 1386234792
transform 1 0 16755 0 1 1042
box 0 0 96 799
use nand4 g8475
timestamp 1386234936
transform 1 0 16851 0 1 1042
box 0 0 144 799
use nand2 g8598
timestamp 1386234792
transform 1 0 16995 0 1 1042
box 0 0 96 799
use nand2 g8555
timestamp 1386234792
transform 1 0 17091 0 1 1042
box 0 0 96 799
use nand2 g8415
timestamp 1386234792
transform 1 0 17187 0 1 1042
box 0 0 96 799
use nand2 g8675
timestamp 1386234792
transform 1 0 17283 0 1 1042
box 0 0 96 799
use nand2 g8725
timestamp 1386234792
transform 1 0 17379 0 1 1042
box 0 0 96 799
use inv g8643
timestamp 1386238110
transform 1 0 17475 0 1 1042
box 0 0 120 799
use inv g8742
timestamp 1386238110
transform 1 0 17595 0 1 1042
box 0 0 120 799
use nand2 g8520
timestamp 1386234792
transform 1 0 17715 0 1 1042
box 0 0 96 799
use nand2 g8708
timestamp 1386234792
transform 1 0 17811 0 1 1042
box 0 0 96 799
use and2 g8617
timestamp 1386234845
transform 1 0 17907 0 1 1042
box 0 0 120 799
use nand3 IRQ1_reg
timestamp 1386234893
transform 1 0 18027 0 1 1042
box 0 0 120 799
use scandtype g8502
timestamp 1386241841
transform 1 0 18147 0 1 1042
box 0 0 624 799
use nand3 g8505
timestamp 1386234893
transform 1 0 18771 0 1 1042
box 0 0 120 799
use nand2 g8419
timestamp 1386234792
transform 1 0 18891 0 1 1042
box 0 0 96 799
use nand4 g8596
timestamp 1386234936
transform 1 0 18987 0 1 1042
box 0 0 144 799
use and2 g8773
timestamp 1386234845
transform 1 0 19131 0 1 1042
box 0 0 120 799
use inv g8463
timestamp 1386238110
transform 1 0 19251 0 1 1042
box 0 0 120 799
use inv g8557
timestamp 1386238110
transform 1 0 19371 0 1 1042
box 0 0 120 799
use nand2 g8757
timestamp 1386234792
transform 1 0 19491 0 1 1042
box 0 0 96 799
use inv g8607
timestamp 1386238110
transform 1 0 19587 0 1 1042
box 0 0 120 799
use nand2 g8727
timestamp 1386234792
transform 1 0 19707 0 1 1042
box 0 0 96 799
use nor2 g8471
timestamp 1386235306
transform 1 0 19803 0 1 1042
box 0 0 120 799
use nand2 g8492
timestamp 1386234792
transform 1 0 19923 0 1 1042
box 0 0 96 799
use nand2 g8583
timestamp 1386234792
transform 1 0 20019 0 1 1042
box 0 0 96 799
use nand2 g8665
timestamp 1386234792
transform 1 0 20115 0 1 1042
box 0 0 96 799
use nor2 g8685
timestamp 1386235306
transform 1 0 20211 0 1 1042
box 0 0 120 799
use and2 g8662
timestamp 1386234845
transform 1 0 20331 0 1 1042
box 0 0 120 799
use inv g8621
timestamp 1386238110
transform 1 0 20451 0 1 1042
box 0 0 120 799
use nor2 g8628
timestamp 1386235306
transform 1 0 20571 0 1 1042
box 0 0 120 799
use and2 g8681
timestamp 1386234845
transform 1 0 20691 0 1 1042
box 0 0 120 799
use nand3 g8657
timestamp 1386234893
transform 1 0 20811 0 1 1042
box 0 0 120 799
use nand2 g8672
timestamp 1386234792
transform 1 0 20931 0 1 1042
box 0 0 96 799
use nand2 g8482
timestamp 1386234792
transform 1 0 21027 0 1 1042
box 0 0 96 799
use nand2 g8711
timestamp 1386234792
transform 1 0 21123 0 1 1042
box 0 0 96 799
use nand3 g8467
timestamp 1386234893
transform 1 0 21219 0 1 1042
box 0 0 120 799
use inv g8722
timestamp 1386238110
transform 1 0 21339 0 1 1042
box 0 0 120 799
use nor2 g8730
timestamp 1386235306
transform 1 0 21459 0 1 1042
box 0 0 120 799
use nor2 g8647
timestamp 1386235306
transform 1 0 21579 0 1 1042
box 0 0 120 799
use and2 g8539
timestamp 1386234845
transform 1 0 21699 0 1 1042
box 0 0 120 799
use nor2 g8565
timestamp 1386235306
transform 1 0 21819 0 1 1042
box 0 0 120 799
use and2 g8551
timestamp 1386234845
transform 1 0 21939 0 1 1042
box 0 0 120 799
use nand2 g8704
timestamp 1386234792
transform 1 0 22059 0 1 1042
box 0 0 96 799
use nand2 g8613
timestamp 1386234792
transform 1 0 22155 0 1 1042
box 0 0 96 799
use inv g8485
timestamp 1386238110
transform 1 0 22251 0 1 1042
box 0 0 120 799
use nand4 g8497
timestamp 1386234936
transform 1 0 22371 0 1 1042
box 0 0 144 799
use inv g8751
timestamp 1386238110
transform 1 0 22515 0 1 1042
box 0 0 120 799
use nand2 g8544
timestamp 1386234792
transform 1 0 22635 0 1 1042
box 0 0 96 799
use nand3 g8569
timestamp 1386234893
transform 1 0 22731 0 1 1042
box 0 0 120 799
use nand2 state_reg_91_0_93_
timestamp 1386234792
transform 1 0 22851 0 1 1042
box 0 0 96 799
use scandtype g8441
timestamp 1386241841
transform 1 0 22947 0 1 1042
box 0 0 624 799
use rowcrosser AluOR_91_0_93_
timestamp 1386086759
transform 1 0 23571 0 1 1042
box 0 0 48 799
use nand3 g8654
timestamp 1386234893
transform 1 0 23619 0 1 1042
box 0 0 120 799
use nand2 stateSub_reg_91_1_93_
timestamp 1386234792
transform 1 0 23739 0 1 1042
box 0 0 96 799
use scandtype g8652
timestamp 1386241841
transform 1 0 23835 0 1 1042
box 0 0 624 799
use nand2 g8693
timestamp 1386234792
transform 1 0 24459 0 1 1042
box 0 0 96 799
use nand2 g8767
timestamp 1386234792
transform 1 0 24555 0 1 1042
box 0 0 96 799
use inv g8525
timestamp 1386238110
transform 1 0 24651 0 1 1042
box 0 0 120 799
use nand2 g8561
timestamp 1386234792
transform 1 0 24771 0 1 1042
box 0 0 96 799
use nand2 g8528
timestamp 1386234792
transform 1 0 24867 0 1 1042
box 0 0 96 799
use nand2 g8689
timestamp 1386234792
transform 1 0 24963 0 1 1042
box 0 0 96 799
use and2 g8448
timestamp 1386234845
transform 1 0 25059 0 1 1042
box 0 0 120 799
use nand2 g8739
timestamp 1386234792
transform 1 0 25179 0 1 1042
box 0 0 96 799
use nor2 g8671
timestamp 1386235306
transform 1 0 25275 0 1 1042
box 0 0 120 799
use nand2 g8606
timestamp 1386234792
transform 1 0 25395 0 1 1042
box 0 0 96 799
use nand2 g8581
timestamp 1386234792
transform 1 0 25491 0 1 1042
box 0 0 96 799
use nand3 g8576
timestamp 1386234893
transform 1 0 25587 0 1 1042
box 0 0 120 799
use nand2 g8709
timestamp 1386234792
transform 1 0 25707 0 1 1042
box 0 0 96 799
use nand2 g8734
timestamp 1386234792
transform 1 0 25803 0 1 1042
box 0 0 96 799
use inv SysBus_91_1_93_
timestamp 1386238110
transform 1 0 25899 0 1 1042
box 0 0 120 799
use rowcrosser SysBus_91_2_93_
timestamp 1386086759
transform 1 0 26019 0 1 1042
box 0 0 48 799
use rowcrosser nWE
timestamp 1386086759
transform 1 0 26067 0 1 1042
box 0 0 48 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 26427 0 1 1042
box 0 0 320 799
<< labels >>
rlabel m2contact 26145 569 26145 569 8 AluOR[0]
rlabel m2contact 26145 65 26145 65 8 AluOR[0]
rlabel m2contact 26121 521 26121 521 8 AluOR[1]
rlabel m2contact 26121 41 26121 41 8 AluOR[1]
rlabel m2contact 26097 425 26097 425 8 ENB
rlabel m2contact 26097 17 26097 17 8 ENB
rlabel m2contact 26097 569 26097 569 8 AluOR[0]
rlabel m2contact 26049 521 26049 521 8 AluOR[1]
rlabel m2contact 25377 353 25377 353 8 n_11
rlabel m2contact 25257 1001 25257 1001 6 n_353
rlabel m2contact 25233 881 25233 881 6 SysBus[0]
rlabel m2contact 24921 401 24921 401 8 n_232
rlabel m2contact 24849 377 24849 377 8 n_129
rlabel m2contact 24633 737 24633 737 8 n_61
rlabel m2contact 24489 161 24489 161 8 n_106
rlabel m2contact 24297 641 24297 641 8 n_486
rlabel m2contact 23937 593 23937 593 8 n_337
rlabel m2contact 23793 689 23793 689 8 n_37
rlabel m2contact 23673 521 23673 521 8 n_316
rlabel m2contact 23649 665 23649 665 8 n_258
rlabel metal2 23619 569 23619 569 8 SysBus[3]
rlabel m2contact 23601 569 23601 569 8 SysBus[3]
rlabel m2contact 22881 209 22881 209 8 n_230
rlabel m2contact 22833 569 22833 569 8 n_181
rlabel m2contact 22761 497 22761 497 8 n_63
rlabel m2contact 22593 113 22593 113 8 n_291
rlabel m2contact 22545 617 22545 617 8 n_279
rlabel m2contact 22497 665 22497 665 8 n_258
rlabel m2contact 22425 401 22425 401 8 n_232
rlabel m2contact 22329 401 22329 401 8 n_232
rlabel m2contact 22233 665 22233 665 8 n_24
rlabel m2contact 22113 473 22113 473 8 n_123
rlabel m2contact 21873 305 21873 305 8 n_228
rlabel m2contact 21753 809 21753 809 6 n_16
rlabel m2contact 21681 761 21681 761 8 n_7
rlabel m2contact 21561 953 21561 953 6 n_46
rlabel m2contact 21417 713 21417 713 8 n_320
rlabel m2contact 21321 89 21321 89 8 n_18
rlabel m2contact 21201 65 21201 65 8 n_330
rlabel m2contact 21105 449 21105 449 8 n_21
rlabel m2contact 20913 977 20913 977 6 n_64
rlabel m2contact 20889 497 20889 497 8 n_63
rlabel m2contact 20265 761 20265 761 8 n_7
rlabel m2contact 20097 761 20097 761 8 n_309
rlabel m2contact 20073 161 20073 161 8 n_106
rlabel m2contact 19449 185 19449 185 8 n_306
rlabel m2contact 19113 593 19113 593 8 n_337
rlabel m2contact 19065 593 19065 593 8 n_287
rlabel m2contact 19017 737 19017 737 8 n_61
rlabel m2contact 18657 281 18657 281 8 IRQ1
rlabel m2contact 18249 41 18249 41 8 n_4
rlabel m2contact 17673 929 17673 929 6 n_132
rlabel m2contact 17505 497 17505 497 8 n_63
rlabel m2contact 17457 689 17457 689 8 n_37
rlabel m2contact 17361 905 17361 905 6 n_297
rlabel m2contact 17265 689 17265 689 8 n_259
rlabel m2contact 17169 785 17169 785 8 n_154
rlabel m2contact 17073 521 17073 521 8 n_316
rlabel m2contact 17025 329 17025 329 8 n_270
rlabel m2contact 16977 521 16977 521 8 n_225
rlabel m2contact 16833 833 16833 833 6 n_118
rlabel m2contact 16737 1025 16737 1025 6 n_71
rlabel m2contact 16713 953 16713 953 6 n_46
rlabel m2contact 16689 857 16689 857 6 n_56
rlabel m2contact 16617 737 16617 737 8 n_245
rlabel m2contact 16545 977 16545 977 6 n_64
rlabel m2contact 16473 809 16473 809 6 n_16
rlabel m2contact 16449 641 16449 641 8 n_486
rlabel m2contact 16377 545 16377 545 8 RegWe
rlabel m2contact 16305 641 16305 641 8 n_278
rlabel m2contact 16089 977 16089 977 6 n_29
rlabel m2contact 16017 545 16017 545 8 n_157
rlabel m2contact 15873 953 15873 953 6 n_46
rlabel m2contact 15825 305 15825 305 8 n_228
rlabel m2contact 15633 809 15633 809 6 IRQ2
rlabel m2contact 15225 281 15225 281 8 IRQ1
rlabel m2contact 15081 305 15081 305 8 n_228
rlabel m2contact 14697 737 14697 737 8 n_245
rlabel m2contact 14649 257 14649 257 8 n_265
rlabel m2contact 14601 737 14601 737 8 n_187
rlabel m2contact 14577 137 14577 137 8 n_102
rlabel m2contact 14505 1001 14505 1001 6 n_353
rlabel m2contact 14457 905 14457 905 6 n_297
rlabel m2contact 14289 737 14289 737 8 n_187
rlabel m2contact 14265 809 14265 809 6 IRQ2
rlabel m2contact 14241 737 14241 737 8 n_128
rlabel m2contact 14193 809 14193 809 6 IntStatus
rlabel m2contact 14097 209 14097 209 8 n_230
rlabel m2contact 14025 785 14025 785 8 n_154
rlabel m2contact 14025 305 14025 305 8 SysBus[2]
rlabel m2contact 14001 569 14001 569 8 n_181
rlabel m2contact 13977 233 13977 233 8 n_240
rlabel m2contact 13953 17 13953 17 8 n_236
rlabel m2contact 13809 569 13809 569 8 n_112
rlabel m2contact 13665 1001 13665 1001 4 n_328
rlabel m2contact 13641 281 13641 281 2 n_295
rlabel m2contact 13425 713 13425 713 2 n_320
rlabel m2contact 13401 785 13401 785 2 n_365
rlabel m2contact 13305 713 13305 713 2 n_125
rlabel m2contact 13281 905 13281 905 4 n_67
rlabel m2contact 13257 1025 13257 1025 4 n_71
rlabel m2contact 12873 1001 12873 1001 4 n_328
rlabel m2contact 12729 857 12729 857 4 n_56
rlabel m2contact 12657 977 12657 977 4 n_29
rlabel m2contact 12609 953 12609 953 4 n_46
rlabel m2contact 12513 377 12513 377 2 n_129
rlabel m2contact 12225 809 12225 809 4 IntStatus
rlabel m2contact 11481 377 11481 377 2 n_138
rlabel m2contact 11337 737 11337 737 2 n_128
rlabel m2contact 11121 161 11121 161 2 n_106
rlabel m2contact 10905 593 10905 593 2 n_287
rlabel m2contact 10809 593 10809 593 2 n_179
rlabel m2contact 10545 209 10545 209 2 n_230
rlabel m2contact 10329 785 10329 785 2 n_365
rlabel m2contact 10209 713 10209 713 2 n_125
rlabel m2contact 10161 737 10161 737 2 n_36
rlabel m2contact 10089 809 10089 809 4 n_192
rlabel m2contact 9969 713 9969 713 2 n_173
rlabel m2contact 9897 929 9897 929 4 n_132
rlabel m2contact 9849 137 9849 137 2 n_102
rlabel m2contact 9705 185 9705 185 2 n_306
rlabel m2contact 9681 809 9681 809 4 n_192
rlabel m2contact 9657 761 9657 761 2 n_309
rlabel m2contact 9393 809 9393 809 4 n_87
rlabel m2contact 9369 377 9369 377 2 n_138
rlabel m2contact 9345 761 9345 761 2 n_218
rlabel m2contact 9321 713 9321 713 2 n_173
rlabel m2contact 9249 137 9249 137 2 n_82
rlabel m2contact 9201 185 9201 185 2 n_107
rlabel m2contact 9129 713 9129 713 2 n_300
rlabel m2contact 8985 329 8985 329 2 n_270
rlabel m2contact 8961 377 8961 377 2 n_204
rlabel m2contact 8769 329 8769 329 2 n_161
rlabel m2contact 8625 65 8625 65 2 n_330
rlabel m2contact 8505 785 8505 785 2 n_365
rlabel m2contact 8265 17 8265 17 2 n_236
rlabel m2contact 8049 905 8049 905 4 n_67
rlabel m2contact 7821 17 7821 17 2 SysBus[1]
rlabel m2contact 7809 905 7809 905 4 n_63
rlabel m2contact 7809 497 7809 497 2 n_63
rlabel m2contact 7785 905 7785 905 4 n_63
rlabel m2contact 7785 881 7785 881 4 SysBus[0]
rlabel m2contact 7497 857 7497 857 4 n_56
rlabel m2contact 7353 833 7353 833 4 n_118
rlabel m2contact 7305 809 7305 809 4 n_87
rlabel m2contact 7137 785 7137 785 2 n_365
rlabel m2contact 7065 17 7065 17 2 SysBus[1]
rlabel m2contact 7017 761 7017 761 2 n_218
rlabel m2contact 6897 737 6897 737 2 n_36
rlabel m2contact 6801 425 6801 425 2 ENB
rlabel m2contact 6753 425 6753 425 2 n_219
rlabel m2contact 6729 713 6729 713 2 n_300
rlabel m2contact 6633 689 6633 689 2 n_259
rlabel m2contact 6609 65 6609 65 2 n_330
rlabel m2contact 6561 65 6561 65 2 n_144
rlabel m2contact 6537 665 6537 665 2 n_24
rlabel m2contact 6513 569 6513 569 2 n_112
rlabel m2contact 6465 569 6465 569 2 n_166
rlabel m2contact 6273 641 6273 641 2 n_278
rlabel m2contact 6153 617 6153 617 2 n_279
rlabel m2contact 6129 593 6129 593 2 n_179
rlabel m2contact 6081 569 6081 569 2 n_166
rlabel m2contact 6009 305 6009 305 2 SysBus[2]
rlabel m2contact 5001 305 5001 305 2 n_274
rlabel m2contact 4977 545 4977 545 2 n_157
rlabel m2contact 4953 521 4953 521 2 n_225
rlabel m2contact 4905 497 4905 497 2 n_63
rlabel m2contact 4665 473 4665 473 2 n_123
rlabel m2contact 4641 449 4641 449 2 n_21
rlabel m2contact 4569 425 4569 425 2 n_219
rlabel m2contact 4545 401 4545 401 2 n_232
rlabel m2contact 4473 377 4473 377 2 n_204
rlabel m2contact 4449 353 4449 353 2 n_11
rlabel m2contact 4377 329 4377 329 2 n_161
rlabel m2contact 4185 305 4185 305 2 n_274
rlabel m2contact 4137 281 4137 281 2 n_295
rlabel m2contact 3537 257 3537 257 2 n_265
rlabel m2contact 3417 233 3417 233 2 n_240
rlabel m2contact 3369 209 3369 209 2 n_230
rlabel m2contact 3321 185 3321 185 2 n_107
rlabel m2contact 3273 161 3273 161 2 n_106
rlabel m2contact 3129 137 3129 137 2 n_82
rlabel m2contact 2985 113 2985 113 2 n_291
rlabel m2contact 2889 41 2889 41 2 n_4
rlabel m2contact 2841 41 2841 41 2 nIRQ
rlabel m2contact 2505 89 2505 89 2 n_18
rlabel m2contact 1953 65 1953 65 2 n_144
rlabel m2contact 1713 65 1713 65 2 nWE
rlabel m2contact 26505 7875 26505 7875 6 Flags[0]
rlabel m2contact 26505 7635 26505 7635 6 Flags[0]
rlabel m2contact 26481 7707 26481 7707 6 Flags[3]
rlabel m2contact 26481 7635 26481 7635 6 Flags[3]
rlabel m2contact 26457 7779 26457 7779 6 Flags[2]
rlabel m2contact 26457 7683 26457 7683 6 Flags[2]
rlabel m2contact 26433 7803 26433 7803 6 CFlag
rlabel m2contact 26433 7731 26433 7731 6 CFlag
rlabel m2contact 26433 7683 26433 7683 6 Flags[1]
rlabel m2contact 26433 7659 26433 7659 6 Flags[1]
rlabel m2contact 26409 7779 26409 7779 6 Flags[2]
rlabel m2contact 25737 7779 25737 7779 6 OpcodeCondIn[0]
rlabel m2contact 25569 7755 25569 7755 6 MemEn
rlabel m2contact 25437 7707 25437 7707 6 StatusRegEn
rlabel m2contact 25017 7659 25017 7659 6 PcSel[0]
rlabel m2contact 24621 7731 24621 7731 6 StatusReg[3]
rlabel m2contact 23961 7635 23961 7635 6 Flags[3]
rlabel m2contact 23805 7947 23805 7947 6 StatusReg[2]
rlabel m2contact 23121 7851 23121 7851 6 Op2Sel[0]
rlabel m2contact 22989 7923 22989 7923 6 StatusReg[1]
rlabel m2contact 22617 7707 22617 7707 6 StatusRegEn
rlabel m2contact 22425 7635 22425 7635 6 PcSel[1]
rlabel m2contact 22173 7707 22173 7707 6 StatusReg[0]
rlabel m2contact 21849 7899 21849 7899 6 AluWe
rlabel m2contact 21705 7707 21705 7707 6 StatusReg[0]
rlabel m2contact 21357 7827 21357 7827 6 AluEn
rlabel m2contact 21333 7899 21333 7899 6 AluWe
rlabel m2contact 20889 7707 20889 7707 6 IrWe
rlabel m2contact 20649 7899 20649 7899 6 Op2Sel[1]
rlabel m2contact 20553 7731 20553 7731 6 StatusReg[3]
rlabel m2contact 20517 7899 20517 7899 6 Op2Sel[1]
rlabel m2contact 19977 7875 19977 7875 6 Flags[0]
rlabel m2contact 19701 7851 19701 7851 6 Op2Sel[0]
rlabel m2contact 19281 7779 19281 7779 6 OpcodeCondIn[0]
rlabel m2contact 18093 7851 18093 7851 6 Op1Sel
rlabel metal2 18003 7875 18003 7875 6 PcEn
rlabel m2contact 17985 7875 17985 7875 6 PcEn
rlabel m2contact 17385 7875 17385 7875 6 WdSel
rlabel m2contact 17253 7875 17253 7875 6 WdSel
rlabel m2contact 17241 7803 17241 7803 6 CFlag
rlabel m2contact 15645 7899 15645 7899 6 PcWe
rlabel m2contact 15633 7803 15633 7803 6 nME
rlabel m2contact 14829 7875 14829 7875 6 PcSel[2]
rlabel m2contact 14805 7635 14805 7635 6 PcSel[1]
rlabel m2contact 14145 7731 14145 7731 6 StatusReg[3]
rlabel m2contact 13989 7659 13989 7659 6 PcSel[0]
rlabel m2contact 13257 7947 13257 7947 4 StatusReg[2]
rlabel m2contact 13089 7683 13089 7683 4 Flags[1]
rlabel m2contact 12873 7875 12873 7875 4 PcSel[2]
rlabel m2contact 12777 7779 12777 7779 4 OpcodeCondIn[0]
rlabel m2contact 12369 7875 12369 7875 4 LrEn
rlabel m2contact 12177 7923 12177 7923 4 StatusReg[1]
rlabel m2contact 12033 7851 12033 7851 4 Op1Sel
rlabel m2contact 11541 7851 11541 7851 4 LrWe
rlabel metal2 11331 7923 11331 7923 4 LrSel
rlabel m2contact 11313 7923 11313 7923 4 LrSel
rlabel metal2 10443 7923 10443 7923 4 ImmSel
rlabel m2contact 10425 7923 10425 7923 4 ImmSel
rlabel m2contact 9849 7707 9849 7707 4 IrWe
rlabel m2contact 9081 7899 9081 7899 4 PcWe
rlabel m2contact 9021 7755 9021 7755 4 MemEn
rlabel m2contact 8961 7755 8961 7755 4 OpcodeCondIn[5]
rlabel m2contact 8889 7875 8889 7875 4 LrEn
rlabel m2contact 8625 7827 8625 7827 4 AluEn
rlabel m2contact 7401 7875 7401 7875 4 OpcodeCondIn[7]
rlabel m2contact 7329 7827 7329 7827 4 ALE
rlabel m2contact 7137 7731 7137 7731 4 StatusReg[3]
rlabel m2contact 6633 7851 6633 7851 4 LrWe
rlabel m2contact 6573 7851 6573 7851 4 OpcodeCondIn[6]
rlabel m2contact 6537 7755 6537 7755 4 OpcodeCondIn[5]
rlabel m2contact 6345 7755 6345 7755 4 OpcodeCondIn[4]
rlabel m2contact 5709 7755 5709 7755 4 OpcodeCondIn[4]
rlabel m2contact 5241 7875 5241 7875 4 OpcodeCondIn[7]
rlabel m2contact 5097 7851 5097 7851 4 OpcodeCondIn[6]
rlabel m2contact 4425 7779 4425 7779 4 OpcodeCondIn[0]
rlabel m2contact 4089 7851 4089 7851 4 OpcodeCondIn[3]
rlabel metal2 3291 7875 3291 7875 4 OpcodeCondIn[2]
rlabel m2contact 3273 7875 3273 7875 4 OpcodeCondIn[2]
rlabel m2contact 3249 7851 3249 7851 4 OpcodeCondIn[3]
rlabel metal2 2883 7851 2883 7851 4 OpcodeCondIn[1]
rlabel m2contact 2865 7851 2865 7851 4 OpcodeCondIn[1]
rlabel m2contact 2331 7779 2331 7779 4 OpcodeCondIn[0]
rlabel m2contact 2313 7779 2313 7779 4 OpcodeCondIn[0]
rlabel m2contact 26457 5962 26457 5962 6 RwSel[0]
rlabel m2contact 26457 1882 26457 1882 6 RwSel[0]
rlabel m2contact 26433 4450 26433 4450 6 RwSel[1]
rlabel m2contact 26433 1858 26433 1858 6 RwSel[1]
rlabel m2contact 26409 2170 26409 2170 6 Flags[2]
rlabel m2contact 26385 5578 26385 5578 6 n_109
rlabel m2contact 26385 2338 26385 2338 6 n_109
rlabel m2contact 26361 4330 26361 4330 6 AluOR[0]
rlabel m2contact 26337 4570 26337 4570 6 n_310
rlabel m2contact 26313 4546 26313 4546 6 n_282
rlabel m2contact 26289 5386 26289 5386 6 n_266
rlabel m2contact 26289 4306 26289 4306 6 n_266
rlabel m2contact 26265 4618 26265 4618 6 n_349
rlabel m2contact 26241 4282 26241 4282 6 SysBus[3]
rlabel m2contact 26217 5290 26217 5290 6 n_351
rlabel m2contact 26181 4426 26181 4426 6 n_25
rlabel m2contact 26181 2530 26181 2530 6 n_25
rlabel m2contact 26169 5770 26169 5770 6 n_253
rlabel m2contact 26145 6394 26145 6394 6 n_163
rlabel m2contact 26121 5458 26121 5458 6 n_188
rlabel m2contact 26097 4330 26097 4330 6 AluOR[0]
rlabel m2contact 26073 5674 26073 5674 6 n_182
rlabel m2contact 26049 4594 26049 4594 6 AluOR[1]
rlabel m2contact 26025 4186 26025 4186 6 n_111
rlabel m2contact 26001 4714 26001 4714 6 n_190
rlabel m2contact 25977 2650 25977 2650 6 n_77
rlabel m2contact 25953 6706 25953 6706 6 n_20
rlabel m2contact 25953 3514 25953 3514 6 n_20
rlabel m2contact 25929 5818 25929 5818 6 n_32
rlabel m2contact 25929 5602 25929 5602 6 n_28
rlabel m2contact 25905 3538 25905 3538 6 stateSub[0]
rlabel m2contact 25881 5146 25881 5146 6 n_79
rlabel m2contact 25857 3322 25857 3322 6 n_81
rlabel m2contact 25857 3730 25857 3730 6 stateSub[1]
rlabel m2contact 25833 4234 25833 4234 6 n_215
rlabel m2contact 25833 4858 25833 4858 6 n_276
rlabel m2contact 25809 5842 25809 5842 6 n_332
rlabel m2contact 25809 4258 25809 4258 6 n_332
rlabel m2contact 25785 5194 25785 5194 6 n_198
rlabel m2contact 25761 4930 25761 4930 6 n_8
rlabel m2contact 25761 4642 25761 4642 6 n_248
rlabel m2contact 25737 5650 25737 5650 6 n_221
rlabel m2contact 25713 4402 25713 4402 6 OpcodeCondIn[1]
rlabel m2contact 25689 6346 25689 6346 6 n_126
rlabel m2contact 25665 2338 25665 2338 6 n_109
rlabel m2contact 25665 2362 25665 2362 6 n_113
rlabel m2contact 25641 6058 25641 6058 6 state[0]
rlabel m2contact 25641 2842 25641 2842 6 n_39
rlabel m2contact 25617 3850 25617 3850 6 n_74
rlabel m2contact 25617 3730 25617 3730 6 stateSub[1]
rlabel m2contact 25593 6250 25593 6250 6 n_91
rlabel m2contact 25593 1954 25593 1954 6 n_91
rlabel m2contact 25569 6514 25569 6514 6 n_374
rlabel m2contact 25545 5386 25545 5386 6 n_266
rlabel m2contact 25545 5362 25545 5362 6 n_85
rlabel m2contact 25521 4834 25521 4834 6 n_318
rlabel m2contact 25521 4330 25521 4330 6 n_185
rlabel m2contact 25497 6226 25497 6226 6 n_224
rlabel m2contact 25497 2386 25497 2386 6 n_224
rlabel m2contact 25473 2530 25473 2530 6 n_25
rlabel m2contact 25473 2554 25473 2554 6 n_89
rlabel m2contact 25449 3514 25449 3514 6 n_20
rlabel m2contact 25449 3538 25449 3538 6 stateSub[0]
rlabel m2contact 25425 5698 25425 5698 6 n_66
rlabel m2contact 25425 3778 25425 3778 6 n_30
rlabel m2contact 25401 3322 25401 3322 6 n_81
rlabel m2contact 25377 6754 25377 6754 6 n_250
rlabel m2contact 25377 4210 25377 4210 6 n_250
rlabel m2contact 25365 3946 25365 3946 6 n_122
rlabel m2contact 25365 3706 25365 3706 6 n_122
rlabel m2contact 25353 5698 25353 5698 6 n_66
rlabel m2contact 25329 3610 25329 3610 6 OpcodeCondIn[7]
rlabel m2contact 25305 3706 25305 3706 6 n_122
rlabel m2contact 25305 3730 25305 3730 6 stateSub[1]
rlabel m2contact 25281 4642 25281 4642 6 n_248
rlabel m2contact 25245 4354 25245 4354 6 n_340
rlabel m2contact 25245 2578 25245 2578 6 n_340
rlabel m2contact 25233 5290 25233 5290 6 n_351
rlabel m2contact 25209 5290 25209 5290 6 n_351
rlabel m2contact 25185 4690 25185 4690 6 OpcodeCondIn[2]
rlabel m2contact 25161 5842 25161 5842 6 n_332
rlabel m2contact 25161 5794 25161 5794 6 n_252
rlabel m2contact 25137 4882 25137 4882 6 n_222
rlabel m2contact 25137 3418 25137 3418 6 n_222
rlabel m2contact 25113 6250 25113 6250 6 n_91
rlabel m2contact 25113 6202 25113 6202 6 n_264
rlabel m2contact 25089 4210 25089 4210 6 n_250
rlabel m2contact 25089 5002 25089 5002 6 n_178
rlabel m2contact 25065 2794 25065 2794 6 n_57
rlabel m2contact 25041 5218 25041 5218 6 n_244
rlabel m2contact 25017 6730 25017 6730 6 n_95
rlabel m2contact 24993 4354 24993 4354 6 n_340
rlabel m2contact 24993 3442 24993 3442 6 n_243
rlabel m2contact 24969 6178 24969 6178 6 n_312
rlabel m2contact 24945 4378 24945 4378 6 n_233
rlabel m2contact 24921 6298 24921 6298 6 n_162
rlabel m2contact 24897 2074 24897 2074 6 n_268
rlabel m2contact 24897 2818 24897 2818 6 OpcodeCondIn[4]
rlabel m2contact 24873 3514 24873 3514 6 n_239
rlabel m2contact 24849 4162 24849 4162 6 n_75
rlabel m2contact 24825 5098 24825 5098 6 OpcodeCondIn[6]
rlabel m2contact 24825 3610 24825 3610 6 OpcodeCondIn[7]
rlabel m2contact 24801 2602 24801 2602 6 n_114
rlabel m2contact 24777 5074 24777 5074 6 n_216
rlabel m2contact 24753 2434 24753 2434 6 n_214
rlabel m2contact 24729 4234 24729 4234 6 n_215
rlabel m2contact 24729 3634 24729 3634 6 n_237
rlabel m2contact 24705 4858 24705 4858 6 n_276
rlabel m2contact 24681 3898 24681 3898 6 OpcodeCondIn[3]
rlabel m2contact 24657 6778 24657 6778 6 n_285
rlabel m2contact 24633 3346 24633 3346 6 n_284
rlabel m2contact 24609 6226 24609 6226 6 n_224
rlabel m2contact 24609 6202 24609 6202 6 n_264
rlabel m2contact 24585 4882 24585 4882 6 n_222
rlabel m2contact 24585 4810 24585 4810 6 n_86
rlabel m2contact 24561 6370 24561 6370 6 n_206
rlabel m2contact 24537 5866 24537 5866 6 n_104
rlabel m2contact 24513 4354 24513 4354 6 n_196
rlabel m2contact 24513 3322 24513 3322 6 n_81
rlabel m2contact 24489 4114 24489 4114 6 n_195
rlabel m2contact 24465 4474 24465 4474 6 n_140
rlabel m2contact 24441 6298 24441 6298 6 n_162
rlabel m2contact 24393 4738 24393 4738 6 n_43
rlabel m2contact 24369 5122 24369 5122 6 n_42
rlabel m2contact 24345 5698 24345 5698 6 n_66
rlabel m2contact 24345 3730 24345 3730 6 stateSub[1]
rlabel m2contact 24297 4066 24297 4066 6 n_101
rlabel m2contact 24273 6538 24273 6538 6 stateSub[2]
rlabel m2contact 24249 3298 24249 3298 6 n_84
rlabel m2contact 24201 3490 24201 3490 6 n_169
rlabel m2contact 24177 2818 24177 2818 6 OpcodeCondIn[4]
rlabel m2contact 24153 4330 24153 4330 6 n_185
rlabel m2contact 24105 3994 24105 3994 6 n_302
rlabel m2contact 24081 4090 24081 4090 6 n_267
rlabel m2contact 24057 2074 24057 2074 6 n_268
rlabel m2contact 24033 4642 24033 4642 6 n_248
rlabel m2contact 23985 4522 23985 4522 6 n_323
rlabel m2contact 23937 2194 23937 2194 6 n_327
rlabel m2contact 23889 6634 23889 6634 6 n_60
rlabel m2contact 23865 5314 23865 5314 6 n_26
rlabel m2contact 23841 6658 23841 6658 6 n_12
rlabel m2contact 23817 4906 23817 4906 6 n_97
rlabel m2contact 23793 6538 23793 6538 6 stateSub[2]
rlabel m2contact 23793 4210 23793 4210 6 stateSub[2]
rlabel m2contact 23769 4210 23769 4210 6 stateSub[2]
rlabel m2contact 23769 5410 23769 5410 6 n_151
rlabel m2contact 23721 4114 23721 4114 6 n_195
rlabel m2contact 23721 2530 23721 2530 6 n_354
rlabel m2contact 23697 3058 23697 3058 6 n_155
rlabel m2contact 23673 4474 23673 4474 6 n_140
rlabel m2contact 23649 4210 23649 4210 6 n_211
rlabel m2contact 23625 6082 23625 6082 6 n_108
rlabel m2contact 23601 4282 23601 4282 6 SysBus[3]
rlabel m2contact 23577 6418 23577 6418 6 n_149
rlabel m2contact 23553 3898 23553 3898 6 OpcodeCondIn[3]
rlabel m2contact 23529 3802 23529 3802 6 n_136
rlabel m2contact 23505 2770 23505 2770 6 n_189
rlabel m2contact 23481 6106 23481 6106 6 n_165
rlabel m2contact 23481 3130 23481 3130 6 n_165
rlabel m2contact 23457 6106 23457 6106 6 n_165
rlabel m2contact 23457 6058 23457 6058 6 state[0]
rlabel m2contact 23433 3514 23433 3514 6 n_239
rlabel m2contact 23409 3226 23409 3226 6 n_53
rlabel m2contact 23409 3730 23409 3730 6 stateSub[1]
rlabel m2contact 23385 1978 23385 1978 6 n_137
rlabel m2contact 23337 4474 23337 4474 6 n_371
rlabel m2contact 23313 4618 23313 4618 6 n_349
rlabel m2contact 23289 4522 23289 4522 6 n_323
rlabel m2contact 23265 6010 23265 6010 6 n_292
rlabel m2contact 23217 5554 23217 5554 6 n_51
rlabel m2contact 23193 5098 23193 5098 6 OpcodeCondIn[6]
rlabel m2contact 23169 6274 23169 6274 6 n_50
rlabel m2contact 23145 5986 23145 5986 6 n_231
rlabel m2contact 23145 4138 23145 4138 6 n_231
rlabel m2contact 23121 5386 23121 5386 6 n_121
rlabel m2contact 23121 3394 23121 3394 6 n_121
rlabel m2contact 23097 4282 23097 4282 6 n_234
rlabel m2contact 23073 4522 23073 4522 6 n_193
rlabel m2contact 23049 5986 23049 5986 6 n_231
rlabel m2contact 23049 5938 23049 5938 6 n_308
rlabel m2contact 23025 5482 23025 5482 6 n_17
rlabel m2contact 23025 3466 23025 3466 6 n_17
rlabel m2contact 23001 5026 23001 5026 6 n_110
rlabel m2contact 22977 6058 22977 6058 6 state[0]
rlabel m2contact 22977 2458 22977 2458 6 state[0]
rlabel m2contact 22953 2290 22953 2290 6 n_31
rlabel m2contact 22929 4138 22929 4138 6 n_231
rlabel m2contact 22929 6154 22929 6154 6 n_69
rlabel m2contact 22905 2770 22905 2770 6 n_189
rlabel m2contact 22881 4522 22881 4522 6 n_193
rlabel m2contact 22857 3946 22857 3946 6 n_122
rlabel m2contact 22833 4714 22833 4714 6 n_190
rlabel m2contact 22809 3394 22809 3394 6 n_121
rlabel m2contact 22809 3514 22809 3514 6 n_239
rlabel m2contact 22785 4330 22785 4330 6 n_185
rlabel m2contact 22761 4498 22761 4498 6 Rs1Sel[1]
rlabel m2contact 22737 4570 22737 4570 6 n_310
rlabel m2contact 22713 3466 22713 3466 6 n_17
rlabel m2contact 22713 3562 22713 3562 6 n_321
rlabel m2contact 22689 2458 22689 2458 6 state[0]
rlabel m2contact 22689 2482 22689 2482 6 n_364
rlabel m2contact 22665 6442 22665 6442 6 n_269
rlabel m2contact 22665 4642 22665 4642 6 n_248
rlabel m2contact 22617 3274 22617 3274 6 StatusRegEn
rlabel m2contact 22569 3106 22569 3106 6 n_294
rlabel m2contact 22545 4114 22545 4114 6 n_195
rlabel m2contact 22521 2146 22521 2146 6 n_172
rlabel m2contact 22497 2074 22497 2074 6 n_268
rlabel m2contact 22473 6802 22473 6802 6 n_105
rlabel m2contact 22473 3706 22473 3706 6 nWait
rlabel m2contact 22449 2986 22449 2986 6 n_257
rlabel m2contact 22425 5626 22425 5626 6 n_340
rlabel m2contact 22425 2578 22425 2578 6 n_340
rlabel m2contact 22401 5626 22401 5626 6 n_340
rlabel m2contact 22401 5530 22401 5530 6 n_288
rlabel m2contact 22377 2098 22377 2098 6 n_345
rlabel m2contact 22353 2314 22353 2314 6 n_335
rlabel m2contact 22305 4450 22305 4450 6 RwSel[1]
rlabel m2contact 22281 3682 22281 3682 6 n_359
rlabel m2contact 22281 3250 22281 3250 6 n_199
rlabel m2contact 22257 2482 22257 2482 6 n_364
rlabel m2contact 22233 4018 22233 4018 6 n_203
rlabel m2contact 22209 6202 22209 6202 6 n_264
rlabel m2contact 22185 4234 22185 4234 6 n_215
rlabel m2contact 22161 5914 22161 5914 6 n_296
rlabel m2contact 22137 4282 22137 4282 6 n_234
rlabel m2contact 22113 5050 22113 5050 6 n_281
rlabel m2contact 22089 4450 22089 4450 6 n_235
rlabel m2contact 22065 5170 22065 5170 6 n_80
rlabel m2contact 22041 3274 22041 3274 6 StatusRegEn
rlabel m2contact 22041 3298 22041 3298 6 n_84
rlabel m2contact 22017 5242 22017 5242 6 n_88
rlabel m2contact 21993 4978 21993 4978 6 n_226
rlabel m2contact 21969 5722 21969 5722 6 n_76
rlabel m2contact 21969 2986 21969 2986 6 n_257
rlabel m2contact 21945 5098 21945 5098 6 OpcodeCondIn[6]
rlabel m2contact 21921 6274 21921 6274 6 n_50
rlabel m2contact 21921 5506 21921 5506 6 n_289
rlabel m2contact 21897 2818 21897 2818 6 OpcodeCondIn[4]
rlabel m2contact 21873 6538 21873 6538 6 stateSub[2]
rlabel m2contact 21873 4282 21873 4282 6 stateSub[2]
rlabel m2contact 21849 4282 21849 4282 6 stateSub[2]
rlabel m2contact 21849 6034 21849 6034 6 AluWe
rlabel m2contact 21801 5890 21801 5890 6 n_314
rlabel m2contact 21729 5794 21729 5794 6 n_252
rlabel m2contact 21705 4786 21705 4786 6 StatusReg[0]
rlabel m2contact 21657 2218 21657 2218 6 n_484
rlabel m2contact 21633 4690 21633 4690 6 OpcodeCondIn[2]
rlabel m2contact 21609 3610 21609 3610 6 OpcodeCondIn[7]
rlabel m2contact 21513 4402 21513 4402 6 OpcodeCondIn[1]
rlabel m2contact 21489 4138 21489 4138 6 n_13
rlabel m2contact 21369 5338 21369 5338 6 n_305
rlabel m2contact 21321 5266 21321 5266 6 n_373
rlabel m2contact 21321 2026 21321 2026 6 n_373
rlabel m2contact 21297 5266 21297 5266 6 n_373
rlabel m2contact 21297 5098 21297 5098 6 OpcodeCondIn[6]
rlabel m2contact 21273 3538 21273 3538 6 stateSub[0]
rlabel m2contact 21249 3898 21249 3898 6 OpcodeCondIn[3]
rlabel m2contact 21225 4522 21225 4522 6 n_122
rlabel m2contact 21225 3946 21225 3946 6 n_122
rlabel m2contact 21201 6106 21201 6106 6 n_99
rlabel m2contact 21201 1930 21201 1930 6 n_99
rlabel m2contact 21177 6754 21177 6754 6 n_250
rlabel m2contact 21177 4954 21177 4954 6 n_209
rlabel m2contact 21153 4858 21153 4858 6 n_276
rlabel m2contact 21153 4042 21153 4042 6 n_313
rlabel m2contact 21129 3226 21129 3226 6 n_53
rlabel m2contact 21105 4498 21105 4498 6 n_189
rlabel m2contact 21105 2770 21105 2770 6 n_189
rlabel m2contact 21081 6802 21081 6802 6 n_105
rlabel m2contact 21081 6706 21081 6706 6 n_20
rlabel m2contact 21057 6106 21057 6106 6 n_99
rlabel m2contact 21057 5386 21057 5386 6 n_121
rlabel m2contact 21033 4642 21033 4642 6 n_248
rlabel m2contact 21009 5626 21009 5626 6 n_130
rlabel m2contact 20985 4162 20985 4162 6 n_75
rlabel m2contact 20985 5746 20985 5746 6 n_78
rlabel m2contact 20961 4522 20961 4522 6 n_122
rlabel m2contact 20961 4210 20961 4210 6 n_211
rlabel m2contact 20937 2650 20937 2650 6 n_77
rlabel m2contact 20913 5386 20913 5386 6 n_121
rlabel m2contact 20913 3658 20913 3658 6 n_121
rlabel m2contact 20889 3970 20889 3970 6 IrWe
rlabel m2contact 20865 4642 20865 4642 6 n_248
rlabel m2contact 20841 6106 20841 6106 6 n_99
rlabel m2contact 20841 6058 20841 6058 6 state[0]
rlabel m2contact 20817 5098 20817 5098 6 OpcodeCondIn[6]
rlabel m2contact 20793 4498 20793 4498 6 n_189
rlabel m2contact 20793 3010 20793 3010 6 n_160
rlabel m2contact 20769 5266 20769 5266 6 n_55
rlabel m2contact 20769 4282 20769 4282 6 n_55
rlabel m2contact 20745 3658 20745 3658 6 n_121
rlabel m2contact 20745 3754 20745 3754 6 n_200
rlabel m2contact 20721 5626 20721 5626 6 n_130
rlabel m2contact 20721 4210 20721 4210 6 n_211
rlabel m2contact 20697 3250 20697 3250 6 n_199
rlabel m2contact 20673 5578 20673 5578 6 n_109
rlabel m2contact 20649 4498 20649 4498 6 Op2Sel[1]
rlabel m2contact 20625 5002 20625 5002 6 n_178
rlabel m2contact 20601 5266 20601 5266 6 n_55
rlabel m2contact 20601 4954 20601 4954 6 n_209
rlabel m2contact 20577 2746 20577 2746 6 n_485
rlabel m2contact 20529 3970 20529 3970 6 IrWe
rlabel m2contact 20505 5266 20505 5266 6 n_156
rlabel m2contact 20481 6490 20481 6490 6 OpcodeCondIn[5]
rlabel m2contact 20481 2554 20481 2554 6 n_89
rlabel m2contact 20457 4330 20457 4330 6 n_185
rlabel m2contact 20433 6106 20433 6106 6 n_72
rlabel m2contact 20409 2050 20409 2050 6 n_103
rlabel m2contact 20385 6538 20385 6538 6 stateSub[2]
rlabel m2contact 20385 4642 20385 4642 6 n_248
rlabel m2contact 20361 6250 20361 6250 6 n_83
rlabel m2contact 20361 6202 20361 6202 6 n_264
rlabel m2contact 20313 5842 20313 5842 6 n_48
rlabel m2contact 20313 3178 20313 3178 6 n_23
rlabel m2contact 20289 5434 20289 5434 6 n_22
rlabel m2contact 20289 3466 20289 3466 6 n_22
rlabel m2contact 20265 3610 20265 3610 6 OpcodeCondIn[7]
rlabel m2contact 20241 3466 20241 3466 6 n_22
rlabel m2contact 20241 3514 20241 3514 6 n_239
rlabel m2contact 20217 6226 20217 6226 6 n_273
rlabel m2contact 20217 3970 20217 3970 6 n_273
rlabel m2contact 20193 4186 20193 4186 6 n_111
rlabel m2contact 20193 4618 20193 4618 6 n_207
rlabel m2contact 20169 4882 20169 4882 6 n_171
rlabel m2contact 20169 3514 20169 3514 6 n_239
rlabel m2contact 20145 5986 20145 5986 6 n_70
rlabel m2contact 20145 6754 20145 6754 6 n_250
rlabel m2contact 20109 4258 20109 4258 6 n_332
rlabel m2contact 20109 2122 20109 2122 6 n_332
rlabel m2contact 20097 4522 20097 4522 6 n_98
rlabel m2contact 20073 5386 20073 5386 6 n_121
rlabel m2contact 20049 3970 20049 3970 6 n_273
rlabel m2contact 20049 4186 20049 4186 6 n_44
rlabel m2contact 20025 6466 20025 6466 6 n_345
rlabel m2contact 20025 2098 20025 2098 6 n_345
rlabel m2contact 20001 2314 20001 2314 6 n_335
rlabel m2contact 20001 2338 20001 2338 6 n_329
rlabel m2contact 19977 5530 19977 5530 6 n_288
rlabel m2contact 19953 2122 19953 2122 6 n_332
rlabel m2contact 19953 2194 19953 2194 6 n_327
rlabel m2contact 19929 4690 19929 4690 6 OpcodeCondIn[2]
rlabel m2contact 19929 3970 19929 3970 6 OpcodeCondIn[2]
rlabel m2contact 19905 6466 19905 6466 6 n_345
rlabel m2contact 19905 6130 19905 6130 6 n_6
rlabel m2contact 19881 1858 19881 1858 6 n_167
rlabel m2contact 19857 3970 19857 3970 6 OpcodeCondIn[2]
rlabel m2contact 19857 4042 19857 4042 6 n_313
rlabel m2contact 19833 5098 19833 5098 6 OpcodeCondIn[6]
rlabel m2contact 19809 5578 19809 5578 6 n_109
rlabel m2contact 19809 3466 19809 3466 6 n_109
rlabel m2contact 19785 3802 19785 3802 6 n_136
rlabel m2contact 19785 4450 19785 4450 6 n_235
rlabel m2contact 19761 3610 19761 3610 6 OpcodeCondIn[7]
rlabel m2contact 19737 3466 19737 3466 6 n_109
rlabel m2contact 19737 3490 19737 3490 6 n_169
rlabel m2contact 19713 4666 19713 4666 6 n_53
rlabel m2contact 19713 3226 19713 3226 6 n_53
rlabel m2contact 19689 3370 19689 3370 6 n_183
rlabel m2contact 19665 5410 19665 5410 6 n_151
rlabel m2contact 19665 2962 19665 2962 6 n_159
rlabel m2contact 19641 3658 19641 3658 6 n_205
rlabel m2contact 19617 3394 19617 3394 6 n_220
rlabel m2contact 19617 3538 19617 3538 6 stateSub[0]
rlabel m2contact 19593 5434 19593 5434 6 n_22
rlabel m2contact 19593 3202 19593 3202 6 n_22
rlabel m2contact 19569 4018 19569 4018 6 n_203
rlabel m2contact 19569 4954 19569 4954 6 n_209
rlabel m2contact 19545 3010 19545 3010 6 n_160
rlabel m2contact 19521 2938 19521 2938 6 n_210
rlabel m2contact 19521 4690 19521 4690 6 OpcodeCondIn[2]
rlabel m2contact 19497 4930 19497 4930 6 n_8
rlabel m2contact 19473 4762 19473 4762 6 n_251
rlabel m2contact 19473 2674 19473 2674 6 n_251
rlabel m2contact 19449 3874 19449 3874 6 n_194
rlabel m2contact 19425 3274 19425 3274 6 n_170
rlabel m2contact 19401 2194 19401 2194 6 n_327
rlabel m2contact 19401 2986 19401 2986 6 n_257
rlabel m2contact 19377 3538 19377 3538 6 stateSub[0]
rlabel m2contact 19341 4330 19341 4330 6 n_185
rlabel m2contact 19341 3586 19341 3586 6 n_185
rlabel m2contact 19329 5002 19329 5002 6 n_178
rlabel m2contact 19329 3514 19329 3514 6 n_239
rlabel m2contact 19305 6754 19305 6754 6 n_250
rlabel m2contact 19305 3826 19305 3826 6 n_250
rlabel m2contact 19281 6490 19281 6490 6 OpcodeCondIn[5]
rlabel m2contact 19257 4402 19257 4402 6 OpcodeCondIn[1]
rlabel m2contact 19233 2938 19233 2938 6 n_210
rlabel m2contact 19209 3970 19209 3970 6 n_15
rlabel m2contact 19185 4666 19185 4666 6 n_53
rlabel m2contact 19185 3898 19185 3898 6 OpcodeCondIn[3]
rlabel m2contact 19161 3586 19161 3586 6 n_185
rlabel m2contact 19161 3730 19161 3730 6 stateSub[1]
rlabel m2contact 19137 4666 19137 4666 6 n_267
rlabel m2contact 19137 4090 19137 4090 6 n_267
rlabel m2contact 19113 2698 19113 2698 6 n_202
rlabel m2contact 19089 3202 19089 3202 6 n_22
rlabel m2contact 19089 3274 19089 3274 6 n_170
rlabel m2contact 19065 2938 19065 2938 6 n_210
rlabel m2contact 19041 3922 19041 3922 6 n_34
rlabel m2contact 19017 2722 19017 2722 6 n_38
rlabel m2contact 18993 3634 18993 3634 6 n_237
rlabel m2contact 18969 2674 18969 2674 6 n_251
rlabel m2contact 18969 2842 18969 2842 6 n_39
rlabel m2contact 18945 6610 18945 6610 6 n_208
rlabel m2contact 18921 3826 18921 3826 6 n_250
rlabel m2contact 18921 4018 18921 4018 6 n_271
rlabel m2contact 18897 3586 18897 3586 6 n_115
rlabel m2contact 18873 3418 18873 3418 6 n_222
rlabel m2contact 18873 3442 18873 3442 6 n_243
rlabel m2contact 18849 3394 18849 3394 6 n_220
rlabel m2contact 18825 6442 18825 6442 6 n_269
rlabel m2contact 18825 5650 18825 5650 6 n_221
rlabel m2contact 18801 4666 18801 4666 6 n_267
rlabel m2contact 18801 4642 18801 4642 6 n_248
rlabel m2contact 18777 2074 18777 2074 6 n_268
rlabel m2contact 18729 4666 18729 4666 6 n_262
rlabel m2contact 18705 3634 18705 3634 6 n_237
rlabel m2contact 18681 4450 18681 4450 6 n_235
rlabel m2contact 18657 5842 18657 5842 6 n_48
rlabel m2contact 18585 4930 18585 4930 6 n_174
rlabel m2contact 18537 5626 18537 5626 6 n_130
rlabel m2contact 18489 5626 18489 5626 6 n_148
rlabel m2contact 18441 2266 18441 2266 6 n_52
rlabel m2contact 18417 6346 18417 6346 6 n_126
rlabel m2contact 18369 4570 18369 4570 6 n_310
rlabel m2contact 18345 5242 18345 5242 6 n_88
rlabel m2contact 18321 4234 18321 4234 6 n_215
rlabel m2contact 18273 2434 18273 2434 6 n_214
rlabel m2contact 18249 4114 18249 4114 6 n_195
rlabel m2contact 18225 2314 18225 2314 6 n_131
rlabel m2contact 18165 4090 18165 4090 6 n_267
rlabel m2contact 18165 2410 18165 2410 6 n_267
rlabel m2contact 18153 6274 18153 6274 6 n_50
rlabel m2contact 18129 3850 18129 3850 6 n_74
rlabel m2contact 18105 3514 18105 3514 6 n_239
rlabel m2contact 18081 6538 18081 6538 6 stateSub[2]
rlabel m2contact 18057 2122 18057 2122 6 n_33
rlabel m2contact 18057 3898 18057 3898 6 OpcodeCondIn[3]
rlabel m2contact 18033 6490 18033 6490 6 OpcodeCondIn[5]
rlabel m2contact 18009 3202 18009 3202 6 n_45
rlabel m2contact 17985 2002 17985 2002 6 PcEn
rlabel m2contact 17961 6538 17961 6538 6 stateSub[2]
rlabel m2contact 17937 6154 17937 6154 6 n_69
rlabel m2contact 17937 3826 17937 3826 6 n_58
rlabel m2contact 17913 5314 17913 5314 6 n_26
rlabel m2contact 17913 3850 17913 3850 6 n_26
rlabel m2contact 17889 4306 17889 4306 6 n_266
rlabel m2contact 17889 6058 17889 6058 6 state[0]
rlabel m2contact 17865 2410 17865 2410 6 n_267
rlabel m2contact 17865 2458 17865 2458 6 n_217
rlabel m2contact 17841 2986 17841 2986 6 n_257
rlabel m2contact 17817 6082 17817 6082 6 n_108
rlabel m2contact 17793 3850 17793 3850 6 n_26
rlabel m2contact 17793 3898 17793 3898 6 OpcodeCondIn[3]
rlabel m2contact 17769 5578 17769 5578 6 n_109
rlabel m2contact 17769 3610 17769 3610 6 OpcodeCondIn[7]
rlabel m2contact 17745 3946 17745 3946 6 n_122
rlabel m2contact 17721 5578 17721 5578 6 n_49
rlabel m2contact 17697 3634 17697 3634 6 n_237
rlabel m2contact 17673 5842 17673 5842 6 n_48
rlabel m2contact 17625 5842 17625 5842 6 n_247
rlabel m2contact 17625 2314 17625 2314 6 n_131
rlabel m2contact 17601 4354 17601 4354 6 n_196
rlabel m2contact 17577 5458 17577 5458 6 n_188
rlabel m2contact 17553 2770 17553 2770 6 n_189
rlabel m2contact 17529 1906 17529 1906 6 n_315
rlabel m2contact 17505 3778 17505 3778 6 n_30
rlabel m2contact 17481 2410 17481 2410 6 n_263
rlabel m2contact 17457 5890 17457 5890 6 n_314
rlabel m2contact 17433 5482 17433 5482 6 n_17
rlabel m2contact 17433 5098 17433 5098 6 OpcodeCondIn[6]
rlabel m2contact 17409 2866 17409 2866 6 n_14
rlabel m2contact 17385 4354 17385 4354 6 WdSel
rlabel m2contact 17337 4786 17337 4786 6 StatusReg[0]
rlabel m2contact 17313 3106 17313 3106 6 n_294
rlabel m2contact 17241 2962 17241 2962 6 n_159
rlabel m2contact 17241 3082 17241 3082 6 CFlag
rlabel m2contact 17217 3418 17217 3418 6 n_255
rlabel m2contact 17145 4306 17145 4306 6 n_153
rlabel m2contact 17121 4330 17121 4330 6 n_185
rlabel m2contact 17049 3514 17049 3514 6 n_239
rlabel m2contact 16953 3898 16953 3898 6 OpcodeCondIn[3]
rlabel m2contact 16929 5650 16929 5650 6 n_221
rlabel m2contact 16905 4642 16905 4642 6 n_248
rlabel m2contact 16881 5530 16881 5530 6 n_288
rlabel m2contact 16833 3034 16833 3034 6 n_372
rlabel m2contact 16809 3538 16809 3538 6 stateSub[0]
rlabel m2contact 16785 2674 16785 2674 6 n_100
rlabel m2contact 16713 3466 16713 3466 6 n_146
rlabel m2contact 16689 6490 16689 6490 6 OpcodeCondIn[5]
rlabel m2contact 16665 4282 16665 4282 6 n_55
rlabel m2contact 16665 5098 16665 5098 6 OpcodeCondIn[6]
rlabel m2contact 16641 6058 16641 6058 6 state[0]
rlabel m2contact 16641 3850 16641 3850 6 state[0]
rlabel m2contact 16617 5458 16617 5458 6 n_188
rlabel m2contact 16593 3970 16593 3970 6 n_15
rlabel m2contact 16569 3154 16569 3154 6 n_96
rlabel m2contact 16569 3226 16569 3226 6 n_53
rlabel m2contact 16545 4642 16545 4642 6 n_248
rlabel m2contact 16521 3130 16521 3130 6 n_165
rlabel m2contact 16497 3970 16497 3970 6 n_142
rlabel m2contact 16473 3898 16473 3898 6 OpcodeCondIn[3]
rlabel m2contact 16449 2458 16449 2458 6 n_217
rlabel m2contact 16425 3850 16425 3850 6 state[0]
rlabel m2contact 16425 5458 16425 5458 6 n_150
rlabel m2contact 16401 5410 16401 5410 6 n_151
rlabel m2contact 16377 6514 16377 6514 6 n_374
rlabel m2contact 16377 3850 16377 3850 6 n_374
rlabel m2contact 16353 3850 16353 3850 6 n_374
rlabel m2contact 16353 5482 16353 5482 6 n_147
rlabel m2contact 16329 2506 16329 2506 6 n_362
rlabel m2contact 16329 3466 16329 3466 6 n_146
rlabel m2contact 16305 4522 16305 4522 6 n_98
rlabel m2contact 16281 4426 16281 4426 6 n_25
rlabel m2contact 16281 3682 16281 3682 6 n_359
rlabel m2contact 16257 4522 16257 4522 6 n_286
rlabel m2contact 16257 3130 16257 3130 6 n_286
rlabel m2contact 16233 2890 16233 2890 6 n_184
rlabel m2contact 16209 4258 16209 4258 6 n_332
rlabel m2contact 16185 3898 16185 3898 6 OpcodeCondIn[3]
rlabel m2contact 16161 3130 16161 3130 6 n_286
rlabel m2contact 16161 3370 16161 3370 6 n_183
rlabel m2contact 16137 4426 16137 4426 6 n_35
rlabel m2contact 16137 3850 16137 3850 6 n_35
rlabel m2contact 16113 6706 16113 6706 6 n_20
rlabel m2contact 16113 6682 16113 6682 6 n_62
rlabel m2contact 16089 6082 16089 6082 6 n_167
rlabel m2contact 16089 1858 16089 1858 6 n_167
rlabel m2contact 16065 3850 16065 3850 6 n_35
rlabel m2contact 16065 3898 16065 3898 6 OpcodeCondIn[3]
rlabel m2contact 16041 6490 16041 6490 6 OpcodeCondIn[5]
rlabel m2contact 16017 6706 16017 6706 6 n_47
rlabel m2contact 16017 1882 16017 1882 6 n_47
rlabel m2contact 15993 6082 15993 6082 6 n_167
rlabel m2contact 15993 3010 15993 3010 6 n_160
rlabel m2contact 15969 3658 15969 3658 6 n_205
rlabel m2contact 15945 5530 15945 5530 6 n_288
rlabel m2contact 15921 1882 15921 1882 6 n_47
rlabel m2contact 15921 2242 15921 2242 6 n_65
rlabel m2contact 15897 5530 15897 5530 6 n_288
rlabel m2contact 15873 5986 15873 5986 6 n_70
rlabel m2contact 15849 2914 15849 2914 6 n_19
rlabel m2contact 15825 4954 15825 4954 6 n_209
rlabel m2contact 15801 5002 15801 5002 6 n_178
rlabel m2contact 15777 5938 15777 5938 6 n_308
rlabel m2contact 15777 4930 15777 4930 6 n_174
rlabel m2contact 15753 6202 15753 6202 6 n_264
rlabel m2contact 15729 5866 15729 5866 6 n_104
rlabel m2contact 15705 5842 15705 5842 6 n_247
rlabel m2contact 15681 4258 15681 4258 6 n_59
rlabel m2contact 15609 5818 15609 5818 6 n_32
rlabel m2contact 15585 5626 15585 5626 6 n_148
rlabel m2contact 15561 6562 15561 6562 6 n_120
rlabel m2contact 15537 6106 15537 6106 6 n_72
rlabel m2contact 15489 5338 15489 5338 6 n_305
rlabel m2contact 15465 4378 15465 4378 6 n_233
rlabel m2contact 15441 5218 15441 5218 6 n_244
rlabel m2contact 15417 4378 15417 4378 6 n_186
rlabel m2contact 15393 4666 15393 4666 6 n_262
rlabel m2contact 15345 3850 15345 3850 6 nWE
rlabel m2contact 15321 6586 15321 6586 6 n_54
rlabel m2contact 15297 4666 15297 4666 6 n_249
rlabel m2contact 15273 5074 15273 5074 6 n_216
rlabel m2contact 15249 5842 15249 5842 6 n_277
rlabel m2contact 15201 5050 15201 5050 6 n_281
rlabel m2contact 15177 6442 15177 6442 6 n_197
rlabel m2contact 15153 5026 15153 5026 6 n_110
rlabel m2contact 15129 6082 15129 6082 6 n_68
rlabel m2contact 15105 4090 15105 4090 6 n_267
rlabel m2contact 15105 4906 15105 4906 6 n_97
rlabel m2contact 15057 3250 15057 3250 6 n_199
rlabel m2contact 15057 4090 15057 4090 6 n_27
rlabel m2contact 15033 3226 15033 3226 6 n_53
rlabel m2contact 15009 2458 15009 2458 6 n_217
rlabel m2contact 15009 3130 15009 3130 6 state[1]
rlabel m2contact 14985 4906 14985 4906 6 n_180
rlabel m2contact 14985 1882 14985 1882 6 n_180
rlabel m2contact 14961 4906 14961 4906 6 n_180
rlabel m2contact 14961 3778 14961 3778 6 n_30
rlabel m2contact 14937 4738 14937 4738 6 n_43
rlabel m2contact 14937 4234 14937 4234 6 n_215
rlabel m2contact 14913 2626 14913 2626 6 n_135
rlabel m2contact 14889 5218 14889 5218 6 n_175
rlabel m2contact 14865 4738 14865 4738 6 n_191
rlabel m2contact 14841 4330 14841 4330 6 n_185
rlabel m2contact 14817 4930 14817 4930 6 n_174
rlabel m2contact 14769 5986 14769 5986 6 n_299
rlabel m2contact 14769 6538 14769 6538 6 stateSub[2]
rlabel m2contact 14721 1882 14721 1882 6 n_180
rlabel m2contact 14721 4642 14721 4642 6 n_248
rlabel m2contact 14625 6202 14625 6202 6 n_264
rlabel m2contact 14529 2026 14529 2026 6 n_373
rlabel m2contact 14481 2338 14481 2338 6 n_329
rlabel m2contact 14409 3274 14409 3274 6 n_170
rlabel m2contact 14385 4906 14385 4906 6 n_280
rlabel m2contact 14385 2026 14385 2026 6 n_280
rlabel m2contact 14361 4906 14361 4906 6 n_280
rlabel m2contact 14361 3946 14361 3946 6 n_122
rlabel m2contact 14337 5410 14337 5410 6 n_151
rlabel m2contact 14217 3298 14217 3298 6 n_84
rlabel m2contact 14145 2386 14145 2386 6 n_224
rlabel m2contact 14121 2650 14121 2650 6 n_77
rlabel m2contact 14097 2386 14097 2386 6 n_487
rlabel m2contact 14049 2194 14049 2194 6 n_327
rlabel m2contact 13905 2650 13905 2650 6 n_119
rlabel m2contact 13881 5938 13881 5938 6 n_127
rlabel m2contact 13857 2722 13857 2722 6 n_38
rlabel m2contact 13785 3538 13785 3538 6 stateSub[0]
rlabel m2contact 13761 2338 13761 2338 6 n_73
rlabel m2contact 13737 4474 13737 4474 6 n_371
rlabel m2contact 13713 3034 13713 3034 6 n_372
rlabel m2contact 13689 5866 13689 5866 6 n_352
rlabel m2contact 13665 5818 13665 5818 4 ImmSel
rlabel m2contact 13665 3034 13665 3034 4 ImmSel
rlabel m2contact 13641 6346 13641 6346 4 n_133
rlabel m2contact 13641 1882 13641 1882 4 n_133
rlabel m2contact 13617 4906 13617 4906 4 n_117
rlabel m2contact 13593 5026 13593 5026 4 n_168
rlabel m2contact 13593 6538 13593 6538 4 stateSub[2]
rlabel m2contact 13569 2074 13569 2074 4 n_268
rlabel m2contact 13545 4930 13545 4930 4 n_174
rlabel m2contact 13521 1858 13521 1858 4 n_167
rlabel m2contact 13521 2074 13521 2074 4 n_268
rlabel m2contact 13497 6154 13497 6154 4 n_164
rlabel m2contact 13497 2722 13497 2722 4 n_164
rlabel m2contact 13473 3034 13473 3034 4 ImmSel
rlabel m2contact 13473 3298 13473 3298 4 n_84
rlabel m2contact 13449 1882 13449 1882 4 n_133
rlabel m2contact 13449 5458 13449 5458 4 n_150
rlabel m2contact 13425 5074 13425 5074 4 n_9
rlabel m2contact 13425 3034 13425 3034 4 n_9
rlabel m2contact 13401 3346 13401 3346 4 n_284
rlabel m2contact 13377 4642 13377 4642 4 n_248
rlabel m2contact 13353 2722 13353 2722 4 n_164
rlabel m2contact 13353 5242 13353 5242 4 n_88
rlabel m2contact 13329 3034 13329 3034 4 n_9
rlabel m2contact 13329 3826 13329 3826 4 n_58
rlabel m2contact 13293 5386 13293 5386 4 n_121
rlabel m2contact 13293 3034 13293 3034 4 n_121
rlabel m2contact 13281 6274 13281 6274 4 n_293
rlabel m2contact 13257 2722 13257 2722 4 StatusReg[2]
rlabel m2contact 13233 3106 13233 3106 4 n_294
rlabel m2contact 13209 4114 13209 4114 4 n_195
rlabel m2contact 13185 2770 13185 2770 4 n_189
rlabel m2contact 13185 5338 13185 5338 4 n_93
rlabel m2contact 13161 3034 13161 3034 4 n_121
rlabel m2contact 13161 3538 13161 3538 4 stateSub[0]
rlabel m2contact 13137 2986 13137 2986 4 n_257
rlabel m2contact 13113 2842 13113 2842 4 n_39
rlabel m2contact 13089 1882 13089 1882 4 Flags[1]
rlabel m2contact 13065 5386 13065 5386 4 n_121
rlabel m2contact 13041 3226 13041 3226 4 n_53
rlabel m2contact 13017 5050 13017 5050 4 n_261
rlabel m2contact 12969 4162 12969 4162 4 n_75
rlabel m2contact 12969 4474 12969 4474 4 n_260
rlabel m2contact 12921 6466 12921 6466 4 n_368
rlabel m2contact 12921 4162 12921 4162 4 n_134
rlabel m2contact 12873 4114 12873 4114 4 PcSel[2]
rlabel m2contact 12849 1882 12849 1882 4 Flags[1]
rlabel m2contact 12849 3034 12849 3034 4 n_348
rlabel m2contact 12825 2194 12825 2194 4 n_327
rlabel m2contact 12801 5074 12801 5074 4 n_9
rlabel m2contact 12777 2794 12777 2794 4 n_57
rlabel m2contact 12753 4282 12753 4282 4 n_55
rlabel m2contact 12753 4786 12753 4786 4 StatusReg[0]
rlabel m2contact 12729 4402 12729 4402 4 OpcodeCondIn[1]
rlabel m2contact 12681 4786 12681 4786 4 n_275
rlabel m2contact 12657 6754 12657 6754 4 n_250
rlabel m2contact 12633 4282 12633 4282 4 n_272
rlabel m2contact 12561 2146 12561 2146 4 n_172
rlabel m2contact 12561 5530 12561 5530 4 n_288
rlabel m2contact 12537 5074 12537 5074 4 n_40
rlabel m2contact 12537 2794 12537 2794 4 n_40
rlabel m2contact 12513 4690 12513 4690 4 OpcodeCondIn[2]
rlabel m2contact 12489 5626 12489 5626 4 n_124
rlabel m2contact 12465 6322 12465 6322 4 Rs1Sel[0]
rlabel m2contact 12441 5794 12441 5794 4 n_252
rlabel m2contact 12441 4810 12441 4810 4 n_86
rlabel m2contact 12417 6322 12417 6322 4 n_176
rlabel m2contact 12393 5986 12393 5986 4 n_299
rlabel m2contact 12393 3538 12393 3538 4 stateSub[0]
rlabel m2contact 12369 5074 12369 5074 4 n_40
rlabel m2contact 12369 4642 12369 4642 4 n_248
rlabel m2contact 12321 5986 12321 5986 4 n_336
rlabel m2contact 12273 2890 12273 2890 4 n_184
rlabel m2contact 12249 5074 12249 5074 4 n_317
rlabel m2contact 12129 3082 12129 3082 4 CFlag
rlabel m2contact 12081 2146 12081 2146 4 n_334
rlabel m2contact 12033 2890 12033 2890 4 Op1Sel
rlabel m2contact 12009 6778 12009 6778 4 n_285
rlabel m2contact 11961 2122 11961 2122 4 n_33
rlabel m2contact 11937 2818 11937 2818 4 OpcodeCondIn[4]
rlabel m2contact 11913 4162 11913 4162 4 n_134
rlabel m2contact 11865 6658 11865 6658 4 n_12
rlabel m2contact 11841 3898 11841 3898 4 OpcodeCondIn[3]
rlabel m2contact 11817 3946 11817 3946 4 n_122
rlabel m2contact 11745 3322 11745 3322 4 n_81
rlabel m2contact 11697 6754 11697 6754 4 n_250
rlabel m2contact 11697 6658 11697 6658 4 n_213
rlabel m2contact 11649 1906 11649 1906 4 n_315
rlabel m2contact 11649 6730 11649 6730 4 n_95
rlabel m2contact 11649 4858 11649 4858 4 n_276
rlabel m2contact 11649 2122 11649 2122 4 n_276
rlabel m2contact 11625 3634 11625 3634 4 n_237
rlabel m2contact 11601 6706 11601 6706 4 n_47
rlabel m2contact 11601 2482 11601 2482 4 n_364
rlabel m2contact 11577 4954 11577 4954 4 n_209
rlabel m2contact 11553 2938 11553 2938 4 n_210
rlabel m2contact 11553 4738 11553 4738 4 n_191
rlabel m2contact 11529 4210 11529 4210 4 n_211
rlabel m2contact 11505 5530 11505 5530 4 n_288
rlabel m2contact 11481 6682 11481 6682 4 n_62
rlabel m2contact 11457 3634 11457 3634 4 n_237
rlabel m2contact 11433 4234 11433 4234 4 n_215
rlabel m2contact 11409 2122 11409 2122 4 n_276
rlabel m2contact 11409 4210 11409 4210 4 n_211
rlabel m2contact 11385 5410 11385 5410 4 n_151
rlabel m2contact 11361 1930 11361 1930 4 n_99
rlabel m2contact 11337 6682 11337 6682 4 LrSel
rlabel m2contact 11337 2122 11337 2122 4 LrSel
rlabel m2contact 11313 6682 11313 6682 4 LrSel
rlabel m2contact 11313 5938 11313 5938 4 n_127
rlabel m2contact 11289 2362 11289 2362 4 n_113
rlabel m2contact 11241 2410 11241 2410 4 n_263
rlabel m2contact 11217 2578 11217 2578 4 n_340
rlabel m2contact 11217 5026 11217 5026 4 n_168
rlabel m2contact 11169 4234 11169 4234 4 n_215
rlabel m2contact 11169 4114 11169 4114 4 PcSel[2]
rlabel m2contact 11145 6058 11145 6058 4 state[0]
rlabel m2contact 11097 5026 11097 5026 4 n_257
rlabel m2contact 11097 2986 11097 2986 4 n_257
rlabel m2contact 11073 5938 11073 5938 4 n_127
rlabel m2contact 11073 4642 11073 4642 4 n_248
rlabel m2contact 11049 5362 11049 5362 4 n_85
rlabel m2contact 11049 3298 11049 3298 4 n_84
rlabel m2contact 11025 6058 11025 6058 4 state[0]
rlabel m2contact 11001 6202 11001 6202 4 n_264
rlabel m2contact 10977 5026 10977 5026 4 n_257
rlabel m2contact 10977 3130 10977 3130 4 state[1]
rlabel m2contact 10953 6058 10953 6058 4 state[0]
rlabel m2contact 10929 5458 10929 5458 4 n_150
rlabel m2contact 10905 5698 10905 5698 4 n_66
rlabel m2contact 10881 3730 10881 3730 4 stateSub[1]
rlabel m2contact 10857 2578 10857 2578 4 n_254
rlabel m2contact 10857 4546 10857 4546 4 n_282
rlabel m2contact 10833 4978 10833 4978 4 n_226
rlabel m2contact 10809 4330 10809 4330 4 n_185
rlabel m2contact 10785 5002 10785 5002 4 n_178
rlabel m2contact 10761 2074 10761 2074 4 n_268
rlabel m2contact 10761 4234 10761 4234 4 n_215
rlabel m2contact 10737 4930 10737 4930 4 n_174
rlabel m2contact 10713 3730 10713 3730 4 stateSub[1]
rlabel m2contact 10689 3682 10689 3682 4 n_359
rlabel m2contact 10689 6538 10689 6538 4 stateSub[2]
rlabel m2contact 10665 5026 10665 5026 4 n_301
rlabel m2contact 10665 2362 10665 2362 4 n_301
rlabel m2contact 10641 5026 10641 5026 4 n_301
rlabel m2contact 10641 2410 10641 2410 4 n_322
rlabel m2contact 10617 3994 10617 3994 4 n_302
rlabel m2contact 10617 4762 10617 4762 4 n_251
rlabel m2contact 10593 2458 10593 2458 4 n_217
rlabel m2contact 10569 6514 10569 6514 4 n_374
rlabel m2contact 10569 1930 10569 1930 4 n_374
rlabel m2contact 10545 5458 10545 5458 4 n_150
rlabel m2contact 10521 4762 10521 4762 4 n_177
rlabel m2contact 10521 3994 10521 3994 4 n_177
rlabel m2contact 10497 1930 10497 1930 4 n_374
rlabel m2contact 10497 3226 10497 3226 4 n_53
rlabel m2contact 10473 3130 10473 3130 4 state[1]
rlabel m2contact 10449 5026 10449 5026 4 n_223
rlabel m2contact 10425 5818 10425 5818 4 ImmSel
rlabel m2contact 10401 2818 10401 2818 4 OpcodeCondIn[4]
rlabel m2contact 10377 3994 10377 3994 4 n_177
rlabel m2contact 10377 4714 10377 4714 4 n_190
rlabel m2contact 10329 4162 10329 4162 4 n_134
rlabel m2contact 10305 4906 10305 4906 4 n_117
rlabel m2contact 10281 6538 10281 6538 4 n_152
rlabel m2contact 10257 6658 10257 6658 4 n_213
rlabel m2contact 10257 5818 10257 5818 4 n_212
rlabel m2contact 10233 2410 10233 2410 4 n_322
rlabel m2contact 10209 5218 10209 5218 4 n_175
rlabel m2contact 10161 3682 10161 3682 4 nOE
rlabel m2contact 10137 1954 10137 1954 4 n_91
rlabel m2contact 10137 5194 10137 5194 4 n_198
rlabel m2contact 10113 3994 10113 3994 4 n_319
rlabel m2contact 10089 5194 10089 5194 4 n_356
rlabel m2contact 10065 2770 10065 2770 4 n_189
rlabel m2contact 10041 5218 10041 5218 4 n_92
rlabel m2contact 10041 4714 10041 4714 4 n_190
rlabel m2contact 10017 6490 10017 6490 4 OpcodeCondIn[5]
rlabel m2contact 10017 4738 10017 4738 4 n_191
rlabel m2contact 9993 6634 9993 6634 4 n_60
rlabel m2contact 9945 5626 9945 5626 4 n_124
rlabel m2contact 9945 4954 9945 4954 4 n_209
rlabel m2contact 9921 2986 9921 2986 4 n_257
rlabel m2contact 9921 4210 9921 4210 4 n_211
rlabel m2contact 9897 5626 9897 5626 4 n_41
rlabel m2contact 9873 6634 9873 6634 4 n_257
rlabel m2contact 9873 2986 9873 2986 4 n_257
rlabel m2contact 9849 2770 9849 2770 4 n_158
rlabel m2contact 9825 3130 9825 3130 4 state[1]
rlabel m2contact 9825 3394 9825 3394 4 n_220
rlabel m2contact 9801 6634 9801 6634 4 n_257
rlabel m2contact 9801 4066 9801 4066 4 n_101
rlabel m2contact 9777 3010 9777 3010 4 n_160
rlabel m2contact 9753 2002 9753 2002 4 PcEn
rlabel m2contact 9729 6610 9729 6610 4 n_208
rlabel m2contact 9729 5194 9729 5194 4 n_356
rlabel m2contact 9705 2434 9705 2434 4 n_214
rlabel m2contact 9681 4858 9681 4858 4 n_276
rlabel m2contact 9633 6586 9633 6586 4 n_54
rlabel m2contact 9633 6058 9633 6058 4 state[0]
rlabel m2contact 9633 2002 9633 2002 4 state[0]
rlabel m2contact 9609 1978 9609 1978 4 n_137
rlabel m2contact 9609 3226 9609 3226 4 n_53
rlabel m2contact 9585 4810 9585 4810 4 n_86
rlabel m2contact 9585 3898 9585 3898 4 OpcodeCondIn[3]
rlabel m2contact 9561 3802 9561 3802 4 n_136
rlabel m2contact 9537 5818 9537 5818 4 n_212
rlabel m2contact 9513 4258 9513 4258 4 n_59
rlabel m2contact 9513 5002 9513 5002 4 n_178
rlabel m2contact 9489 2002 9489 2002 4 state[0]
rlabel m2contact 9489 2938 9489 2938 4 n_210
rlabel m2contact 9465 4210 9465 4210 4 n_211
rlabel m2contact 9465 3826 9465 3826 4 n_58
rlabel m2contact 9417 5818 9417 5818 4 n_242
rlabel m2contact 9417 3802 9417 3802 4 n_304
rlabel m2contact 9393 3538 9393 3538 4 stateSub[0]
rlabel m2contact 9369 5698 9369 5698 4 n_66
rlabel m2contact 9345 4258 9345 4258 4 n_238
rlabel m2contact 9273 2026 9273 2026 4 n_280
rlabel m2contact 9273 6562 9273 6562 4 n_120
rlabel m2contact 9225 2050 9225 2050 4 n_103
rlabel m2contact 9225 2650 9225 2650 4 n_119
rlabel m2contact 9177 6538 9177 6538 4 n_152
rlabel m2contact 9177 5770 9177 5770 4 n_253
rlabel m2contact 9153 5410 9153 5410 4 n_151
rlabel m2contact 9129 4330 9129 4330 4 n_185
rlabel m2contact 9105 4858 9105 4858 4 n_276
rlabel m2contact 9081 5506 9081 5506 4 n_289
rlabel m2contact 9057 6514 9057 6514 4 n_374
rlabel m2contact 9057 3538 9057 3538 4 stateSub[0]
rlabel m2contact 9033 6466 9033 6466 4 n_368
rlabel m2contact 9033 3730 9033 3730 4 stateSub[1]
rlabel m2contact 8985 5602 8985 5602 4 n_28
rlabel m2contact 8961 6490 8961 6490 4 OpcodeCondIn[5]
rlabel m2contact 8961 6466 8961 6466 4 n_19
rlabel m2contact 8961 2914 8961 2914 4 n_19
rlabel m2contact 8937 6466 8937 6466 4 n_19
rlabel m2contact 8937 4474 8937 4474 4 n_260
rlabel m2contact 8889 6466 8889 6466 4 LrEn
rlabel m2contact 8889 4522 8889 4522 4 n_286
rlabel m2contact 8865 5506 8865 5506 4 n_289
rlabel m2contact 8841 2074 8841 2074 4 n_268
rlabel m2contact 8817 2242 8817 2242 4 n_65
rlabel m2contact 8793 6466 8793 6466 4 LrEn
rlabel m2contact 8769 4426 8769 4426 4 n_35
rlabel m2contact 8745 2098 8745 2098 4 n_345
rlabel m2contact 8721 6442 8721 6442 4 n_197
rlabel m2contact 8697 6418 8697 6418 4 n_149
rlabel m2contact 8673 2122 8673 2122 4 LrSel
rlabel m2contact 8673 6058 8673 6058 4 state[0]
rlabel m2contact 8625 2122 8625 2122 4 AluEn
rlabel m2contact 8577 2122 8577 2122 4 AluEn
rlabel m2contact 8577 3658 8577 3658 4 n_205
rlabel m2contact 8553 2482 8553 2482 4 n_364
rlabel m2contact 8529 2146 8529 2146 4 n_334
rlabel m2contact 8529 5458 8529 5458 4 n_150
rlabel m2contact 8505 4234 8505 4234 4 n_215
rlabel m2contact 8457 6394 8457 6394 4 n_163
rlabel m2contact 8457 6370 8457 6370 4 n_206
rlabel m2contact 8433 2434 8433 2434 4 n_214
rlabel m2contact 8433 4234 8433 4234 4 n_116
rlabel m2contact 8409 6298 8409 6298 4 n_162
rlabel m2contact 8409 3658 8409 3658 4 n_205
rlabel m2contact 8361 6346 8361 6346 4 n_133
rlabel m2contact 8361 6298 8361 6298 4 n_324
rlabel m2contact 8337 2170 8337 2170 4 Flags[2]
rlabel m2contact 8337 5410 8337 5410 4 n_151
rlabel m2contact 8313 2194 8313 2194 4 n_327
rlabel m2contact 8313 2458 8313 2458 4 n_217
rlabel m2contact 8289 5458 8289 5458 4 n_150
rlabel m2contact 8241 6322 8241 6322 4 n_176
rlabel m2contact 8241 5554 8241 5554 4 n_51
rlabel m2contact 8217 6058 8217 6058 4 state[0]
rlabel m2contact 8217 4450 8217 4450 4 n_235
rlabel m2contact 8193 5482 8193 5482 4 n_147
rlabel m2contact 8145 5482 8145 5482 4 n_370
rlabel m2contact 8145 2914 8145 2914 4 n_19
rlabel m2contact 8121 5554 8121 5554 4 n_350
rlabel m2contact 8097 6298 8097 6298 4 n_324
rlabel m2contact 8097 2818 8097 2818 4 OpcodeCondIn[4]
rlabel m2contact 8073 6274 8073 6274 4 n_293
rlabel m2contact 8025 6250 8025 6250 4 n_83
rlabel m2contact 8025 4690 8025 4690 4 OpcodeCondIn[2]
rlabel m2contact 8001 2218 8001 2218 4 n_484
rlabel m2contact 8001 3298 8001 3298 4 n_84
rlabel m2contact 7977 6202 7977 6202 4 n_264
rlabel m2contact 7977 2242 7977 2242 4 n_65
rlabel m2contact 7929 6226 7929 6226 4 n_273
rlabel m2contact 7929 6202 7929 6202 4 n_3
rlabel m2contact 7929 2242 7929 2242 4 n_3
rlabel m2contact 7905 2242 7905 2242 4 n_3
rlabel m2contact 7905 6058 7905 6058 4 state[0]
rlabel m2contact 7881 4282 7881 4282 4 n_272
rlabel m2contact 7857 3706 7857 3706 4 nWait
rlabel m2contact 7833 2290 7833 2290 4 n_31
rlabel m2contact 7809 2266 7809 2266 4 n_52
rlabel m2contact 7797 6058 7797 6058 4 state[0]
rlabel m2contact 7797 2290 7797 2290 4 state[0]
rlabel m2contact 7785 6130 7785 6130 4 n_6
rlabel m2contact 7761 2290 7761 2290 4 state[0]
rlabel m2contact 7761 3778 7761 3778 4 n_30
rlabel m2contact 7713 6130 7713 6130 4 n_10
rlabel m2contact 7689 6202 7689 6202 4 n_3
rlabel m2contact 7689 3562 7689 3562 4 n_321
rlabel m2contact 7665 4858 7665 4858 4 n_276
rlabel m2contact 7641 3562 7641 3562 4 n_307
rlabel m2contact 7617 6178 7617 6178 4 n_312
rlabel m2contact 7593 2314 7593 2314 4 n_131
rlabel m2contact 7593 4042 7593 4042 4 n_313
rlabel m2contact 7569 6154 7569 6154 4 n_164
rlabel m2contact 7569 3898 7569 3898 4 OpcodeCondIn[3]
rlabel m2contact 7545 4210 7545 4210 4 n_211
rlabel m2contact 7521 2338 7521 2338 4 n_73
rlabel m2contact 7497 6130 7497 6130 4 n_10
rlabel m2contact 7473 6106 7473 6106 4 n_72
rlabel m2contact 7473 2386 7473 2386 4 n_487
rlabel m2contact 7449 2722 7449 2722 4 StatusReg[2]
rlabel m2contact 7425 2410 7425 2410 4 n_322
rlabel m2contact 7401 2386 7401 2386 4 ALE
rlabel m2contact 7401 5242 7401 5242 4 n_88
rlabel m2contact 7377 2362 7377 2362 4 n_301
rlabel m2contact 7377 2458 7377 2458 4 n_217
rlabel m2contact 7329 2386 7329 2386 4 ALE
rlabel m2contact 7281 6082 7281 6082 4 n_68
rlabel m2contact 7281 5242 7281 5242 4 n_88
rlabel m2contact 7257 5122 7257 5122 4 n_42
rlabel m2contact 7257 4810 7257 4810 4 n_86
rlabel m2contact 7233 4642 7233 4642 4 n_248
rlabel m2contact 7209 6058 7209 6058 4 state[0]
rlabel m2contact 7209 6034 7209 6034 4 AluWe
rlabel m2contact 7185 2410 7185 2410 4 n_322
rlabel m2contact 7161 6010 7161 6010 4 n_292
rlabel m2contact 7161 5986 7161 5986 4 n_336
rlabel m2contact 7113 2482 7113 2482 4 n_364
rlabel m2contact 7113 3106 7113 3106 4 n_294
rlabel m2contact 7065 5962 7065 5962 4 RwSel[0]
rlabel m2contact 7065 2482 7065 2482 4 SysBus[1]
rlabel m2contact 7041 5938 7041 5938 4 n_127
rlabel m2contact 7017 5914 7017 5914 4 n_296
rlabel m2contact 6993 5890 6993 5890 4 n_314
rlabel m2contact 6993 2434 6993 2434 4 n_214
rlabel m2contact 6969 2458 6969 2458 4 n_217
rlabel m2contact 6945 5866 6945 5866 4 n_352
rlabel m2contact 6945 4858 6945 4858 4 n_276
rlabel m2contact 6921 2482 6921 2482 4 SysBus[1]
rlabel m2contact 6897 5290 6897 5290 4 n_351
rlabel m2contact 6873 5530 6873 5530 4 n_288
rlabel m2contact 6849 5842 6849 5842 4 n_277
rlabel m2contact 6849 4426 6849 4426 4 n_35
rlabel m2contact 6825 4858 6825 4858 4 n_276
rlabel m2contact 6801 5506 6801 5506 4 n_289
rlabel m2contact 6777 5818 6777 5818 4 n_242
rlabel m2contact 6729 2506 6729 2506 4 n_362
rlabel m2contact 6705 2554 6705 2554 4 n_89
rlabel m2contact 6681 2530 6681 2530 4 n_354
rlabel m2contact 6657 2554 6657 2554 4 LrWe
rlabel m2contact 6633 2554 6633 2554 4 LrWe
rlabel m2contact 6585 2578 6585 2578 4 n_254
rlabel m2contact 6561 5794 6561 5794 4 n_252
rlabel m2contact 6537 5770 6537 5770 4 n_253
rlabel m2contact 6489 2602 6489 2602 4 n_114
rlabel m2contact 6465 5746 6465 5746 4 n_78
rlabel m2contact 6441 5722 6441 5722 4 n_76
rlabel m2contact 6441 4930 6441 4930 4 n_174
rlabel m2contact 6417 3658 6417 3658 4 n_205
rlabel m2contact 6393 4306 6393 4306 4 n_153
rlabel m2contact 6369 2626 6369 2626 4 n_135
rlabel m2contact 6369 5722 6369 5722 4 OpcodeCondIn[4]
rlabel m2contact 6369 2818 6369 2818 4 OpcodeCondIn[4]
rlabel m2contact 6345 5722 6345 5722 4 OpcodeCondIn[4]
rlabel m2contact 6345 3514 6345 3514 4 n_239
rlabel m2contact 6321 2650 6321 2650 4 n_119
rlabel m2contact 6321 3466 6321 3466 4 n_146
rlabel m2contact 6273 3922 6273 3922 4 n_34
rlabel m2contact 6249 3226 6249 3226 4 n_53
rlabel m2contact 6225 5698 6225 5698 4 n_66
rlabel m2contact 6225 5674 6225 5674 4 n_182
rlabel m2contact 6201 3922 6201 3922 4 n_241
rlabel m2contact 6153 2674 6153 2674 4 n_100
rlabel m2contact 6105 2698 6105 2698 4 n_202
rlabel m2contact 6105 4570 6105 4570 4 n_310
rlabel m2contact 6057 5650 6057 5650 4 n_221
rlabel m2contact 6057 2770 6057 2770 4 n_158
rlabel m2contact 6009 2770 6009 2770 4 SysBus[2]
rlabel m2contact 6009 3010 6009 3010 4 n_160
rlabel m2contact 5985 5458 5985 5458 4 n_150
rlabel m2contact 5937 5626 5937 5626 4 n_41
rlabel m2contact 5913 5002 5913 5002 4 n_178
rlabel m2contact 5889 4642 5889 4642 4 n_248
rlabel m2contact 5865 2722 5865 2722 4 StatusReg[2]
rlabel m2contact 5865 2962 5865 2962 4 n_159
rlabel m2contact 5817 2746 5817 2746 4 n_485
rlabel m2contact 5817 5002 5817 5002 4 n_94
rlabel m2contact 5793 5602 5793 5602 4 n_28
rlabel m2contact 5769 5578 5769 5578 4 n_49
rlabel m2contact 5697 3418 5697 3418 4 n_255
rlabel m2contact 5649 3874 5649 3874 4 n_194
rlabel m2contact 5601 5554 5601 5554 4 n_350
rlabel m2contact 5577 2770 5577 2770 4 SysBus[2]
rlabel m2contact 5553 5290 5553 5290 4 n_351
rlabel m2contact 5505 5290 5505 5290 4 n_290
rlabel m2contact 5481 5530 5481 5530 4 n_288
rlabel m2contact 5457 5506 5457 5506 4 n_289
rlabel m2contact 5457 5482 5457 5482 4 n_370
rlabel m2contact 5433 5458 5433 5458 4 n_150
rlabel m2contact 5409 3730 5409 3730 4 stateSub[1]
rlabel m2contact 5361 5434 5361 5434 4 n_22
rlabel m2contact 5337 2794 5337 2794 4 n_40
rlabel m2contact 5337 3730 5337 3730 4 stateSub[1]
rlabel m2contact 5313 2818 5313 2818 4 OpcodeCondIn[4]
rlabel m2contact 5313 3538 5313 3538 4 stateSub[0]
rlabel m2contact 5289 2842 5289 2842 4 n_39
rlabel m2contact 5265 2866 5265 2866 4 n_14
rlabel m2contact 5241 2890 5241 2890 4 Op1Sel
rlabel m2contact 5241 3610 5241 3610 4 OpcodeCondIn[7]
rlabel m2contact 5217 4138 5217 4138 4 n_13
rlabel m2contact 5193 4738 5193 4738 4 n_191
rlabel m2contact 5169 4018 5169 4018 4 n_271
rlabel m2contact 5145 3946 5145 3946 4 n_122
rlabel m2contact 5097 5098 5097 5098 4 OpcodeCondIn[6]
rlabel m2contact 5097 3298 5097 3298 4 n_84
rlabel m2contact 5049 3826 5049 3826 4 n_58
rlabel m2contact 5025 5386 5025 5386 4 n_121
rlabel m2contact 4977 3610 4977 3610 4 OpcodeCondIn[7]
rlabel m2contact 4929 3946 4929 3946 4 n_201
rlabel m2contact 4905 5410 4905 5410 4 n_151
rlabel m2contact 4905 5386 4905 5386 4 n_210
rlabel m2contact 4905 2938 4905 2938 4 n_210
rlabel m2contact 4881 5386 4881 5386 4 n_210
rlabel m2contact 4881 3514 4881 3514 4 n_239
rlabel m2contact 4857 2914 4857 2914 4 n_19
rlabel m2contact 4809 5362 4809 5362 4 n_85
rlabel m2contact 4809 3034 4809 3034 4 n_348
rlabel m2contact 4785 5338 4785 5338 4 n_93
rlabel m2contact 4761 5314 4761 5314 4 n_26
rlabel m2contact 4761 3034 4761 3034 4 n_303
rlabel m2contact 4737 5290 4737 5290 4 n_290
rlabel m2contact 4713 5266 4713 5266 4 n_156
rlabel m2contact 4689 5242 4689 5242 4 n_88
rlabel m2contact 4641 4090 4641 4090 4 n_27
rlabel m2contact 4617 5218 4617 5218 4 n_92
rlabel m2contact 4593 5194 4593 5194 4 n_356
rlabel m2contact 4545 5170 4545 5170 4 n_80
rlabel m2contact 4521 5146 4521 5146 4 n_79
rlabel m2contact 4521 2986 4521 2986 4 n_257
rlabel m2contact 4449 5122 4449 5122 4 n_42
rlabel m2contact 4425 2938 4425 2938 4 n_210
rlabel m2contact 4377 5098 4377 5098 4 OpcodeCondIn[6]
rlabel m2contact 4353 2962 4353 2962 4 n_159
rlabel m2contact 4353 3610 4353 3610 4 OpcodeCondIn[7]
rlabel m2contact 4329 2986 4329 2986 4 n_257
rlabel m2contact 4305 3010 4305 3010 4 n_160
rlabel m2contact 4281 3034 4281 3034 4 n_303
rlabel m2contact 4257 5074 4257 5074 4 n_317
rlabel m2contact 4233 5050 4233 5050 4 n_261
rlabel m2contact 4209 5026 4209 5026 4 n_223
rlabel m2contact 4209 3538 4209 3538 4 stateSub[0]
rlabel m2contact 4161 3058 4161 3058 4 n_155
rlabel m2contact 4137 5002 4137 5002 4 n_94
rlabel m2contact 4113 3082 4113 3082 4 CFlag
rlabel m2contact 4113 4330 4113 4330 4 n_185
rlabel m2contact 4089 3106 4089 3106 4 n_294
rlabel m2contact 4065 4978 4065 4978 4 n_226
rlabel m2contact 4017 4954 4017 4954 4 n_209
rlabel m2contact 3993 4930 3993 4930 4 n_174
rlabel m2contact 3945 3130 3945 3130 4 state[1]
rlabel m2contact 3921 4258 3921 4258 4 n_238
rlabel m2contact 3897 4858 3897 4858 4 n_276
rlabel m2contact 3873 4882 3873 4882 4 n_171
rlabel m2contact 3801 4330 3801 4330 4 n_185
rlabel m2contact 3753 4906 3753 4906 4 n_117
rlabel m2contact 3705 4882 3705 4882 4 n_171
rlabel m2contact 3681 3274 3681 3274 4 n_170
rlabel m2contact 3657 4858 3657 4858 4 n_276
rlabel m2contact 3609 4834 3609 4834 4 n_318
rlabel m2contact 3585 4810 3585 4810 4 n_86
rlabel m2contact 3561 4786 3561 4786 4 n_275
rlabel m2contact 3513 3154 3513 3154 4 n_96
rlabel m2contact 3465 3178 3465 3178 4 n_23
rlabel m2contact 3441 3202 3441 3202 4 n_45
rlabel m2contact 3393 4762 3393 4762 4 n_177
rlabel m2contact 3393 3514 3393 3514 4 n_239
rlabel m2contact 3369 4738 3369 4738 4 n_191
rlabel m2contact 3345 4714 3345 4714 4 n_190
rlabel m2contact 3297 3226 3297 3226 4 n_53
rlabel m2contact 3297 3394 3297 3394 4 n_220
rlabel m2contact 3273 4690 3273 4690 4 OpcodeCondIn[2]
rlabel m2contact 3249 3898 3249 3898 4 OpcodeCondIn[3]
rlabel m2contact 3225 3250 3225 3250 4 n_199
rlabel m2contact 3201 4666 3201 4666 4 n_249
rlabel m2contact 3201 3898 3201 3898 4 OpcodeCondIn[3]
rlabel m2contact 3177 4642 3177 4642 4 n_248
rlabel m2contact 3177 3274 3177 3274 4 n_170
rlabel m2contact 3153 4618 3153 4618 4 n_207
rlabel m2contact 3105 4594 3105 4594 4 AluOR[1]
rlabel m2contact 3105 3298 3105 3298 4 n_84
rlabel m2contact 3081 4570 3081 4570 4 n_310
rlabel m2contact 3081 3322 3081 3322 4 n_81
rlabel m2contact 3057 4546 3057 4546 4 n_282
rlabel m2contact 3033 4522 3033 4522 4 n_286
rlabel m2contact 3033 4498 3033 4498 4 Op2Sel[1]
rlabel m2contact 3009 3346 3009 3346 4 n_284
rlabel m2contact 2985 4474 2985 4474 4 n_260
rlabel m2contact 2961 3370 2961 3370 4 n_183
rlabel m2contact 2961 4162 2961 4162 4 n_134
rlabel m2contact 2937 4450 2937 4450 4 n_235
rlabel m2contact 2889 4426 2889 4426 4 n_35
rlabel m2contact 2865 4402 2865 4402 4 OpcodeCondIn[1]
rlabel m2contact 2841 4138 2841 4138 4 n_13
rlabel m2contact 2793 4378 2793 4378 4 n_186
rlabel m2contact 2793 4354 2793 4354 4 WdSel
rlabel m2contact 2769 3610 2769 3610 4 OpcodeCondIn[7]
rlabel m2contact 2745 4330 2745 4330 4 n_185
rlabel m2contact 2745 3394 2745 3394 4 n_220
rlabel m2contact 2721 4306 2721 4306 4 n_153
rlabel m2contact 2721 3418 2721 3418 4 n_255
rlabel m2contact 2673 4282 2673 4282 4 n_272
rlabel m2contact 2673 3442 2673 3442 4 n_243
rlabel m2contact 2649 3634 2649 3634 4 n_237
rlabel m2contact 2625 4258 2625 4258 4 n_238
rlabel m2contact 2625 3466 2625 3466 4 n_146
rlabel m2contact 2601 3490 2601 3490 4 n_169
rlabel m2contact 2577 4234 2577 4234 4 n_116
rlabel m2contact 2553 4210 2553 4210 4 n_211
rlabel m2contact 2553 4186 2553 4186 4 n_44
rlabel m2contact 2529 3514 2529 3514 4 n_239
rlabel m2contact 2529 3586 2529 3586 4 n_115
rlabel m2contact 2481 4162 2481 4162 4 n_134
rlabel m2contact 2457 3898 2457 3898 4 OpcodeCondIn[3]
rlabel m2contact 2433 3610 2433 3610 4 OpcodeCondIn[7]
rlabel m2contact 2361 4138 2361 4138 4 n_13
rlabel m2contact 2361 3538 2361 3538 4 stateSub[0]
rlabel m2contact 2313 3778 2313 3778 4 n_30
rlabel m2contact 2265 4114 2265 4114 4 PcSel[2]
rlabel m2contact 2217 4090 2217 4090 4 n_27
rlabel m2contact 2193 4066 2193 4066 4 n_101
rlabel m2contact 2121 4042 2121 4042 4 n_313
rlabel m2contact 2073 4018 2073 4018 4 n_271
rlabel m2contact 2001 3994 2001 3994 4 n_319
rlabel m2contact 1953 3802 1953 3802 4 n_304
rlabel m2contact 1905 3562 1905 3562 4 n_307
rlabel m2contact 1881 3802 1881 3802 4 n_246
rlabel m2contact 1857 3970 1857 3970 4 n_142
rlabel m2contact 1833 3946 1833 3946 4 n_201
rlabel m2contact 1833 3586 1833 3586 4 n_115
rlabel m2contact 1785 3922 1785 3922 4 n_241
rlabel m2contact 1785 3610 1785 3610 4 OpcodeCondIn[7]
rlabel m2contact 1761 3634 1761 3634 4 n_237
rlabel m2contact 1737 3898 1737 3898 4 OpcodeCondIn[3]
rlabel m2contact 1713 3874 1713 3874 4 n_194
rlabel m2contact 1713 3850 1713 3850 4 nWE
rlabel m2contact 1665 3826 1665 3826 4 n_58
rlabel m2contact 1665 3802 1665 3802 4 n_246
rlabel m2contact 1641 3778 1641 3778 4 n_30
rlabel m2contact 1641 3754 1641 3754 4 n_200
rlabel m2contact 1617 3658 1617 3658 4 n_205
rlabel m2contact 1617 3730 1617 3730 4 stateSub[1]
rlabel metal2 25431 7964 25443 7964 6 StatusRegEn
rlabel metal2 24615 7964 24627 7964 6 StatusReg[3]
rlabel metal2 23799 7964 23811 7964 6 StatusReg[2]
rlabel metal2 22983 7964 22995 7964 6 StatusReg[1]
rlabel metal2 22167 7964 22179 7964 6 StatusReg[0]
rlabel metal2 21351 7964 21363 7964 6 AluEn
rlabel metal2 21327 7964 21339 7964 6 AluWe
rlabel metal2 20511 7964 20523 7964 6 Op2Sel[1]
rlabel metal2 19695 7964 19707 7964 6 Op2Sel[0]
rlabel metal2 18087 7964 18099 7964 6 Op1Sel
rlabel metal2 17991 7964 18003 7964 6 PcEn
rlabel metal2 17247 7964 17259 7964 6 WdSel
rlabel metal2 15639 7964 15651 7964 6 PcWe
rlabel metal2 14823 7964 14835 7964 6 PcSel[2]
rlabel metal2 14799 7964 14811 7964 6 PcSel[1]
rlabel metal2 13983 7964 13995 7964 6 PcSel[0]
rlabel metal2 12363 7964 12375 7964 4 LrEn
rlabel metal2 11535 7964 11547 7964 4 LrWe
rlabel metal2 11319 7964 11331 7964 4 LrSel
rlabel metal2 10431 7964 10443 7964 4 ImmSel
rlabel metal2 9843 7964 9855 7964 4 IrWe
rlabel metal2 9015 7964 9027 7964 4 MemEn
rlabel metal2 7395 7964 7407 7964 4 OpcodeCondIn[7]
rlabel metal2 6567 7964 6579 7964 4 OpcodeCondIn[6]
rlabel metal2 6531 7964 6543 7964 4 OpcodeCondIn[5]
rlabel metal2 5703 7964 5715 7964 4 OpcodeCondIn[4]
rlabel metal2 4083 7964 4095 7964 4 OpcodeCondIn[3]
rlabel metal2 3279 7964 3291 7964 4 OpcodeCondIn[2]
rlabel metal2 2871 7964 2883 7964 4 OpcodeCondIn[1]
rlabel metal2 2319 7964 2331 7964 4 OpcodeCondIn[0]
rlabel metal2 23607 0 23619 0 8 SysBus[3]
rlabel metal2 14019 0 14031 0 8 SysBus[2]
rlabel metal2 7815 0 7827 0 2 SysBus[1]
rlabel metal2 7779 0 7791 0 2 SysBus[0]
rlabel metal2 0 59 0 71 2 nWE
rlabel metal2 0 35 0 47 2 nIRQ
rlabel metal2 0 3700 0 3712 4 nWait
rlabel metal2 0 3676 0 3688 4 nOE
rlabel metal2 0 7821 0 7833 4 ALE
rlabel metal2 0 7797 0 7809 4 nME
rlabel metal2 123 7964 323 7964 5 Vdd!
rlabel metal2 339 7964 351 7964 5 SDO
rlabel metal2 363 7964 375 7964 5 Test
rlabel metal2 387 7964 399 7964 5 Clock
rlabel metal2 411 7964 423 7964 5 nReset
rlabel metal2 123 0 323 0 1 Vdd!
rlabel metal2 339 0 351 0 1 SDI
rlabel metal2 363 0 375 0 1 Test
rlabel metal2 387 0 399 0 1 Clock
rlabel metal2 411 0 423 0 1 nReset
rlabel metal2 26905 539 26905 551 8 RegWe
rlabel metal2 26905 59 26905 71 8 AluOR[0]
rlabel metal2 26905 35 26905 47 8 AluOR[1]
rlabel metal2 26905 11 26905 23 8 ENB
rlabel metal2 26905 6316 26905 6328 6 Rs1Sel[0]
rlabel metal2 26905 4492 26905 4504 6 Rs1Sel[1]
rlabel metal2 26905 1876 26905 1888 6 RwSel[0]
rlabel metal2 26905 1852 26905 1864 6 RwSel[1]
rlabel metal2 26905 7725 26905 7737 6 CFlag
rlabel metal2 26905 7701 26905 7713 6 Flags[3]
rlabel metal2 26905 7677 26905 7689 6 Flags[2]
rlabel metal2 26905 7653 26905 7665 6 Flags[1]
rlabel metal2 26905 7629 26905 7641 6 Flags[0]
rlabel metal2 26547 0 26747 0 1 GND!
rlabel metal2 26547 7964 26747 7964 5 GND!
<< end >>
