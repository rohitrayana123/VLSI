magic
tech c035u
timestamp 1395354352
<< nwell >>
rect 24759 7676 25239 8074
<< pwell >>
rect 24759 7275 25239 7676
<< nohmic >>
rect 24759 8011 24766 8021
rect 25231 8011 25239 8021
<< nsubstratetap >>
rect 24766 8005 25231 8021
<< metal1 >>
rect -1416 8254 21302 8264
rect 21340 8254 25599 8264
rect -1416 8230 230 8240
rect 5620 8230 21470 8240
rect -1416 8206 422 8216
rect 436 8206 3398 8216
rect 6316 8206 21374 8216
rect 21412 8206 25599 8216
rect 13492 8182 21422 8192
rect 21460 8182 25599 8192
rect 14260 8158 21350 8168
rect 21388 8158 25599 8168
rect 16036 8134 21326 8144
rect 21364 8134 25599 8144
rect 16780 8110 21398 8120
rect 21436 8110 25599 8120
rect 18772 8086 21446 8096
rect 21484 8086 25599 8096
rect 24759 8057 25239 8067
rect 24759 8034 25239 8044
rect 24759 8005 24766 8021
rect 25231 8005 25239 8021
rect 24759 7996 25239 8005
rect 11740 7253 11750 7263
rect 14956 7253 15614 7263
rect 22828 7253 23702 7263
rect 11620 7229 11846 7239
rect 14764 7229 15398 7239
rect 15412 7229 19238 7239
rect 19252 7229 20702 7239
rect 20716 7229 22814 7239
rect 22828 7229 24614 7239
rect 11140 7205 11798 7215
rect 12484 7205 14750 7215
rect 14908 7205 20390 7215
rect 10516 7181 11126 7191
rect 11356 7181 17270 7191
rect 10468 7157 17054 7167
rect 17068 7157 18422 7167
rect 10420 7133 23726 7143
rect 23740 7133 24470 7143
rect 10156 7109 15806 7119
rect 15820 7109 20294 7119
rect 20308 7109 24062 7119
rect 10156 7085 21782 7095
rect 9532 7061 19838 7071
rect 9220 7037 16454 7047
rect 9052 7013 18110 7023
rect 18124 7013 20462 7023
rect 8860 6989 18710 6999
rect 8812 6965 21302 6975
rect 8764 6941 9038 6951
rect 9148 6941 15254 6951
rect 15268 6941 22358 6951
rect 22372 6941 22838 6951
rect 8692 6917 9302 6927
rect 9532 6917 18254 6927
rect 8668 6893 19334 6903
rect 8452 6869 21398 6879
rect 8404 6845 18326 6855
rect 8332 6821 10118 6831
rect 10132 6821 10982 6831
rect 10996 6821 17462 6831
rect 17476 6821 18134 6831
rect 8308 6797 9182 6807
rect 9196 6797 15446 6807
rect 15460 6797 19310 6807
rect 8308 6773 21710 6783
rect 8260 6749 8438 6759
rect 8500 6749 13598 6759
rect 14428 6749 17582 6759
rect 8212 6725 18398 6735
rect 8140 6701 8174 6711
rect 8236 6701 9686 6711
rect 9700 6701 13838 6711
rect 13852 6701 14510 6711
rect 14524 6701 22382 6711
rect 22396 6701 24014 6711
rect 7996 6677 21206 6687
rect 7948 6653 21230 6663
rect 24460 6653 24662 6663
rect 7900 6629 12470 6639
rect 12484 6629 24446 6639
rect 7804 6605 11006 6615
rect 11188 6605 19046 6615
rect 19060 6605 20990 6615
rect 7732 6581 18686 6591
rect 7636 6557 9086 6567
rect 9100 6557 18350 6567
rect 7564 6533 9566 6543
rect 9580 6533 17798 6543
rect 7396 6509 17390 6519
rect 7372 6485 9326 6495
rect 9484 6485 19934 6495
rect 7324 6461 11990 6471
rect 12004 6461 20294 6471
rect 20308 6461 22118 6471
rect 22132 6461 23486 6471
rect 7228 6437 14894 6447
rect 14908 6437 15494 6447
rect 7180 6413 7694 6423
rect 7708 6413 17294 6423
rect 17308 6413 20918 6423
rect 7036 6389 16694 6399
rect 6676 6365 21902 6375
rect 6460 6341 21494 6351
rect 6316 6317 6326 6327
rect 6388 6317 7238 6327
rect 7252 6317 7598 6327
rect 7612 6317 12062 6327
rect 12076 6317 15734 6327
rect 15748 6317 19094 6327
rect 19108 6317 22790 6327
rect 22804 6317 23198 6327
rect 6220 6293 8198 6303
rect 8212 6293 12398 6303
rect 12412 6293 17798 6303
rect 17812 6293 18326 6303
rect 6172 6269 20702 6279
rect 6124 6245 6758 6255
rect 6772 6245 9542 6255
rect 9556 6245 10550 6255
rect 10564 6245 15014 6255
rect 15028 6245 20342 6255
rect 5764 6221 21614 6231
rect 5404 6197 14918 6207
rect 5404 6173 12494 6183
rect 14188 6173 18878 6183
rect 5380 6149 7166 6159
rect 7180 6149 8678 6159
rect 8692 6149 22622 6159
rect 22636 6149 23318 6159
rect 5380 6125 15278 6135
rect 5356 6101 21590 6111
rect 21604 6101 25262 6111
rect 5308 6077 22910 6087
rect 5284 6053 5942 6063
rect 5956 6053 23078 6063
rect 5284 6029 17342 6039
rect 5236 6005 5918 6015
rect 5932 6005 21974 6015
rect 5188 5981 8726 5991
rect 8740 5981 14198 5991
rect 14380 5981 15158 5991
rect 5068 5957 22886 5967
rect 22900 5957 24398 5967
rect 5020 5933 14126 5943
rect 14140 5933 16694 5943
rect 21892 5933 23606 5943
rect 4972 5909 21014 5919
rect 21028 5909 21878 5919
rect 4972 5885 6806 5895
rect 6964 5885 11462 5895
rect 11476 5885 15230 5895
rect 18676 5885 18758 5895
rect 19396 5885 19466 5895
rect 20236 5885 20270 5895
rect 22084 5885 22574 5895
rect 4924 5861 5174 5871
rect 5188 5861 5990 5871
rect 6004 5861 18542 5871
rect 18556 5861 20654 5871
rect 20668 5861 22070 5871
rect 4900 5837 18038 5847
rect 18052 5837 22454 5847
rect 22468 5837 23390 5847
rect 23404 5837 23678 5847
rect 4900 5813 7430 5823
rect 7492 5813 9062 5823
rect 9076 5813 12326 5823
rect 12340 5813 14774 5823
rect 14788 5813 23558 5823
rect 4828 5789 22598 5799
rect 22612 5789 25238 5799
rect 4684 5765 13646 5775
rect 13660 5765 19958 5775
rect 19972 5765 20222 5775
rect 21868 5765 21914 5775
rect 22420 5765 24110 5775
rect 4492 5741 23318 5751
rect 4492 5717 22958 5727
rect 4420 5693 4718 5703
rect 4732 5693 9374 5703
rect 9388 5693 10190 5703
rect 10204 5693 10478 5703
rect 10492 5693 12206 5703
rect 12220 5693 17438 5703
rect 17452 5693 17918 5703
rect 17932 5693 18134 5703
rect 18148 5693 18230 5703
rect 18244 5693 19142 5703
rect 19156 5693 24374 5703
rect 24388 5693 24398 5703
rect 24412 5693 24686 5703
rect 24700 5693 25118 5703
rect 4324 5669 21854 5679
rect 21868 5669 22526 5679
rect 4228 5645 5246 5655
rect 5260 5645 21950 5655
rect 22324 5645 22670 5655
rect 4204 5621 13190 5631
rect 13468 5621 24734 5631
rect 4180 5597 4190 5607
rect 4276 5597 8654 5607
rect 8668 5597 17006 5607
rect 18628 5597 23030 5607
rect 23044 5597 24422 5607
rect 4084 5573 14378 5583
rect 14392 5573 17678 5583
rect 18532 5573 22406 5583
rect 4036 5549 14990 5559
rect 15004 5549 22310 5559
rect 3820 5525 21134 5535
rect 3796 5501 5726 5511
rect 5740 5501 8942 5511
rect 8956 5501 15134 5511
rect 15148 5501 23990 5511
rect 3772 5477 10166 5487
rect 10324 5477 11990 5487
rect 12844 5477 20750 5487
rect 3700 5453 5678 5463
rect 5692 5453 8870 5463
rect 8884 5453 10070 5463
rect 10084 5453 14534 5463
rect 14548 5453 19262 5463
rect 19276 5453 24086 5463
rect 3676 5429 8846 5439
rect 8860 5429 13886 5439
rect 13900 5429 16142 5439
rect 16156 5429 19886 5439
rect 3364 5405 18662 5415
rect 18676 5405 20534 5415
rect 3340 5381 11726 5391
rect 11740 5381 17966 5391
rect 17980 5381 18158 5391
rect 18172 5381 18566 5391
rect 18580 5381 19190 5391
rect 19204 5381 19382 5391
rect 19396 5381 22262 5391
rect 22276 5381 22334 5391
rect 22348 5381 23150 5391
rect 23164 5381 25166 5391
rect 3220 5357 8366 5367
rect 8476 5357 13598 5367
rect 13612 5357 15614 5367
rect 17908 5357 21326 5367
rect 23356 5357 23534 5367
rect 3100 5333 11150 5343
rect 11164 5333 23342 5343
rect 3028 5309 3062 5319
rect 3148 5309 9806 5319
rect 9916 5309 22766 5319
rect 3004 5285 17750 5295
rect 17764 5285 20630 5295
rect 2980 5261 12110 5271
rect 12700 5261 21686 5271
rect 2908 5237 20174 5247
rect 2788 5213 11582 5223
rect 11956 5213 18734 5223
rect 2740 5189 10322 5199
rect 10336 5189 15758 5199
rect 17044 5189 17102 5199
rect 17860 5189 19214 5199
rect 20380 5189 20630 5199
rect 2692 5165 7694 5175
rect 7708 5165 17030 5175
rect 17500 5165 23366 5175
rect 2668 5141 9398 5151
rect 9460 5141 20822 5151
rect 2620 5117 5822 5127
rect 6076 5117 11954 5127
rect 12460 5117 13334 5127
rect 13420 5117 16310 5127
rect 17332 5117 18806 5127
rect 18820 5117 22022 5127
rect 2620 5093 21278 5103
rect 2572 5069 9614 5079
rect 9628 5069 24302 5079
rect 2548 5045 3518 5055
rect 3532 5045 10958 5055
rect 10972 5045 11246 5055
rect 11260 5045 12350 5055
rect 12364 5045 15926 5055
rect 15940 5045 24518 5055
rect 2452 5021 6206 5031
rect 6268 5021 21914 5031
rect 2404 4997 4622 5007
rect 4636 4997 12542 5007
rect 12556 4997 20438 5007
rect 2308 4973 3302 4983
rect 3316 4973 4646 4983
rect 4660 4973 11918 4983
rect 12292 4973 21038 4983
rect 2284 4949 4862 4959
rect 4876 4949 7622 4959
rect 7636 4949 7934 4959
rect 7948 4949 8126 4959
rect 8140 4949 10286 4959
rect 10300 4949 11678 4959
rect 11692 4949 12110 4959
rect 12124 4949 14942 4959
rect 14956 4949 15830 4959
rect 15844 4949 19118 4959
rect 19132 4949 20870 4959
rect 2284 4925 16910 4935
rect 17260 4925 17534 4935
rect 17716 4925 23438 4935
rect 2188 4901 20726 4911
rect 21076 4901 21410 4911
rect 21820 4901 21830 4911
rect 2116 4877 5558 4887
rect 5572 4877 10670 4887
rect 10732 4877 25598 4887
rect 2092 4853 2510 4863
rect 2524 4853 4814 4863
rect 4828 4853 5966 4863
rect 5980 4853 15518 4863
rect 15532 4853 16478 4863
rect 16492 4853 20414 4863
rect 20428 4853 21470 4863
rect 21484 4853 21806 4863
rect 21820 4853 24494 4863
rect 2068 4829 6014 4839
rect 6028 4829 6350 4839
rect 6364 4829 21062 4839
rect 1996 4805 4742 4815
rect 4756 4805 12662 4815
rect 12676 4805 21470 4815
rect 21484 4805 23582 4815
rect 1948 4781 2030 4791
rect 2044 4781 14678 4791
rect 14692 4781 18062 4791
rect 18076 4781 20486 4791
rect 20500 4781 22274 4791
rect 1852 4757 6422 4767
rect 6436 4757 8150 4767
rect 8164 4757 15134 4767
rect 15196 4757 15290 4767
rect 16036 4757 16070 4767
rect 17212 4757 18614 4767
rect 18988 4757 21758 4767
rect 23140 4757 23246 4767
rect 23308 4757 23654 4767
rect 23668 4757 25214 4767
rect 1804 4733 3974 4743
rect 3988 4733 6398 4743
rect 6412 4733 15182 4743
rect 15196 4733 16022 4743
rect 16396 4733 16430 4743
rect 16636 4733 24494 4743
rect 1732 4709 3110 4719
rect 3196 4709 19430 4719
rect 19444 4709 20798 4719
rect 23020 4709 23654 4719
rect 1708 4685 3446 4695
rect 3556 4685 4574 4695
rect 4588 4685 8174 4695
rect 8188 4685 11750 4695
rect 11764 4685 18854 4695
rect 18964 4685 19442 4695
rect 19924 4685 20018 4695
rect 20260 4685 20606 4695
rect 20692 4685 20834 4695
rect 22876 4685 23270 4695
rect 23428 4685 23630 4695
rect 1684 4661 1694 4671
rect 1708 4661 2462 4671
rect 2476 4661 2582 4671
rect 2596 4661 4214 4671
rect 4228 4661 4382 4671
rect 4396 4661 7574 4671
rect 7588 4661 11606 4671
rect 11620 4661 15326 4671
rect 15340 4661 16598 4671
rect 16612 4661 18350 4671
rect 18364 4661 22742 4671
rect 22756 4661 23870 4671
rect 24388 4661 24470 4671
rect 1636 4637 11438 4647
rect 11572 4637 11750 4647
rect 11884 4637 19166 4647
rect 19324 4637 19334 4647
rect 19996 4637 22550 4647
rect 22636 4637 22790 4647
rect 1612 4613 3254 4623
rect 3268 4613 12638 4623
rect 13684 4613 21086 4623
rect 21100 4613 22574 4623
rect 22756 4613 23030 4623
rect 1588 4589 8990 4599
rect 9004 4589 11462 4599
rect 11476 4589 18782 4599
rect 19132 4589 19238 4599
rect 20452 4589 20654 4599
rect 20740 4589 23534 4599
rect 1516 4565 5870 4575
rect 5884 4565 13238 4575
rect 13252 4565 23510 4575
rect 1492 4541 3158 4551
rect 3172 4541 10502 4551
rect 10516 4541 16166 4551
rect 16180 4541 20198 4551
rect 20500 4541 24278 4551
rect 1444 4517 14438 4527
rect 15340 4517 16982 4527
rect 18412 4517 18422 4527
rect 18532 4517 22934 4527
rect 1420 4493 3566 4503
rect 3580 4493 5438 4503
rect 5452 4493 6038 4503
rect 6052 4493 8630 4503
rect 8644 4493 11102 4503
rect 11116 4493 12014 4503
rect 12028 4493 12254 4503
rect 12268 4493 16886 4503
rect 16900 4493 18590 4503
rect 21916 4493 22358 4503
rect 22444 4493 23462 4503
rect 1396 4469 2390 4479
rect 2404 4469 2894 4479
rect 2908 4469 6878 4479
rect 6892 4469 7286 4479
rect 7300 4469 11414 4479
rect 11428 4469 16382 4479
rect 16396 4469 20558 4479
rect 20572 4469 22694 4479
rect 1324 4445 22166 4455
rect 1276 4421 14462 4431
rect 15436 4421 23222 4431
rect 1228 4397 13430 4407
rect 13708 4397 22982 4407
rect 23236 4397 23438 4407
rect 1180 4373 2198 4383
rect 2260 4373 3854 4383
rect 3868 4373 18086 4383
rect 1156 4349 22214 4359
rect 1156 4325 17126 4335
rect 1108 4301 2102 4311
rect 2164 4301 3038 4311
rect 3100 4301 3446 4311
rect 3460 4301 6278 4311
rect 6292 4301 6926 4311
rect 6940 4301 8222 4311
rect 8236 4301 10262 4311
rect 10276 4301 16862 4311
rect 1084 4277 4586 4287
rect 4600 4277 8150 4287
rect 8260 4277 10646 4287
rect 10660 4277 14150 4287
rect 14164 4277 16670 4287
rect 16684 4277 16922 4287
rect 1060 4253 1190 4263
rect 1204 4253 1286 4263
rect 1300 4253 4550 4263
rect 4564 4253 4838 4263
rect 4852 4253 7766 4263
rect 7780 4253 8534 4263
rect 8548 4253 8918 4263
rect 8932 4253 10022 4263
rect 10036 4253 11030 4263
rect 11044 4253 13958 4263
rect 13972 4253 16574 4263
rect 16588 4253 22838 4263
rect 1036 4229 4526 4239
rect 4540 4229 11486 4239
rect 11500 4229 13526 4239
rect 13540 4229 16598 4239
rect 16612 4229 17414 4239
rect 17428 4229 17870 4239
rect 17884 4229 18566 4239
rect 18580 4229 18998 4239
rect 19012 4229 19598 4239
rect 19612 4229 23846 4239
rect 23860 4229 24230 4239
rect 964 4205 1166 4215
rect 1180 4205 6686 4215
rect 6700 4205 6854 4215
rect 6868 4205 12566 4215
rect 12580 4205 17894 4215
rect 17908 4205 23918 4215
rect 916 4181 1862 4191
rect 1924 4181 9110 4191
rect 9172 4181 14630 4191
rect 14644 4181 21974 4191
rect 21988 4181 22094 4191
rect 844 4157 9854 4167
rect 9940 4157 20966 4167
rect 820 4133 10910 4143
rect 11188 4133 14822 4143
rect 15460 4133 18062 4143
rect 18076 4133 18494 4143
rect 20980 4133 21086 4143
rect 772 4109 8006 4119
rect 8092 4109 11822 4119
rect 11932 4109 11954 4119
rect 12028 4109 23174 4119
rect 748 4085 11654 4095
rect 11668 4085 12182 4095
rect 12196 4085 12806 4095
rect 12820 4085 18710 4095
rect 18724 4085 19046 4095
rect 19060 4085 19910 4095
rect 19924 4085 21734 4095
rect 21748 4085 22238 4095
rect 22252 4085 22550 4095
rect 724 4061 2486 4071
rect 2500 4061 4286 4071
rect 4300 4061 4934 4071
rect 4948 4061 5198 4071
rect 5212 4061 5486 4071
rect 5500 4061 6158 4071
rect 6172 4061 17822 4071
rect 17836 4061 20318 4071
rect 20332 4061 22046 4071
rect 22060 4061 23054 4071
rect 652 4037 2222 4047
rect 2236 4037 6494 4047
rect 6580 4037 16982 4047
rect 23068 4037 23198 4047
rect 604 4013 11630 4023
rect 11644 4013 21254 4023
rect 556 3989 18470 3999
rect 21268 3989 21326 3999
rect 532 3965 8966 3975
rect 8980 3965 9734 3975
rect 9748 3965 10094 3975
rect 10108 3965 11486 3975
rect 11500 3965 20150 3975
rect 508 3941 4622 3951
rect 4636 3941 6974 3951
rect 6988 3941 9254 3951
rect 9268 3941 14582 3951
rect 15916 3941 21998 3951
rect 460 3917 2846 3927
rect 2932 3917 9758 3927
rect 9964 3917 16622 3927
rect 16876 3917 17006 3927
rect 18484 3917 20018 3927
rect 20164 3917 20174 3927
rect 412 3893 5126 3903
rect 5140 3893 7430 3903
rect 7444 3893 8750 3903
rect 8812 3893 16358 3903
rect 388 3869 1358 3879
rect 1372 3869 5654 3879
rect 5668 3869 7118 3879
rect 7132 3869 7790 3879
rect 7804 3869 8726 3879
rect 8740 3869 11054 3879
rect 11068 3869 17942 3879
rect 17956 3869 21566 3879
rect 364 3845 878 3855
rect 940 3845 2366 3855
rect 2380 3845 6110 3855
rect 6124 3845 8054 3855
rect 8068 3845 16838 3855
rect 16852 3845 19142 3855
rect 19156 3845 21542 3855
rect 316 3821 12590 3831
rect 13756 3821 16502 3831
rect 21556 3821 21590 3831
rect 292 3797 974 3807
rect 988 3797 7358 3807
rect 7372 3797 9590 3807
rect 9652 3797 9854 3807
rect 9868 3797 12230 3807
rect 12244 3797 12278 3807
rect 12292 3797 14078 3807
rect 14092 3797 14318 3807
rect 14332 3797 22910 3807
rect 244 3773 23414 3783
rect 244 3749 6134 3759
rect 6196 3749 16430 3759
rect 196 3725 19550 3735
rect 172 3701 22646 3711
rect 148 3677 10598 3687
rect 10828 3677 24518 3687
rect -1416 3653 662 3663
rect 724 3653 6230 3663
rect 6244 3653 10214 3663
rect 10228 3653 11078 3663
rect 11092 3653 11390 3663
rect 11404 3653 18590 3663
rect -1416 3629 14030 3639
rect 16324 3629 16718 3639
rect -1416 3605 11294 3615
rect 11716 3605 17102 3615
rect 17116 3605 21446 3615
rect -1416 3581 7550 3591
rect 7684 3581 7838 3591
rect 7852 3581 9350 3591
rect 9412 3581 9566 3591
rect 9676 3581 10238 3591
rect 10300 3581 10322 3591
rect 10420 3581 11510 3591
rect 11956 3581 24662 3591
rect 124 3557 20246 3567
rect 124 3533 3014 3543
rect 3028 3533 11774 3543
rect 12196 3533 16526 3543
rect 16540 3533 16958 3543
rect 16972 3533 22214 3543
rect 148 3509 3470 3519
rect 3484 3509 5294 3519
rect 5308 3509 7982 3519
rect 7996 3509 9302 3519
rect 9316 3509 12086 3519
rect 12100 3509 13550 3519
rect 13564 3509 14006 3519
rect 14020 3509 16286 3519
rect 16300 3509 17774 3519
rect 17788 3509 20798 3519
rect 20812 3509 20894 3519
rect 20908 3509 21374 3519
rect 172 3485 5558 3495
rect 5572 3485 9278 3495
rect 9292 3485 20606 3495
rect 20620 3485 23102 3495
rect 196 3461 22190 3471
rect 340 3437 1046 3447
rect 1108 3437 18446 3447
rect 20908 3437 20990 3447
rect 22204 3437 22274 3447
rect 628 3413 19502 3423
rect 772 3389 974 3399
rect 988 3389 4454 3399
rect 4468 3389 4742 3399
rect 4756 3389 7910 3399
rect 7924 3389 9830 3399
rect 9844 3389 11894 3399
rect 11908 3389 12302 3399
rect 12316 3389 14342 3399
rect 14356 3389 14798 3399
rect 14812 3389 16550 3399
rect 16564 3389 18902 3399
rect 18916 3389 18974 3399
rect 868 3365 22862 3375
rect 964 3341 2006 3351
rect 2020 3341 18014 3351
rect 18028 3341 23774 3351
rect 1084 3317 10886 3327
rect 10900 3317 11366 3327
rect 11380 3317 15350 3327
rect 15364 3317 17222 3327
rect 17236 3317 21134 3327
rect 21148 3317 23582 3327
rect 23596 3317 25070 3327
rect 1540 3293 20678 3303
rect 1756 3269 2630 3279
rect 2644 3269 3062 3279
rect 3076 3269 9422 3279
rect 9436 3269 10382 3279
rect 10396 3269 19574 3279
rect 1780 3245 22766 3255
rect 1828 3221 22478 3231
rect 1900 3197 16046 3207
rect 16060 3197 17990 3207
rect 18004 3197 21158 3207
rect 1948 3173 3638 3183
rect 3652 3173 5150 3183
rect 5164 3173 6086 3183
rect 6100 3173 9878 3183
rect 9892 3173 16814 3183
rect 17236 3173 17270 3183
rect 17788 3173 17966 3183
rect 17980 3173 18110 3183
rect 18460 3173 18542 3183
rect 2044 3149 2534 3159
rect 2548 3149 11558 3159
rect 11572 3149 22934 3159
rect 22948 3149 24206 3159
rect 2068 3125 14222 3135
rect 14236 3125 15206 3135
rect 15220 3125 16742 3135
rect 16756 3125 20006 3135
rect 2332 3101 2774 3111
rect 2884 3101 22262 3111
rect 2356 3077 2438 3087
rect 2452 3077 2558 3087
rect 2572 3077 5774 3087
rect 5788 3077 8606 3087
rect 8620 3077 10358 3087
rect 10372 3077 10766 3087
rect 10780 3077 10862 3087
rect 10876 3077 18878 3087
rect 18892 3077 20834 3087
rect 20848 3077 22718 3087
rect 2380 3053 2390 3063
rect 2500 3053 17630 3063
rect 22732 3053 22886 3063
rect 2404 3029 8414 3039
rect 8620 3029 8654 3039
rect 8716 3029 15038 3039
rect 16732 3029 20510 3039
rect 2692 3005 4766 3015
rect 4780 3005 7382 3015
rect 7396 3005 7502 3015
rect 7516 3005 17078 3015
rect 17092 3005 17654 3015
rect 17668 3005 24566 3015
rect 2956 2981 16238 2991
rect 16828 2981 16922 2991
rect 17644 2981 17678 2991
rect 3004 2957 5846 2967
rect 5860 2957 7334 2967
rect 7348 2957 19070 2967
rect 19084 2957 23462 2967
rect 3124 2933 21182 2943
rect 3220 2909 3494 2919
rect 3508 2909 15110 2919
rect 15124 2909 16454 2919
rect 19084 2909 22142 2919
rect 3268 2885 7886 2895
rect 7900 2885 8102 2895
rect 8116 2885 9710 2895
rect 9724 2885 18830 2895
rect 18844 2885 19790 2895
rect 19804 2885 21662 2895
rect 21676 2885 23966 2895
rect 3340 2861 11750 2871
rect 11764 2861 15290 2871
rect 15304 2861 20774 2871
rect 20788 2861 23126 2871
rect 3604 2837 9758 2847
rect 9988 2837 11006 2847
rect 11020 2837 19622 2847
rect 21196 2837 21206 2847
rect 3724 2813 11246 2823
rect 11308 2813 11846 2823
rect 12220 2813 24326 2823
rect 3916 2789 4166 2799
rect 4252 2789 6398 2799
rect 6412 2789 7094 2799
rect 7108 2789 8558 2799
rect 8572 2789 20582 2799
rect 20596 2789 24182 2799
rect 24196 2789 24710 2799
rect 3988 2765 5894 2775
rect 5980 2765 6206 2775
rect 6268 2765 6710 2775
rect 6724 2765 15398 2775
rect 4012 2741 22958 2751
rect 4036 2717 4190 2727
rect 4204 2717 12590 2727
rect 12604 2717 16190 2727
rect 4108 2693 14702 2703
rect 4132 2669 5414 2679
rect 5596 2669 6302 2679
rect 6316 2669 10694 2679
rect 10708 2669 12518 2679
rect 13780 2669 24542 2679
rect 4348 2645 13382 2655
rect 13396 2645 15638 2655
rect 15652 2645 16358 2655
rect 16372 2645 18758 2655
rect 4564 2621 4586 2631
rect 4684 2621 9494 2631
rect 9748 2621 10022 2631
rect 10108 2621 10118 2631
rect 10324 2621 23246 2631
rect 4948 2597 16214 2607
rect 5068 2573 10646 2583
rect 10660 2573 19022 2583
rect 5140 2549 5174 2559
rect 5236 2549 15278 2559
rect 15292 2549 23630 2559
rect 5716 2525 12398 2535
rect 13396 2525 22502 2535
rect 5788 2501 15470 2511
rect 15484 2501 15542 2511
rect 15556 2501 19358 2511
rect 5908 2477 5942 2487
rect 6028 2477 11582 2487
rect 11596 2477 24590 2487
rect 6148 2453 6278 2463
rect 6388 2453 7718 2463
rect 7732 2453 10790 2463
rect 10804 2453 11414 2463
rect 11428 2453 24158 2463
rect 6244 2429 6422 2439
rect 6484 2429 15062 2439
rect 19036 2429 19094 2439
rect 6532 2405 9950 2415
rect 10012 2405 23822 2415
rect 6604 2381 15854 2391
rect 6628 2357 13574 2367
rect 13972 2357 24638 2367
rect 6796 2333 7094 2343
rect 7156 2333 12734 2343
rect 12748 2333 25190 2343
rect 7252 2309 10238 2319
rect 10252 2309 16262 2319
rect 16276 2309 18038 2319
rect 7276 2285 12374 2295
rect 14356 2285 14378 2295
rect 16276 2285 16406 2295
rect 7852 2261 11822 2271
rect 11836 2261 18926 2271
rect 18940 2261 19466 2271
rect 19480 2261 20102 2271
rect 7924 2237 7934 2247
rect 8044 2237 14294 2247
rect 16420 2237 21350 2247
rect 8788 2213 9998 2223
rect 10012 2213 17558 2223
rect 17572 2213 19166 2223
rect 19180 2213 20270 2223
rect 20284 2213 20942 2223
rect 20956 2213 22670 2223
rect 9244 2189 10598 2199
rect 10612 2189 11198 2199
rect 11212 2189 20918 2199
rect 20932 2189 25142 2199
rect 9268 2165 9326 2175
rect 9508 2165 9686 2175
rect 9796 2165 21110 2175
rect 21364 2165 21410 2175
rect 25276 2165 25599 2175
rect 9340 2141 21830 2151
rect 25252 2141 25599 2151
rect 10060 2117 19406 2127
rect 19420 2117 21614 2127
rect 25228 2117 25599 2127
rect 10540 2093 16070 2103
rect 16084 2093 21398 2103
rect 25204 2093 25599 2103
rect 10564 2069 14870 2079
rect 19420 2069 19442 2079
rect 25180 2069 25599 2079
rect 10588 2045 10838 2055
rect 11092 2045 11150 2055
rect 25156 2045 25599 2055
rect 10372 1212 16166 1222
rect 16780 1212 19454 1222
rect 9916 1188 19694 1198
rect 9580 1164 20078 1174
rect 8932 1140 16262 1150
rect 16756 1140 19190 1150
rect 8884 1116 10022 1126
rect 10036 1116 10118 1126
rect 10132 1116 12830 1126
rect 12844 1116 16478 1126
rect 16492 1116 16958 1126
rect 16972 1116 22574 1126
rect 22588 1116 24734 1126
rect 8644 1092 9206 1102
rect 9220 1092 18494 1102
rect 18508 1092 20462 1102
rect 20476 1092 24806 1102
rect 8572 1068 8942 1078
rect 9052 1068 20690 1078
rect 8524 1044 8894 1054
rect 9004 1044 11270 1054
rect 12436 1044 19814 1054
rect 8500 1020 23174 1030
rect 8356 996 11750 1006
rect 12340 996 18206 1006
rect 8332 972 17846 982
rect 7948 948 8534 958
rect 8548 948 21014 958
rect 6436 924 21278 934
rect 6292 900 19742 910
rect 5980 876 11318 886
rect 12244 876 19262 886
rect 5500 852 7814 862
rect 7828 852 10094 862
rect 10108 852 11678 862
rect 11692 852 20558 862
rect 20572 852 21758 862
rect 21772 852 21998 862
rect 22012 852 23006 862
rect 23020 852 24782 862
rect 5452 828 6542 838
rect 7756 828 11150 838
rect 11212 828 23618 838
rect 5332 804 21230 814
rect 5188 780 23510 790
rect 4996 756 7190 766
rect 7492 756 13982 766
rect 13996 756 17102 766
rect 4660 732 5510 742
rect 5524 732 5606 742
rect 5620 732 14102 742
rect 14116 732 14198 742
rect 14212 732 24758 742
rect 4588 708 23390 718
rect 4504 684 15470 694
rect 15676 684 18110 694
rect 18172 684 24542 694
rect 4444 660 20366 670
rect 4420 636 15974 646
rect 16204 636 19238 646
rect 19684 636 22358 646
rect 23236 634 23254 648
rect 24604 636 24710 646
rect 3628 612 5006 622
rect 5092 612 20894 622
rect 20908 612 24710 622
rect 3412 588 20102 598
rect 3364 564 22646 574
rect 3148 540 7646 550
rect 7660 540 8006 550
rect 8116 540 20582 550
rect 3076 516 20846 526
rect 3028 492 15230 502
rect 15724 492 21662 502
rect 2932 468 16574 478
rect 17752 468 21350 478
rect 2884 444 18830 454
rect 2860 420 12134 430
rect 12988 420 20030 430
rect 2812 396 20822 406
rect 2764 372 10886 382
rect 10900 372 15566 382
rect 16288 372 23270 382
rect 2716 348 14174 358
rect 14824 348 21926 358
rect 2188 324 9350 334
rect 9460 324 10430 334
rect 10732 324 16094 334
rect 2164 300 14222 310
rect 2140 276 11510 286
rect 13804 276 18806 286
rect 1348 252 10454 262
rect 10756 252 18278 262
rect 1228 228 8366 238
rect 8452 228 10430 238
rect 10804 228 11966 238
rect 14020 228 18926 238
rect -1416 204 20630 214
rect -1416 180 230 190
rect 916 178 934 192
rect 1012 180 16670 190
rect -1416 156 7094 166
rect 7456 156 22430 166
rect -1416 132 10838 142
rect 10948 132 16934 142
rect 24724 132 25599 142
rect 2308 108 17762 118
rect 24820 108 25599 118
rect 4180 84 19226 94
rect 24796 84 25599 94
rect 5740 60 24710 70
rect 24772 60 25599 70
rect 9100 36 11906 46
rect 24748 36 25599 46
rect 9964 10 9982 24
rect 10348 12 12854 22
rect 24724 12 25599 22
<< m2contact >>
rect -1430 8252 -1416 8266
rect 21302 8252 21316 8266
rect 21326 8252 21340 8266
rect 25599 8252 25613 8266
rect -1430 8228 -1416 8242
rect 230 8228 244 8242
rect 5606 8228 5620 8242
rect 21470 8228 21484 8242
rect -1430 8204 -1416 8218
rect 422 8204 436 8218
rect 3398 8204 3412 8218
rect 6302 8204 6316 8218
rect 21374 8204 21388 8218
rect 21398 8204 21412 8218
rect 25599 8204 25613 8218
rect 13478 8180 13492 8194
rect 21422 8180 21436 8194
rect 21446 8180 21460 8194
rect 25599 8180 25613 8194
rect 14246 8156 14260 8170
rect 21350 8156 21364 8170
rect 21374 8156 21388 8170
rect 25599 8156 25613 8170
rect 16022 8132 16036 8146
rect 21326 8132 21340 8146
rect 21350 8132 21364 8146
rect 25599 8132 25613 8146
rect 16766 8108 16780 8122
rect 21398 8108 21412 8122
rect 21422 8108 21436 8122
rect 25599 8108 25613 8122
rect 18758 8084 18772 8098
rect 21446 8084 21460 8098
rect 21470 8084 21484 8098
rect 25599 8084 25613 8098
rect 11726 7251 11740 7265
rect 11750 7251 11764 7265
rect 14942 7251 14956 7265
rect 15614 7251 15628 7265
rect 22814 7251 22828 7265
rect 23702 7251 23716 7265
rect 11606 7227 11620 7241
rect 11846 7227 11860 7241
rect 14750 7227 14764 7241
rect 15398 7227 15412 7241
rect 19238 7227 19252 7241
rect 20702 7227 20716 7241
rect 22814 7227 22828 7241
rect 24614 7227 24628 7241
rect 11126 7203 11140 7217
rect 11798 7203 11812 7217
rect 12470 7203 12484 7217
rect 14750 7203 14764 7217
rect 14894 7203 14908 7217
rect 20390 7203 20404 7217
rect 10502 7179 10516 7193
rect 11126 7179 11140 7193
rect 11342 7179 11356 7193
rect 17270 7179 17284 7193
rect 10454 7155 10468 7169
rect 17054 7155 17068 7169
rect 18422 7155 18436 7169
rect 10406 7131 10420 7145
rect 23726 7131 23740 7145
rect 24470 7131 24484 7145
rect 10142 7107 10156 7121
rect 15806 7107 15820 7121
rect 20294 7107 20308 7121
rect 24062 7107 24076 7121
rect 10142 7083 10156 7097
rect 21782 7083 21796 7097
rect 9518 7059 9532 7073
rect 19838 7059 19852 7073
rect 9206 7035 9220 7049
rect 16454 7035 16468 7049
rect 9038 7011 9052 7025
rect 18110 7011 18124 7025
rect 20462 7011 20476 7025
rect 8846 6987 8860 7001
rect 18710 6987 18724 7001
rect 8798 6963 8812 6977
rect 21302 6963 21316 6977
rect 8750 6939 8764 6953
rect 9038 6939 9052 6953
rect 9134 6939 9148 6953
rect 15254 6939 15268 6953
rect 22358 6939 22372 6953
rect 22838 6939 22852 6953
rect 8678 6915 8692 6929
rect 9302 6915 9316 6929
rect 9518 6915 9532 6929
rect 18254 6915 18268 6929
rect 8654 6891 8668 6905
rect 19334 6891 19348 6905
rect 8438 6867 8452 6881
rect 21398 6867 21412 6881
rect 8390 6843 8404 6857
rect 18326 6843 18340 6857
rect 8318 6819 8332 6833
rect 10118 6819 10132 6833
rect 10982 6819 10996 6833
rect 17462 6819 17476 6833
rect 18134 6819 18148 6833
rect 8294 6795 8308 6809
rect 9182 6795 9196 6809
rect 15446 6795 15460 6809
rect 19310 6795 19324 6809
rect 8294 6771 8308 6785
rect 21710 6771 21724 6785
rect 8246 6747 8260 6761
rect 8438 6747 8452 6761
rect 8486 6747 8500 6761
rect 13598 6747 13612 6761
rect 14414 6747 14428 6761
rect 17582 6747 17596 6761
rect 8198 6723 8212 6737
rect 18398 6723 18412 6737
rect 8126 6699 8140 6713
rect 8174 6699 8188 6713
rect 8222 6699 8236 6713
rect 9686 6699 9700 6713
rect 13838 6699 13852 6713
rect 14510 6699 14524 6713
rect 22382 6699 22396 6713
rect 24014 6699 24028 6713
rect 7982 6675 7996 6689
rect 21206 6675 21220 6689
rect 7934 6651 7948 6665
rect 21230 6651 21244 6665
rect 24446 6651 24460 6665
rect 24662 6651 24676 6665
rect 7886 6627 7900 6641
rect 12470 6627 12484 6641
rect 24446 6627 24460 6641
rect 7790 6603 7804 6617
rect 11006 6603 11020 6617
rect 11174 6603 11188 6617
rect 19046 6603 19060 6617
rect 20990 6603 21004 6617
rect 7718 6579 7732 6593
rect 18686 6579 18700 6593
rect 7622 6555 7636 6569
rect 9086 6555 9100 6569
rect 18350 6555 18364 6569
rect 7550 6531 7564 6545
rect 9566 6531 9580 6545
rect 17798 6531 17812 6545
rect 7382 6507 7396 6521
rect 17390 6507 17404 6521
rect 7358 6483 7372 6497
rect 9326 6483 9340 6497
rect 9470 6483 9484 6497
rect 19934 6483 19948 6497
rect 7310 6459 7324 6473
rect 11990 6459 12004 6473
rect 20294 6459 20308 6473
rect 22118 6459 22132 6473
rect 23486 6459 23500 6473
rect 7214 6435 7228 6449
rect 14894 6435 14908 6449
rect 15494 6435 15508 6449
rect 7166 6411 7180 6425
rect 7694 6411 7708 6425
rect 17294 6411 17308 6425
rect 20918 6411 20932 6425
rect 7022 6387 7036 6401
rect 16694 6387 16708 6401
rect 6662 6363 6676 6377
rect 21902 6363 21916 6377
rect 6446 6339 6460 6353
rect 21494 6339 21508 6353
rect 6302 6315 6316 6329
rect 6326 6315 6340 6329
rect 6374 6315 6388 6329
rect 7238 6315 7252 6329
rect 7598 6315 7612 6329
rect 12062 6315 12076 6329
rect 15734 6315 15748 6329
rect 19094 6315 19108 6329
rect 22790 6315 22804 6329
rect 23198 6315 23212 6329
rect 6206 6291 6220 6305
rect 8198 6291 8212 6305
rect 12398 6291 12412 6305
rect 17798 6291 17812 6305
rect 18326 6291 18340 6305
rect 6158 6267 6172 6281
rect 20702 6267 20716 6281
rect 6110 6243 6124 6257
rect 6758 6243 6772 6257
rect 9542 6243 9556 6257
rect 10550 6243 10564 6257
rect 15014 6243 15028 6257
rect 20342 6243 20356 6257
rect 5750 6219 5764 6233
rect 21614 6219 21628 6233
rect 5390 6195 5404 6209
rect 14918 6195 14932 6209
rect 5390 6171 5404 6185
rect 12494 6171 12508 6185
rect 14174 6171 14188 6185
rect 18878 6171 18892 6185
rect 5366 6147 5380 6161
rect 7166 6147 7180 6161
rect 8678 6147 8692 6161
rect 22622 6147 22636 6161
rect 23318 6147 23332 6161
rect 5366 6123 5380 6137
rect 15278 6123 15292 6137
rect 5342 6099 5356 6113
rect 21590 6099 21604 6113
rect 25262 6099 25276 6113
rect 5294 6075 5308 6089
rect 22910 6075 22924 6089
rect 5270 6051 5284 6065
rect 5942 6051 5956 6065
rect 23078 6051 23092 6065
rect 5270 6027 5284 6041
rect 17342 6027 17356 6041
rect 5222 6003 5236 6017
rect 5918 6003 5932 6017
rect 21974 6003 21988 6017
rect 5174 5979 5188 5993
rect 8726 5979 8740 5993
rect 14198 5979 14212 5993
rect 14366 5979 14380 5993
rect 15158 5979 15172 5993
rect 5054 5955 5068 5969
rect 22886 5955 22900 5969
rect 24398 5955 24412 5969
rect 5006 5931 5020 5945
rect 14126 5931 14140 5945
rect 16694 5931 16708 5945
rect 21878 5931 21892 5945
rect 23606 5931 23620 5945
rect 4958 5907 4972 5921
rect 21014 5907 21028 5921
rect 21878 5907 21892 5921
rect 4958 5883 4972 5897
rect 6806 5883 6820 5897
rect 6950 5883 6964 5897
rect 11462 5883 11476 5897
rect 15230 5883 15244 5897
rect 18662 5883 18676 5897
rect 18758 5883 18772 5897
rect 19382 5883 19396 5897
rect 19466 5883 19480 5897
rect 20222 5883 20236 5897
rect 20270 5883 20284 5897
rect 22070 5883 22084 5897
rect 22574 5883 22588 5897
rect 4910 5859 4924 5873
rect 5174 5859 5188 5873
rect 5990 5859 6004 5873
rect 18542 5859 18556 5873
rect 20654 5859 20668 5873
rect 22070 5859 22084 5873
rect 4886 5835 4900 5849
rect 18038 5835 18052 5849
rect 22454 5835 22468 5849
rect 23390 5835 23404 5849
rect 23678 5835 23692 5849
rect 4886 5811 4900 5825
rect 7430 5811 7444 5825
rect 7478 5811 7492 5825
rect 9062 5811 9076 5825
rect 12326 5811 12340 5825
rect 14774 5811 14788 5825
rect 23558 5811 23572 5825
rect 4814 5787 4828 5801
rect 22598 5787 22612 5801
rect 25238 5787 25252 5801
rect 4670 5763 4684 5777
rect 13646 5763 13660 5777
rect 19958 5763 19972 5777
rect 20222 5763 20236 5777
rect 21854 5763 21868 5777
rect 21914 5763 21928 5777
rect 22406 5763 22420 5777
rect 24110 5763 24124 5777
rect 4478 5739 4492 5753
rect 23318 5739 23332 5753
rect 4478 5715 4492 5729
rect 22958 5715 22972 5729
rect 4406 5691 4420 5705
rect 4718 5691 4732 5705
rect 9374 5691 9388 5705
rect 10190 5691 10204 5705
rect 10478 5691 10492 5705
rect 12206 5691 12220 5705
rect 17438 5691 17452 5705
rect 17918 5691 17932 5705
rect 18134 5691 18148 5705
rect 18230 5691 18244 5705
rect 19142 5691 19156 5705
rect 24374 5691 24388 5705
rect 24398 5691 24412 5705
rect 24686 5691 24700 5705
rect 25118 5691 25132 5705
rect 4310 5667 4324 5681
rect 21854 5667 21868 5681
rect 22526 5667 22540 5681
rect 4214 5643 4228 5657
rect 5246 5643 5260 5657
rect 21950 5643 21964 5657
rect 22310 5643 22324 5657
rect 22670 5643 22684 5657
rect 4190 5619 4204 5633
rect 13190 5619 13204 5633
rect 13454 5619 13468 5633
rect 24734 5619 24748 5633
rect 4166 5595 4180 5609
rect 4190 5595 4204 5609
rect 4262 5595 4276 5609
rect 8654 5595 8668 5609
rect 17006 5595 17020 5609
rect 18614 5595 18628 5609
rect 23030 5595 23044 5609
rect 24422 5595 24436 5609
rect 4070 5571 4084 5585
rect 14378 5571 14392 5585
rect 17678 5571 17692 5585
rect 18518 5571 18532 5585
rect 22406 5571 22420 5585
rect 4022 5547 4036 5561
rect 14990 5547 15004 5561
rect 22310 5547 22324 5561
rect 3806 5523 3820 5537
rect 21134 5523 21148 5537
rect 3782 5499 3796 5513
rect 5726 5499 5740 5513
rect 8942 5499 8956 5513
rect 15134 5499 15148 5513
rect 23990 5499 24004 5513
rect 3758 5475 3772 5489
rect 10166 5475 10180 5489
rect 10310 5475 10324 5489
rect 11990 5475 12004 5489
rect 12830 5475 12844 5489
rect 20750 5475 20764 5489
rect 3686 5451 3700 5465
rect 5678 5451 5692 5465
rect 8870 5451 8884 5465
rect 10070 5451 10084 5465
rect 14534 5451 14548 5465
rect 19262 5451 19276 5465
rect 24086 5451 24100 5465
rect 3662 5427 3676 5441
rect 8846 5427 8860 5441
rect 13886 5427 13900 5441
rect 16142 5427 16156 5441
rect 19886 5427 19900 5441
rect 3350 5403 3364 5417
rect 18662 5403 18676 5417
rect 20534 5403 20548 5417
rect 3326 5379 3340 5393
rect 11726 5379 11740 5393
rect 17966 5379 17980 5393
rect 18158 5379 18172 5393
rect 18566 5379 18580 5393
rect 19190 5379 19204 5393
rect 19382 5379 19396 5393
rect 22262 5379 22276 5393
rect 22334 5379 22348 5393
rect 23150 5379 23164 5393
rect 25166 5379 25180 5393
rect 3206 5355 3220 5369
rect 8366 5355 8380 5369
rect 8462 5355 8476 5369
rect 13598 5355 13612 5369
rect 15614 5355 15628 5369
rect 17894 5355 17908 5369
rect 21326 5355 21340 5369
rect 23342 5355 23356 5369
rect 23534 5355 23548 5369
rect 3086 5331 3100 5345
rect 11150 5331 11164 5345
rect 23342 5331 23356 5345
rect 3014 5307 3028 5321
rect 3062 5307 3076 5321
rect 3134 5307 3148 5321
rect 9806 5307 9820 5321
rect 9902 5307 9916 5321
rect 22766 5307 22780 5321
rect 2990 5283 3004 5297
rect 17750 5283 17764 5297
rect 20630 5283 20644 5297
rect 2966 5259 2980 5273
rect 12110 5259 12124 5273
rect 12686 5259 12700 5273
rect 21686 5259 21700 5273
rect 2894 5235 2908 5249
rect 20174 5235 20188 5249
rect 2774 5211 2788 5225
rect 11582 5211 11596 5225
rect 11942 5211 11956 5225
rect 18734 5211 18748 5225
rect 2726 5187 2740 5201
rect 10322 5187 10336 5201
rect 15758 5187 15772 5201
rect 17030 5187 17044 5201
rect 17102 5187 17116 5201
rect 17846 5187 17860 5201
rect 19214 5187 19228 5201
rect 20366 5187 20380 5201
rect 20630 5187 20644 5201
rect 2678 5163 2692 5177
rect 7694 5163 7708 5177
rect 17030 5163 17044 5177
rect 17486 5163 17500 5177
rect 23366 5163 23380 5177
rect 2654 5139 2668 5153
rect 9398 5139 9412 5153
rect 9446 5139 9460 5153
rect 20822 5139 20836 5153
rect 2606 5115 2620 5129
rect 5822 5115 5836 5129
rect 6062 5115 6076 5129
rect 11954 5115 11968 5129
rect 12446 5115 12460 5129
rect 13334 5115 13348 5129
rect 13406 5115 13420 5129
rect 16310 5115 16324 5129
rect 17318 5115 17332 5129
rect 18806 5115 18820 5129
rect 22022 5115 22036 5129
rect 2606 5091 2620 5105
rect 21278 5091 21292 5105
rect 2558 5067 2572 5081
rect 9614 5067 9628 5081
rect 24302 5067 24316 5081
rect 2534 5043 2548 5057
rect 3518 5043 3532 5057
rect 10958 5043 10972 5057
rect 11246 5043 11260 5057
rect 12350 5043 12364 5057
rect 15926 5043 15940 5057
rect 24518 5043 24532 5057
rect 2438 5019 2452 5033
rect 6206 5019 6220 5033
rect 6254 5019 6268 5033
rect 21914 5019 21928 5033
rect 2390 4995 2404 5009
rect 4622 4995 4636 5009
rect 12542 4995 12556 5009
rect 20438 4995 20452 5009
rect 2294 4971 2308 4985
rect 3302 4971 3316 4985
rect 4646 4971 4660 4985
rect 11918 4971 11932 4985
rect 12278 4971 12292 4985
rect 21038 4971 21052 4985
rect 2270 4947 2284 4961
rect 4862 4947 4876 4961
rect 7622 4947 7636 4961
rect 7934 4947 7948 4961
rect 8126 4947 8140 4961
rect 10286 4947 10300 4961
rect 11678 4947 11692 4961
rect 12110 4947 12124 4961
rect 14942 4947 14956 4961
rect 15830 4947 15844 4961
rect 19118 4947 19132 4961
rect 20870 4947 20884 4961
rect 2270 4923 2284 4937
rect 16910 4923 16924 4937
rect 17246 4923 17260 4937
rect 17534 4923 17548 4937
rect 17702 4923 17716 4937
rect 23438 4923 23452 4937
rect 2174 4899 2188 4913
rect 20726 4899 20740 4913
rect 21062 4899 21076 4913
rect 21410 4899 21424 4913
rect 21806 4899 21820 4913
rect 21830 4899 21844 4913
rect 2102 4875 2116 4889
rect 5558 4875 5572 4889
rect 10670 4875 10684 4889
rect 10718 4875 10732 4889
rect 25598 4875 25612 4889
rect 2078 4851 2092 4865
rect 2510 4851 2524 4865
rect 4814 4851 4828 4865
rect 5966 4851 5980 4865
rect 15518 4851 15532 4865
rect 16478 4851 16492 4865
rect 20414 4851 20428 4865
rect 21470 4851 21484 4865
rect 21806 4851 21820 4865
rect 24494 4851 24508 4865
rect 2054 4827 2068 4841
rect 6014 4827 6028 4841
rect 6350 4827 6364 4841
rect 21062 4827 21076 4841
rect 1982 4803 1996 4817
rect 4742 4803 4756 4817
rect 12662 4803 12676 4817
rect 21470 4803 21484 4817
rect 23582 4803 23596 4817
rect 1934 4779 1948 4793
rect 2030 4779 2044 4793
rect 14678 4779 14692 4793
rect 18062 4779 18076 4793
rect 20486 4779 20500 4793
rect 22274 4779 22288 4793
rect 1838 4755 1852 4769
rect 6422 4755 6436 4769
rect 8150 4755 8164 4769
rect 15134 4755 15148 4769
rect 15182 4755 15196 4769
rect 15290 4755 15304 4769
rect 16022 4755 16036 4769
rect 16070 4755 16084 4769
rect 17198 4755 17212 4769
rect 18614 4755 18628 4769
rect 18974 4755 18988 4769
rect 21758 4755 21772 4769
rect 23126 4755 23140 4769
rect 23246 4755 23260 4769
rect 23294 4755 23308 4769
rect 23654 4755 23668 4769
rect 25214 4755 25228 4769
rect 1790 4731 1804 4745
rect 3974 4731 3988 4745
rect 6398 4731 6412 4745
rect 15182 4731 15196 4745
rect 16022 4731 16036 4745
rect 16382 4731 16396 4745
rect 16430 4731 16444 4745
rect 16622 4731 16636 4745
rect 24494 4731 24508 4745
rect 1718 4707 1732 4721
rect 3110 4707 3124 4721
rect 3182 4707 3196 4721
rect 19430 4707 19444 4721
rect 20798 4707 20812 4721
rect 23006 4707 23020 4721
rect 23654 4707 23668 4721
rect 1694 4683 1708 4697
rect 3446 4683 3460 4697
rect 3542 4683 3556 4697
rect 4574 4683 4588 4697
rect 8174 4683 8188 4697
rect 11750 4683 11764 4697
rect 18854 4683 18868 4697
rect 18950 4683 18964 4697
rect 19442 4683 19456 4697
rect 19910 4683 19924 4697
rect 20018 4683 20032 4697
rect 20246 4683 20260 4697
rect 20606 4683 20620 4697
rect 20678 4683 20692 4697
rect 20834 4683 20848 4697
rect 22862 4683 22876 4697
rect 23270 4683 23284 4697
rect 23414 4683 23428 4697
rect 23630 4683 23644 4697
rect 1670 4659 1684 4673
rect 1694 4659 1708 4673
rect 2462 4659 2476 4673
rect 2582 4659 2596 4673
rect 4214 4659 4228 4673
rect 4382 4659 4396 4673
rect 7574 4659 7588 4673
rect 11606 4659 11620 4673
rect 15326 4659 15340 4673
rect 16598 4659 16612 4673
rect 18350 4659 18364 4673
rect 22742 4659 22756 4673
rect 23870 4659 23884 4673
rect 24374 4659 24388 4673
rect 24470 4659 24484 4673
rect 1622 4635 1636 4649
rect 11438 4635 11452 4649
rect 11558 4635 11572 4649
rect 11750 4635 11764 4649
rect 11870 4635 11884 4649
rect 19166 4635 19180 4649
rect 19310 4635 19324 4649
rect 19334 4635 19348 4649
rect 19982 4635 19996 4649
rect 22550 4635 22564 4649
rect 22622 4635 22636 4649
rect 22790 4635 22804 4649
rect 1598 4611 1612 4625
rect 3254 4611 3268 4625
rect 12638 4611 12652 4625
rect 13670 4611 13684 4625
rect 21086 4611 21100 4625
rect 22574 4611 22588 4625
rect 22742 4611 22756 4625
rect 23030 4611 23044 4625
rect 1574 4587 1588 4601
rect 8990 4587 9004 4601
rect 11462 4587 11476 4601
rect 18782 4587 18796 4601
rect 19118 4587 19132 4601
rect 19238 4587 19252 4601
rect 20438 4587 20452 4601
rect 20654 4587 20668 4601
rect 20726 4587 20740 4601
rect 23534 4587 23548 4601
rect 1502 4563 1516 4577
rect 5870 4563 5884 4577
rect 13238 4563 13252 4577
rect 23510 4563 23524 4577
rect 1478 4539 1492 4553
rect 3158 4539 3172 4553
rect 10502 4539 10516 4553
rect 16166 4539 16180 4553
rect 20198 4539 20212 4553
rect 20486 4539 20500 4553
rect 24278 4539 24292 4553
rect 1430 4515 1444 4529
rect 14438 4515 14452 4529
rect 15326 4515 15340 4529
rect 16982 4515 16996 4529
rect 18398 4515 18412 4529
rect 18422 4515 18436 4529
rect 18518 4515 18532 4529
rect 22934 4515 22948 4529
rect 1406 4491 1420 4505
rect 3566 4491 3580 4505
rect 5438 4491 5452 4505
rect 6038 4491 6052 4505
rect 8630 4491 8644 4505
rect 11102 4491 11116 4505
rect 12014 4491 12028 4505
rect 12254 4491 12268 4505
rect 16886 4491 16900 4505
rect 18590 4491 18604 4505
rect 21902 4491 21916 4505
rect 22358 4491 22372 4505
rect 22430 4491 22444 4505
rect 23462 4491 23476 4505
rect 1382 4467 1396 4481
rect 2390 4467 2404 4481
rect 2894 4467 2908 4481
rect 6878 4467 6892 4481
rect 7286 4467 7300 4481
rect 11414 4467 11428 4481
rect 16382 4467 16396 4481
rect 20558 4467 20572 4481
rect 22694 4467 22708 4481
rect 1310 4443 1324 4457
rect 22166 4443 22180 4457
rect 1262 4419 1276 4433
rect 14462 4419 14476 4433
rect 15422 4419 15436 4433
rect 23222 4419 23236 4433
rect 1214 4395 1228 4409
rect 13430 4395 13444 4409
rect 13694 4395 13708 4409
rect 22982 4395 22996 4409
rect 23222 4395 23236 4409
rect 23438 4395 23452 4409
rect 1166 4371 1180 4385
rect 2198 4371 2212 4385
rect 2246 4371 2260 4385
rect 3854 4371 3868 4385
rect 18086 4371 18100 4385
rect 1142 4347 1156 4361
rect 22214 4347 22228 4361
rect 1142 4323 1156 4337
rect 17126 4323 17140 4337
rect 1094 4299 1108 4313
rect 2102 4299 2116 4313
rect 2150 4299 2164 4313
rect 3038 4299 3052 4313
rect 3086 4299 3100 4313
rect 3446 4299 3460 4313
rect 6278 4299 6292 4313
rect 6926 4299 6940 4313
rect 8222 4299 8236 4313
rect 10262 4299 10276 4313
rect 16862 4299 16876 4313
rect 1070 4275 1084 4289
rect 4586 4275 4600 4289
rect 8150 4275 8164 4289
rect 8246 4275 8260 4289
rect 10646 4275 10660 4289
rect 14150 4275 14164 4289
rect 16670 4275 16684 4289
rect 16922 4275 16936 4289
rect 1046 4251 1060 4265
rect 1190 4251 1204 4265
rect 1286 4251 1300 4265
rect 4550 4251 4564 4265
rect 4838 4251 4852 4265
rect 7766 4251 7780 4265
rect 8534 4251 8548 4265
rect 8918 4251 8932 4265
rect 10022 4251 10036 4265
rect 11030 4251 11044 4265
rect 13958 4251 13972 4265
rect 16574 4251 16588 4265
rect 22838 4251 22852 4265
rect 1022 4227 1036 4241
rect 4526 4227 4540 4241
rect 11486 4227 11500 4241
rect 13526 4227 13540 4241
rect 16598 4227 16612 4241
rect 17414 4227 17428 4241
rect 17870 4227 17884 4241
rect 18566 4227 18580 4241
rect 18998 4227 19012 4241
rect 19598 4227 19612 4241
rect 23846 4227 23860 4241
rect 24230 4227 24244 4241
rect 950 4203 964 4217
rect 1166 4203 1180 4217
rect 6686 4203 6700 4217
rect 6854 4203 6868 4217
rect 12566 4203 12580 4217
rect 17894 4203 17908 4217
rect 23918 4203 23932 4217
rect 902 4179 916 4193
rect 1862 4179 1876 4193
rect 1910 4179 1924 4193
rect 9110 4179 9124 4193
rect 9158 4179 9172 4193
rect 14630 4179 14644 4193
rect 21974 4179 21988 4193
rect 22094 4179 22108 4193
rect 830 4155 844 4169
rect 9854 4155 9868 4169
rect 9926 4155 9940 4169
rect 20966 4155 20980 4169
rect 806 4131 820 4145
rect 10910 4131 10924 4145
rect 11174 4131 11188 4145
rect 14822 4131 14836 4145
rect 15446 4131 15460 4145
rect 18062 4131 18076 4145
rect 18494 4131 18508 4145
rect 20966 4131 20980 4145
rect 21086 4131 21100 4145
rect 758 4107 772 4121
rect 8006 4107 8020 4121
rect 8078 4107 8092 4121
rect 11822 4107 11836 4121
rect 11918 4107 11932 4121
rect 11954 4107 11968 4121
rect 12014 4107 12028 4121
rect 23174 4107 23188 4121
rect 734 4083 748 4097
rect 11654 4083 11668 4097
rect 12182 4083 12196 4097
rect 12806 4083 12820 4097
rect 18710 4083 18724 4097
rect 19046 4083 19060 4097
rect 19910 4083 19924 4097
rect 21734 4083 21748 4097
rect 22238 4083 22252 4097
rect 22550 4083 22564 4097
rect 710 4059 724 4073
rect 2486 4059 2500 4073
rect 4286 4059 4300 4073
rect 4934 4059 4948 4073
rect 5198 4059 5212 4073
rect 5486 4059 5500 4073
rect 6158 4059 6172 4073
rect 17822 4059 17836 4073
rect 20318 4059 20332 4073
rect 22046 4059 22060 4073
rect 23054 4059 23068 4073
rect 638 4035 652 4049
rect 2222 4035 2236 4049
rect 6494 4035 6508 4049
rect 6566 4035 6580 4049
rect 16982 4035 16996 4049
rect 23054 4035 23068 4049
rect 23198 4035 23212 4049
rect 590 4011 604 4025
rect 11630 4011 11644 4025
rect 21254 4011 21268 4025
rect 542 3987 556 4001
rect 18470 3987 18484 4001
rect 21254 3987 21268 4001
rect 21326 3987 21340 4001
rect 518 3963 532 3977
rect 8966 3963 8980 3977
rect 9734 3963 9748 3977
rect 10094 3963 10108 3977
rect 11486 3963 11500 3977
rect 20150 3963 20164 3977
rect 494 3939 508 3953
rect 4622 3939 4636 3953
rect 6974 3939 6988 3953
rect 9254 3939 9268 3953
rect 14582 3939 14596 3953
rect 15902 3939 15916 3953
rect 21998 3939 22012 3953
rect 446 3915 460 3929
rect 2846 3915 2860 3929
rect 2918 3915 2932 3929
rect 9758 3915 9772 3929
rect 9950 3915 9964 3929
rect 16622 3915 16636 3929
rect 16862 3915 16876 3929
rect 17006 3915 17020 3929
rect 18470 3915 18484 3929
rect 20018 3915 20032 3929
rect 20150 3915 20164 3929
rect 20174 3915 20188 3929
rect 398 3891 412 3905
rect 5126 3891 5140 3905
rect 7430 3891 7444 3905
rect 8750 3891 8764 3905
rect 8798 3891 8812 3905
rect 16358 3891 16372 3905
rect 374 3867 388 3881
rect 1358 3867 1372 3881
rect 5654 3867 5668 3881
rect 7118 3867 7132 3881
rect 7790 3867 7804 3881
rect 8726 3867 8740 3881
rect 11054 3867 11068 3881
rect 17942 3867 17956 3881
rect 21566 3867 21580 3881
rect 350 3843 364 3857
rect 878 3843 892 3857
rect 926 3843 940 3857
rect 2366 3843 2380 3857
rect 6110 3843 6124 3857
rect 8054 3843 8068 3857
rect 16838 3843 16852 3857
rect 19142 3843 19156 3857
rect 21542 3843 21556 3857
rect 302 3819 316 3833
rect 12590 3819 12604 3833
rect 13742 3819 13756 3833
rect 16502 3819 16516 3833
rect 21542 3819 21556 3833
rect 21590 3819 21604 3833
rect 278 3795 292 3809
rect 974 3795 988 3809
rect 7358 3795 7372 3809
rect 9590 3795 9604 3809
rect 9638 3795 9652 3809
rect 9854 3795 9868 3809
rect 12230 3795 12244 3809
rect 12278 3795 12292 3809
rect 14078 3795 14092 3809
rect 14318 3795 14332 3809
rect 22910 3795 22924 3809
rect 230 3771 244 3785
rect 23414 3771 23428 3785
rect 230 3747 244 3761
rect 6134 3747 6148 3761
rect 6182 3747 6196 3761
rect 16430 3747 16444 3761
rect 182 3723 196 3737
rect 19550 3723 19564 3737
rect 158 3699 172 3713
rect 22646 3699 22660 3713
rect 134 3675 148 3689
rect 10598 3675 10612 3689
rect 10814 3675 10828 3689
rect 24518 3675 24532 3689
rect -1430 3651 -1416 3665
rect 662 3651 676 3665
rect 710 3651 724 3665
rect 6230 3651 6244 3665
rect 10214 3651 10228 3665
rect 11078 3651 11092 3665
rect 11390 3651 11404 3665
rect 18590 3651 18604 3665
rect -1430 3627 -1416 3641
rect 14030 3627 14044 3641
rect 16310 3627 16324 3641
rect 16718 3627 16732 3641
rect -1430 3603 -1416 3617
rect 11294 3603 11308 3617
rect 11702 3603 11716 3617
rect 17102 3603 17116 3617
rect 21446 3603 21460 3617
rect -1430 3579 -1416 3593
rect 7550 3579 7564 3593
rect 7670 3579 7684 3593
rect 7838 3579 7852 3593
rect 9350 3579 9364 3593
rect 9398 3579 9412 3593
rect 9566 3579 9580 3593
rect 9662 3579 9676 3593
rect 10238 3579 10252 3593
rect 10286 3579 10300 3593
rect 10322 3579 10336 3593
rect 10406 3579 10420 3593
rect 11510 3579 11524 3593
rect 11942 3579 11956 3593
rect 24662 3579 24676 3593
rect 110 3555 124 3569
rect 20246 3555 20260 3569
rect 110 3531 124 3545
rect 3014 3531 3028 3545
rect 11774 3531 11788 3545
rect 12182 3531 12196 3545
rect 16526 3531 16540 3545
rect 16958 3531 16972 3545
rect 22214 3531 22228 3545
rect 134 3507 148 3521
rect 3470 3507 3484 3521
rect 5294 3507 5308 3521
rect 7982 3507 7996 3521
rect 9302 3507 9316 3521
rect 12086 3507 12100 3521
rect 13550 3507 13564 3521
rect 14006 3507 14020 3521
rect 16286 3507 16300 3521
rect 17774 3507 17788 3521
rect 20798 3507 20812 3521
rect 20894 3507 20908 3521
rect 21374 3507 21388 3521
rect 158 3483 172 3497
rect 5558 3483 5572 3497
rect 9278 3483 9292 3497
rect 20606 3483 20620 3497
rect 23102 3483 23116 3497
rect 182 3459 196 3473
rect 22190 3459 22204 3473
rect 326 3435 340 3449
rect 1046 3435 1060 3449
rect 1094 3435 1108 3449
rect 18446 3435 18460 3449
rect 20894 3435 20908 3449
rect 20990 3435 21004 3449
rect 22190 3435 22204 3449
rect 22274 3435 22288 3449
rect 614 3411 628 3425
rect 19502 3411 19516 3425
rect 758 3387 772 3401
rect 974 3387 988 3401
rect 4454 3387 4468 3401
rect 4742 3387 4756 3401
rect 7910 3387 7924 3401
rect 9830 3387 9844 3401
rect 11894 3387 11908 3401
rect 12302 3387 12316 3401
rect 14342 3387 14356 3401
rect 14798 3387 14812 3401
rect 16550 3387 16564 3401
rect 18902 3387 18916 3401
rect 18974 3387 18988 3401
rect 854 3363 868 3377
rect 22862 3363 22876 3377
rect 950 3339 964 3353
rect 2006 3339 2020 3353
rect 18014 3339 18028 3353
rect 23774 3339 23788 3353
rect 1070 3315 1084 3329
rect 10886 3315 10900 3329
rect 11366 3315 11380 3329
rect 15350 3315 15364 3329
rect 17222 3315 17236 3329
rect 21134 3315 21148 3329
rect 23582 3315 23596 3329
rect 25070 3315 25084 3329
rect 1526 3291 1540 3305
rect 20678 3291 20692 3305
rect 1742 3267 1756 3281
rect 2630 3267 2644 3281
rect 3062 3267 3076 3281
rect 9422 3267 9436 3281
rect 10382 3267 10396 3281
rect 19574 3267 19588 3281
rect 1766 3243 1780 3257
rect 22766 3243 22780 3257
rect 1814 3219 1828 3233
rect 22478 3219 22492 3233
rect 1886 3195 1900 3209
rect 16046 3195 16060 3209
rect 17990 3195 18004 3209
rect 21158 3195 21172 3209
rect 1934 3171 1948 3185
rect 3638 3171 3652 3185
rect 5150 3171 5164 3185
rect 6086 3171 6100 3185
rect 9878 3171 9892 3185
rect 16814 3171 16828 3185
rect 17222 3171 17236 3185
rect 17270 3171 17284 3185
rect 17774 3171 17788 3185
rect 17966 3171 17980 3185
rect 18110 3171 18124 3185
rect 18446 3171 18460 3185
rect 18542 3171 18556 3185
rect 2030 3147 2044 3161
rect 2534 3147 2548 3161
rect 11558 3147 11572 3161
rect 22934 3147 22948 3161
rect 24206 3147 24220 3161
rect 2054 3123 2068 3137
rect 14222 3123 14236 3137
rect 15206 3123 15220 3137
rect 16742 3123 16756 3137
rect 20006 3123 20020 3137
rect 2318 3099 2332 3113
rect 2774 3099 2788 3113
rect 2870 3099 2884 3113
rect 22262 3099 22276 3113
rect 2342 3075 2356 3089
rect 2438 3075 2452 3089
rect 2558 3075 2572 3089
rect 5774 3075 5788 3089
rect 8606 3075 8620 3089
rect 10358 3075 10372 3089
rect 10766 3075 10780 3089
rect 10862 3075 10876 3089
rect 18878 3075 18892 3089
rect 20834 3075 20848 3089
rect 22718 3075 22732 3089
rect 2366 3051 2380 3065
rect 2390 3051 2404 3065
rect 2486 3051 2500 3065
rect 17630 3051 17644 3065
rect 22718 3051 22732 3065
rect 22886 3051 22900 3065
rect 2390 3027 2404 3041
rect 8414 3027 8428 3041
rect 8606 3027 8620 3041
rect 8654 3027 8668 3041
rect 8702 3027 8716 3041
rect 15038 3027 15052 3041
rect 16718 3027 16732 3041
rect 20510 3027 20524 3041
rect 2678 3003 2692 3017
rect 4766 3003 4780 3017
rect 7382 3003 7396 3017
rect 7502 3003 7516 3017
rect 17078 3003 17092 3017
rect 17654 3003 17668 3017
rect 24566 3003 24580 3017
rect 2942 2979 2956 2993
rect 16238 2979 16252 2993
rect 16814 2979 16828 2993
rect 16922 2979 16936 2993
rect 17630 2979 17644 2993
rect 17678 2979 17692 2993
rect 2990 2955 3004 2969
rect 5846 2955 5860 2969
rect 7334 2955 7348 2969
rect 19070 2955 19084 2969
rect 23462 2955 23476 2969
rect 3110 2931 3124 2945
rect 21182 2931 21196 2945
rect 3206 2907 3220 2921
rect 3494 2907 3508 2921
rect 15110 2907 15124 2921
rect 16454 2907 16468 2921
rect 19070 2907 19084 2921
rect 22142 2907 22156 2921
rect 3254 2883 3268 2897
rect 7886 2883 7900 2897
rect 8102 2883 8116 2897
rect 9710 2883 9724 2897
rect 18830 2883 18844 2897
rect 19790 2883 19804 2897
rect 21662 2883 21676 2897
rect 23966 2883 23980 2897
rect 3326 2859 3340 2873
rect 11750 2859 11764 2873
rect 15290 2859 15304 2873
rect 20774 2859 20788 2873
rect 23126 2859 23140 2873
rect 3590 2835 3604 2849
rect 9758 2835 9772 2849
rect 9974 2835 9988 2849
rect 11006 2835 11020 2849
rect 19622 2835 19636 2849
rect 21182 2835 21196 2849
rect 21206 2835 21220 2849
rect 3710 2811 3724 2825
rect 11246 2811 11260 2825
rect 11294 2811 11308 2825
rect 11846 2811 11860 2825
rect 12206 2811 12220 2825
rect 24326 2811 24340 2825
rect 3902 2787 3916 2801
rect 4166 2787 4180 2801
rect 4238 2787 4252 2801
rect 6398 2787 6412 2801
rect 7094 2787 7108 2801
rect 8558 2787 8572 2801
rect 20582 2787 20596 2801
rect 24182 2787 24196 2801
rect 24710 2787 24724 2801
rect 3974 2763 3988 2777
rect 5894 2763 5908 2777
rect 5966 2763 5980 2777
rect 6206 2763 6220 2777
rect 6254 2763 6268 2777
rect 6710 2763 6724 2777
rect 15398 2763 15412 2777
rect 3998 2739 4012 2753
rect 22958 2739 22972 2753
rect 4022 2715 4036 2729
rect 4190 2715 4204 2729
rect 12590 2715 12604 2729
rect 16190 2715 16204 2729
rect 4094 2691 4108 2705
rect 14702 2691 14716 2705
rect 4118 2667 4132 2681
rect 5414 2667 5428 2681
rect 5582 2667 5596 2681
rect 6302 2667 6316 2681
rect 10694 2667 10708 2681
rect 12518 2667 12532 2681
rect 13766 2667 13780 2681
rect 24542 2667 24556 2681
rect 4334 2643 4348 2657
rect 13382 2643 13396 2657
rect 15638 2643 15652 2657
rect 16358 2643 16372 2657
rect 18758 2643 18772 2657
rect 4550 2619 4564 2633
rect 4586 2619 4600 2633
rect 4670 2619 4684 2633
rect 9494 2619 9508 2633
rect 9734 2619 9748 2633
rect 10022 2619 10036 2633
rect 10094 2619 10108 2633
rect 10118 2619 10132 2633
rect 10310 2619 10324 2633
rect 23246 2619 23260 2633
rect 4934 2595 4948 2609
rect 16214 2595 16228 2609
rect 5054 2571 5068 2585
rect 10646 2571 10660 2585
rect 19022 2571 19036 2585
rect 5126 2547 5140 2561
rect 5174 2547 5188 2561
rect 5222 2547 5236 2561
rect 15278 2547 15292 2561
rect 23630 2547 23644 2561
rect 5702 2523 5716 2537
rect 12398 2523 12412 2537
rect 13382 2523 13396 2537
rect 22502 2523 22516 2537
rect 5774 2499 5788 2513
rect 15470 2499 15484 2513
rect 15542 2499 15556 2513
rect 19358 2499 19372 2513
rect 5894 2475 5908 2489
rect 5942 2475 5956 2489
rect 6014 2475 6028 2489
rect 11582 2475 11596 2489
rect 24590 2475 24604 2489
rect 6134 2451 6148 2465
rect 6278 2451 6292 2465
rect 6374 2451 6388 2465
rect 7718 2451 7732 2465
rect 10790 2451 10804 2465
rect 11414 2451 11428 2465
rect 24158 2451 24172 2465
rect 6230 2427 6244 2441
rect 6422 2427 6436 2441
rect 6470 2427 6484 2441
rect 15062 2427 15076 2441
rect 19022 2427 19036 2441
rect 19094 2427 19108 2441
rect 6518 2403 6532 2417
rect 9950 2403 9964 2417
rect 9998 2403 10012 2417
rect 23822 2403 23836 2417
rect 6590 2379 6604 2393
rect 15854 2379 15868 2393
rect 6614 2355 6628 2369
rect 13574 2355 13588 2369
rect 13958 2355 13972 2369
rect 24638 2355 24652 2369
rect 6782 2331 6796 2345
rect 7094 2331 7108 2345
rect 7142 2331 7156 2345
rect 12734 2331 12748 2345
rect 25190 2331 25204 2345
rect 7238 2307 7252 2321
rect 10238 2307 10252 2321
rect 16262 2307 16276 2321
rect 18038 2307 18052 2321
rect 7262 2283 7276 2297
rect 12374 2283 12388 2297
rect 14342 2283 14356 2297
rect 14378 2283 14392 2297
rect 16262 2283 16276 2297
rect 16406 2283 16420 2297
rect 7838 2259 7852 2273
rect 11822 2259 11836 2273
rect 18926 2259 18940 2273
rect 19466 2259 19480 2273
rect 20102 2259 20116 2273
rect 7910 2235 7924 2249
rect 7934 2235 7948 2249
rect 8030 2235 8044 2249
rect 14294 2235 14308 2249
rect 16406 2235 16420 2249
rect 21350 2235 21364 2249
rect 8774 2211 8788 2225
rect 9998 2211 10012 2225
rect 17558 2211 17572 2225
rect 19166 2211 19180 2225
rect 20270 2211 20284 2225
rect 20942 2211 20956 2225
rect 22670 2211 22684 2225
rect 9230 2187 9244 2201
rect 10598 2187 10612 2201
rect 11198 2187 11212 2201
rect 20918 2187 20932 2201
rect 25142 2187 25156 2201
rect 9254 2163 9268 2177
rect 9326 2163 9340 2177
rect 9494 2163 9508 2177
rect 9686 2163 9700 2177
rect 9782 2163 9796 2177
rect 21110 2163 21124 2177
rect 21350 2163 21364 2177
rect 21410 2163 21424 2177
rect 25262 2163 25276 2177
rect 25599 2163 25613 2177
rect 9326 2139 9340 2153
rect 21830 2139 21844 2153
rect 25238 2139 25252 2153
rect 25599 2139 25613 2153
rect 10046 2115 10060 2129
rect 19406 2115 19420 2129
rect 21614 2115 21628 2129
rect 25214 2115 25228 2129
rect 25599 2115 25613 2129
rect 10526 2091 10540 2105
rect 16070 2091 16084 2105
rect 21398 2091 21412 2105
rect 25190 2091 25204 2105
rect 25599 2091 25613 2105
rect 10550 2067 10564 2081
rect 14870 2067 14884 2081
rect 19406 2067 19420 2081
rect 19442 2067 19456 2081
rect 25166 2067 25180 2081
rect 25599 2067 25613 2081
rect 10574 2043 10588 2057
rect 10838 2043 10852 2057
rect 11078 2043 11092 2057
rect 11150 2043 11164 2057
rect 25142 2043 25156 2057
rect 25599 2043 25613 2057
rect 10358 1210 10372 1224
rect 16166 1210 16180 1224
rect 16766 1210 16780 1224
rect 19454 1210 19468 1224
rect 9902 1186 9916 1200
rect 19694 1186 19708 1200
rect 9566 1162 9580 1176
rect 20078 1162 20092 1176
rect 8918 1138 8932 1152
rect 16262 1138 16276 1152
rect 16742 1138 16756 1152
rect 19190 1138 19204 1152
rect 8870 1114 8884 1128
rect 10022 1114 10036 1128
rect 10118 1114 10132 1128
rect 12830 1114 12844 1128
rect 16478 1114 16492 1128
rect 16958 1114 16972 1128
rect 22574 1114 22588 1128
rect 24734 1114 24748 1128
rect 8630 1090 8644 1104
rect 9206 1090 9220 1104
rect 18494 1090 18508 1104
rect 20462 1090 20476 1104
rect 24806 1090 24820 1104
rect 8558 1066 8572 1080
rect 8942 1066 8956 1080
rect 9038 1066 9052 1080
rect 20690 1066 20704 1080
rect 8510 1042 8524 1056
rect 8894 1042 8908 1056
rect 8990 1042 9004 1056
rect 11270 1042 11284 1056
rect 12422 1042 12436 1056
rect 19814 1042 19828 1056
rect 8486 1018 8500 1032
rect 23174 1018 23188 1032
rect 8342 994 8356 1008
rect 11750 994 11764 1008
rect 12326 994 12340 1008
rect 18206 994 18220 1008
rect 8318 970 8332 984
rect 17846 970 17860 984
rect 7934 946 7948 960
rect 8534 946 8548 960
rect 21014 946 21028 960
rect 6422 922 6436 936
rect 21278 922 21292 936
rect 6278 898 6292 912
rect 19742 898 19756 912
rect 5966 874 5980 888
rect 11318 874 11332 888
rect 12230 874 12244 888
rect 19262 874 19276 888
rect 5486 850 5500 864
rect 7814 850 7828 864
rect 10094 850 10108 864
rect 11678 850 11692 864
rect 20558 850 20572 864
rect 21758 850 21772 864
rect 21998 850 22012 864
rect 23006 850 23020 864
rect 24782 850 24796 864
rect 5438 826 5452 840
rect 6542 826 6556 840
rect 7742 826 7756 840
rect 11150 826 11164 840
rect 11198 826 11212 840
rect 23618 826 23632 840
rect 5318 802 5332 816
rect 21230 802 21244 816
rect 5174 778 5188 792
rect 23510 778 23524 792
rect 4982 754 4996 768
rect 7190 754 7204 768
rect 7478 754 7492 768
rect 13982 754 13996 768
rect 17102 754 17116 768
rect 4646 730 4660 744
rect 5510 730 5524 744
rect 5606 730 5620 744
rect 14102 730 14116 744
rect 14198 730 14212 744
rect 24758 730 24772 744
rect 4574 706 4588 720
rect 23390 706 23404 720
rect 4490 682 4504 696
rect 15470 682 15484 696
rect 15662 682 15676 696
rect 18110 682 18124 696
rect 18158 682 18172 696
rect 24542 682 24556 696
rect 4430 658 4444 672
rect 20366 658 20380 672
rect 4406 634 4420 648
rect 15974 634 15988 648
rect 16190 634 16204 648
rect 19238 634 19252 648
rect 19670 634 19684 648
rect 22358 634 22372 648
rect 23222 634 23236 648
rect 24590 634 24604 648
rect 24710 634 24724 648
rect 3614 610 3628 624
rect 5006 610 5020 624
rect 5078 610 5092 624
rect 20894 610 20908 624
rect 24710 610 24724 624
rect 3398 586 3412 600
rect 20102 586 20116 600
rect 3350 562 3364 576
rect 22646 562 22660 576
rect 3134 538 3148 552
rect 7646 538 7660 552
rect 8006 538 8020 552
rect 8102 538 8116 552
rect 20582 538 20596 552
rect 3062 514 3076 528
rect 20846 514 20860 528
rect 3014 490 3028 504
rect 15230 490 15244 504
rect 15710 490 15724 504
rect 21662 490 21676 504
rect 2918 466 2932 480
rect 16574 466 16588 480
rect 17738 466 17752 480
rect 21350 466 21364 480
rect 2870 442 2884 456
rect 18830 442 18844 456
rect 2846 418 2860 432
rect 12134 418 12148 432
rect 12974 418 12988 432
rect 20030 418 20044 432
rect 2798 394 2812 408
rect 20822 394 20836 408
rect 2750 370 2764 384
rect 10886 370 10900 384
rect 15566 370 15580 384
rect 16274 370 16288 384
rect 23270 370 23284 384
rect 2702 346 2716 360
rect 14174 346 14188 360
rect 14810 346 14824 360
rect 21926 346 21940 360
rect 2174 322 2188 336
rect 9350 322 9364 336
rect 9446 322 9460 336
rect 10430 322 10444 336
rect 10718 322 10732 336
rect 16094 322 16108 336
rect 2150 298 2164 312
rect 14222 298 14236 312
rect 2126 274 2140 288
rect 11510 274 11524 288
rect 13790 274 13804 288
rect 18806 274 18820 288
rect 1334 250 1348 264
rect 10454 250 10468 264
rect 10742 250 10756 264
rect 18278 250 18292 264
rect 1214 226 1228 240
rect 8366 226 8380 240
rect 8438 226 8452 240
rect 10430 226 10444 240
rect 10790 226 10804 240
rect 11966 226 11980 240
rect 14006 226 14020 240
rect 18926 226 18940 240
rect -1430 202 -1416 216
rect 20630 202 20644 216
rect -1430 178 -1416 192
rect 230 178 244 192
rect 902 178 916 192
rect 998 178 1012 192
rect 16670 178 16684 192
rect -1430 154 -1416 168
rect 7094 154 7108 168
rect 7442 154 7456 168
rect 22430 154 22444 168
rect -1430 130 -1416 144
rect 10838 130 10852 144
rect 10934 130 10948 144
rect 16934 130 16948 144
rect 24710 130 24724 144
rect 25599 130 25613 144
rect 2294 106 2308 120
rect 17762 106 17776 120
rect 24806 106 24820 120
rect 25599 106 25613 120
rect 4166 82 4180 96
rect 19226 82 19240 96
rect 24782 82 24796 96
rect 25599 82 25613 96
rect 5726 58 5740 72
rect 24710 58 24724 72
rect 24758 58 24772 72
rect 25599 58 25613 72
rect 9086 34 9100 48
rect 11906 34 11920 48
rect 24734 34 24748 48
rect 25599 34 25613 48
rect 9950 10 9964 24
rect 10334 10 10348 24
rect 12854 10 12868 24
rect 24710 10 24724 24
rect 25599 10 25613 24
<< metal2 >>
rect -1500 8253 -1430 8265
rect -1500 8229 -1430 8241
rect -1500 8205 -1430 8217
rect -1377 8074 -1177 8276
rect -1161 8074 -1149 8276
rect -1137 8074 -1125 8276
rect -1113 8074 -1101 8276
rect -1089 8074 -1077 8276
rect 231 8074 243 8228
rect 423 8074 435 8204
rect 3399 8074 3411 8204
rect 5607 8074 5619 8228
rect 6303 8074 6315 8204
rect 13479 8074 13491 8180
rect 14247 8074 14259 8156
rect 16023 8074 16035 8132
rect 16767 8074 16779 8108
rect 18759 8074 18771 8084
rect 21303 8074 21315 8252
rect 21327 8146 21339 8252
rect 21375 8170 21387 8204
rect 21351 8146 21363 8156
rect 21399 8122 21411 8204
rect 21423 8122 21435 8180
rect 21447 8098 21459 8180
rect 21471 8098 21483 8228
rect 25359 8074 25559 8276
rect 25613 8253 25683 8265
rect 25613 8205 25683 8217
rect 25613 8181 25683 8193
rect 25613 8157 25683 8169
rect 25613 8133 25683 8145
rect 25613 8109 25683 8121
rect 25613 8085 25683 8097
rect -1500 3652 -1430 3664
rect -1500 3628 -1430 3640
rect -1500 3604 -1430 3616
rect -1500 3580 -1430 3592
rect -1377 2033 -1177 7275
rect -1161 2033 -1149 7275
rect -1137 2033 -1125 7275
rect -1113 2033 -1101 7275
rect -1089 2033 -1077 7275
rect 111 3569 123 7275
rect 135 3689 147 7275
rect 159 3713 171 7275
rect 183 3737 195 7275
rect 231 3785 243 7275
rect 279 3809 291 7275
rect 303 3833 315 7275
rect 111 2033 123 3531
rect 135 2033 147 3507
rect 159 2033 171 3483
rect 183 2033 195 3459
rect 231 2033 243 3747
rect 327 3449 339 7275
rect 375 3881 387 7275
rect 399 3905 411 7275
rect 447 3929 459 7275
rect 495 3953 507 7275
rect 519 3977 531 7275
rect 543 4001 555 7275
rect 591 4025 603 7275
rect 351 2033 363 3843
rect 615 3425 627 7275
rect 639 4049 651 7275
rect 663 3665 675 7275
rect 711 4073 723 7275
rect 735 4097 747 7275
rect 759 4121 771 7275
rect 807 4145 819 7275
rect 831 4169 843 7275
rect 711 2033 723 3651
rect 759 2033 771 3387
rect 855 3377 867 7275
rect 879 3857 891 7275
rect 903 2033 915 4179
rect 927 3857 939 7275
rect 951 4217 963 7275
rect 975 3809 987 7275
rect 1023 4241 1035 7275
rect 1047 4265 1059 7275
rect 1071 4289 1083 7275
rect 1095 4313 1107 7275
rect 1143 4361 1155 7275
rect 1167 4385 1179 7275
rect 1215 4409 1227 7275
rect 1263 4433 1275 7275
rect 951 2033 963 3339
rect 975 2033 987 3387
rect 1047 2033 1059 3435
rect 1071 2033 1083 3315
rect 1095 2033 1107 3435
rect 1143 2033 1155 4323
rect 1287 4265 1299 7275
rect 1311 4457 1323 7275
rect 1167 2033 1179 4203
rect 1191 2033 1203 4251
rect 1359 3881 1371 7275
rect 1383 4481 1395 7275
rect 1407 4505 1419 7275
rect 1431 4529 1443 7275
rect 1479 4553 1491 7275
rect 1503 4577 1515 7275
rect 1527 3305 1539 7275
rect 1575 4601 1587 7275
rect 1599 4625 1611 7275
rect 1623 4649 1635 7275
rect 1671 4673 1683 7275
rect 1695 4697 1707 7275
rect 1719 4721 1731 7275
rect 1695 2033 1707 4659
rect 1743 2033 1755 3267
rect 1767 3257 1779 7275
rect 1791 4745 1803 7275
rect 1815 3233 1827 7275
rect 1839 4769 1851 7275
rect 1863 4193 1875 7275
rect 1911 4193 1923 7275
rect 1935 4793 1947 7275
rect 1983 4817 1995 7275
rect 2031 4793 2043 7275
rect 2055 4841 2067 7275
rect 2079 4865 2091 7275
rect 2103 4889 2115 7275
rect 2151 4313 2163 7275
rect 2175 4913 2187 7275
rect 1887 2033 1899 3195
rect 1935 2033 1947 3171
rect 2007 2033 2019 3339
rect 2031 2033 2043 3147
rect 2055 2033 2067 3123
rect 2103 2033 2115 4299
rect 2199 2033 2211 4371
rect 2223 4049 2235 7275
rect 2271 4961 2283 7275
rect 2295 4985 2307 7275
rect 2247 2033 2259 4371
rect 2271 2033 2283 4923
rect 2319 3113 2331 7275
rect 2367 3857 2379 7275
rect 2391 5009 2403 7275
rect 2439 5033 2451 7275
rect 2343 2033 2355 3075
rect 2391 3065 2403 4467
rect 2367 2033 2379 3051
rect 2391 2033 2403 3027
rect 2439 2033 2451 3075
rect 2463 2033 2475 4659
rect 2487 4073 2499 7275
rect 2511 4865 2523 7275
rect 2535 5057 2547 7275
rect 2559 5081 2571 7275
rect 2607 5129 2619 7275
rect 2487 2033 2499 3051
rect 2535 2033 2547 3147
rect 2559 2033 2571 3075
rect 2583 2033 2595 4659
rect 2607 2033 2619 5091
rect 2631 3281 2643 7275
rect 2679 5177 2691 7275
rect 2727 5201 2739 7275
rect 2775 5225 2787 7275
rect 2655 2033 2667 5139
rect 2847 3929 2859 7275
rect 2871 3113 2883 7275
rect 2895 5249 2907 7275
rect 2679 2033 2691 3003
rect 2775 2033 2787 3099
rect 2895 2033 2907 4467
rect 2919 3929 2931 7275
rect 2943 2993 2955 7275
rect 2991 5297 3003 7275
rect 3015 5321 3027 7275
rect 2967 2033 2979 5259
rect 3039 4313 3051 7275
rect 3087 5345 3099 7275
rect 2991 2033 3003 2955
rect 3015 2033 3027 3531
rect 3063 3281 3075 5307
rect 3111 4721 3123 7275
rect 3135 5321 3147 7275
rect 3183 4721 3195 7275
rect 3207 5369 3219 7275
rect 3255 4625 3267 7275
rect 3303 4985 3315 7275
rect 3327 5393 3339 7275
rect 3351 5417 3363 7275
rect 3447 4697 3459 7275
rect 3519 5057 3531 7275
rect 3543 4697 3555 7275
rect 3087 2033 3099 4299
rect 3111 2033 3123 2931
rect 3159 2033 3171 4539
rect 3567 4505 3579 7275
rect 3207 2033 3219 2907
rect 3255 2033 3267 2883
rect 3327 2033 3339 2859
rect 3447 2033 3459 4299
rect 3471 2033 3483 3507
rect 3495 2033 3507 2907
rect 3591 2849 3603 7275
rect 3639 3185 3651 7275
rect 3663 5441 3675 7275
rect 3687 5465 3699 7275
rect 3711 2825 3723 7275
rect 3759 5489 3771 7275
rect 3783 5513 3795 7275
rect 3807 5537 3819 7275
rect 3855 4385 3867 7275
rect 3903 2801 3915 7275
rect 3975 4745 3987 7275
rect 3975 2033 3987 2763
rect 3999 2753 4011 7275
rect 4023 5561 4035 7275
rect 4071 5585 4083 7275
rect 4023 2033 4035 2715
rect 4095 2705 4107 7275
rect 4119 2681 4131 7275
rect 4167 5609 4179 7275
rect 4191 5633 4203 7275
rect 4215 5657 4227 7275
rect 4263 5609 4275 7275
rect 4167 2033 4179 2787
rect 4191 2729 4203 5595
rect 4215 2033 4227 4659
rect 4287 4073 4299 7275
rect 4311 5681 4323 7275
rect 4383 4673 4395 7275
rect 4407 5705 4419 7275
rect 4455 3401 4467 7275
rect 4479 5753 4491 7275
rect 4239 2033 4251 2787
rect 4335 2033 4347 2643
rect 4479 2033 4491 5715
rect 4551 4265 4563 7275
rect 4575 4697 4587 7275
rect 4623 5009 4635 7275
rect 4671 5777 4683 7275
rect 4527 2033 4539 4227
rect 4587 2633 4599 4275
rect 4551 2033 4563 2619
rect 4623 2033 4635 3939
rect 4647 2033 4659 4971
rect 4671 2033 4683 2619
rect 4719 2033 4731 5691
rect 4743 4817 4755 7275
rect 4815 5801 4827 7275
rect 4887 5849 4899 7275
rect 4911 5873 4923 7275
rect 4743 2033 4755 3387
rect 4767 2033 4779 3003
rect 4815 2033 4827 4851
rect 4839 2033 4851 4251
rect 4863 2033 4875 4947
rect 4887 2033 4899 5811
rect 4935 4073 4947 7275
rect 4959 5921 4971 7275
rect 5007 5945 5019 7275
rect 5055 5969 5067 7275
rect 4935 2033 4947 2595
rect 4959 2033 4971 5883
rect 5127 3905 5139 7275
rect 5151 3185 5163 7275
rect 5175 5993 5187 7275
rect 5223 6017 5235 7275
rect 5055 2033 5067 2571
rect 5175 2561 5187 5859
rect 5247 5657 5259 7275
rect 5271 6065 5283 7275
rect 5295 6089 5307 7275
rect 5343 6113 5355 7275
rect 5367 6161 5379 7275
rect 5391 6209 5403 7275
rect 5127 2033 5139 2547
rect 5199 2033 5211 4059
rect 5223 2033 5235 2547
rect 5271 2033 5283 6027
rect 5295 2033 5307 3507
rect 5367 2033 5379 6123
rect 5391 2033 5403 6171
rect 5439 4505 5451 7275
rect 5487 4073 5499 7275
rect 5559 4889 5571 7275
rect 5415 2033 5427 2667
rect 5559 2033 5571 3483
rect 5583 2681 5595 7275
rect 5655 3881 5667 7275
rect 5679 5465 5691 7275
rect 5655 2033 5667 3867
rect 5703 2537 5715 7275
rect 5751 6233 5763 7275
rect 5727 2033 5739 5499
rect 5775 3089 5787 7275
rect 5823 5129 5835 7275
rect 5871 4577 5883 7275
rect 5775 2033 5787 2499
rect 5847 2033 5859 2955
rect 5895 2777 5907 7275
rect 5919 6017 5931 7275
rect 5943 2489 5955 6051
rect 5967 4865 5979 7275
rect 5991 5873 6003 7275
rect 6015 4841 6027 7275
rect 6039 4505 6051 7275
rect 6063 5129 6075 7275
rect 6111 6257 6123 7275
rect 5895 2033 5907 2475
rect 5967 2033 5979 2763
rect 6015 2033 6027 2475
rect 6087 2033 6099 3171
rect 6111 2033 6123 3843
rect 6135 3761 6147 7275
rect 6159 6281 6171 7275
rect 6207 6305 6219 7275
rect 6135 2033 6147 2451
rect 6159 2033 6171 4059
rect 6183 2033 6195 3747
rect 6207 2777 6219 5019
rect 6231 3665 6243 7275
rect 6255 5033 6267 7275
rect 6303 6329 6315 7275
rect 6231 2033 6243 2427
rect 6255 2033 6267 2763
rect 6279 2465 6291 4299
rect 6303 2033 6315 2667
rect 6327 2033 6339 6315
rect 6351 4841 6363 7275
rect 6375 6329 6387 7275
rect 6399 4745 6411 7275
rect 6447 6353 6459 7275
rect 6375 2033 6387 2451
rect 6399 2033 6411 2787
rect 6423 2441 6435 4755
rect 6471 2441 6483 7275
rect 6495 4049 6507 7275
rect 6519 2417 6531 7275
rect 6567 4049 6579 7275
rect 6591 2393 6603 7275
rect 6615 2369 6627 7275
rect 6663 6377 6675 7275
rect 6687 4217 6699 7275
rect 6711 2777 6723 7275
rect 6759 6257 6771 7275
rect 6783 2345 6795 7275
rect 6807 5897 6819 7275
rect 6855 4217 6867 7275
rect 6879 4481 6891 7275
rect 6927 4313 6939 7275
rect 6951 2033 6963 5883
rect 6975 3953 6987 7275
rect 7023 6401 7035 7275
rect 7095 2801 7107 7275
rect 7119 3881 7131 7275
rect 7167 6425 7179 7275
rect 7215 6449 7227 7275
rect 7239 6329 7251 7275
rect 7095 2033 7107 2331
rect 7143 2033 7155 2331
rect 7167 2033 7179 6147
rect 7239 2033 7251 2307
rect 7263 2297 7275 7275
rect 7311 6473 7323 7275
rect 7287 2033 7299 4467
rect 7335 2969 7347 7275
rect 7359 6497 7371 7275
rect 7383 6521 7395 7275
rect 7431 5825 7443 7275
rect 7479 5825 7491 7275
rect 7551 6545 7563 7275
rect 7575 4673 7587 7275
rect 7623 6569 7635 7275
rect 7359 2033 7371 3795
rect 7383 2033 7395 3003
rect 7431 2033 7443 3891
rect 7503 2033 7515 3003
rect 7551 2033 7563 3579
rect 7599 2033 7611 6315
rect 7623 2033 7635 4947
rect 7671 3593 7683 7275
rect 7695 6425 7707 7275
rect 7719 6593 7731 7275
rect 7695 2033 7707 5163
rect 7767 4265 7779 7275
rect 7791 6617 7803 7275
rect 7719 2033 7731 2451
rect 7791 2033 7803 3867
rect 7839 3593 7851 7275
rect 7887 6641 7899 7275
rect 7911 3401 7923 7275
rect 7935 6665 7947 7275
rect 7983 6689 7995 7275
rect 7839 2033 7851 2259
rect 7887 2033 7899 2883
rect 7935 2249 7947 4947
rect 8007 4121 8019 7275
rect 7911 2033 7923 2235
rect 7983 2033 7995 3507
rect 8031 2249 8043 7275
rect 8079 4121 8091 7275
rect 8055 2033 8067 3843
rect 8103 2897 8115 7275
rect 8127 6713 8139 7275
rect 8127 2033 8139 4947
rect 8151 4769 8163 7275
rect 8199 6737 8211 7275
rect 8223 6713 8235 7275
rect 8247 6761 8259 7275
rect 8295 6809 8307 7275
rect 8319 6833 8331 7275
rect 8175 4697 8187 6699
rect 8151 2033 8163 4275
rect 8199 2033 8211 6291
rect 8223 2033 8235 4299
rect 8247 2033 8259 4275
rect 8295 2033 8307 6771
rect 8367 5369 8379 7275
rect 8391 2033 8403 6843
rect 8415 3041 8427 7275
rect 8439 6881 8451 7275
rect 8439 2033 8451 6747
rect 8463 5369 8475 7275
rect 8487 6761 8499 7275
rect 8535 4265 8547 7275
rect 8559 2801 8571 7275
rect 8607 3089 8619 7275
rect 8655 6905 8667 7275
rect 8679 6929 8691 7275
rect 8607 2033 8619 3027
rect 8631 2033 8643 4491
rect 8655 3041 8667 5595
rect 8679 2033 8691 6147
rect 8703 3041 8715 7275
rect 8727 5993 8739 7275
rect 8751 6953 8763 7275
rect 8799 6977 8811 7275
rect 8847 7001 8859 7275
rect 8727 2033 8739 3867
rect 8751 2033 8763 3891
rect 8775 2033 8787 2211
rect 8799 2033 8811 3891
rect 8847 2033 8859 5427
rect 8871 2033 8883 5451
rect 8919 4265 8931 7275
rect 8943 5513 8955 7275
rect 8991 4601 9003 7275
rect 9039 7025 9051 7275
rect 8967 2033 8979 3963
rect 9039 2033 9051 6939
rect 9063 5825 9075 7275
rect 9087 2033 9099 6555
rect 9111 4193 9123 7275
rect 9135 2033 9147 6939
rect 9159 4193 9171 7275
rect 9183 6809 9195 7275
rect 9207 7049 9219 7275
rect 9255 3953 9267 7275
rect 9279 3497 9291 7275
rect 9303 6929 9315 7275
rect 9231 2033 9243 2187
rect 9255 2033 9267 2163
rect 9303 2033 9315 3507
rect 9327 2177 9339 6483
rect 9351 3593 9363 7275
rect 9375 5705 9387 7275
rect 9399 5153 9411 7275
rect 9447 5153 9459 7275
rect 9471 6497 9483 7275
rect 9327 2033 9339 2139
rect 9399 2033 9411 3579
rect 9423 2033 9435 3267
rect 9495 2633 9507 7275
rect 9519 7073 9531 7275
rect 9495 2033 9507 2163
rect 9519 2033 9531 6915
rect 9543 6257 9555 7275
rect 9567 3593 9579 6531
rect 9591 3809 9603 7275
rect 9615 2033 9627 5067
rect 9639 3809 9651 7275
rect 9663 2033 9675 3579
rect 9687 2177 9699 6699
rect 9711 2897 9723 7275
rect 9735 3977 9747 7275
rect 9759 3929 9771 7275
rect 9807 5321 9819 7275
rect 9831 3401 9843 7275
rect 9855 4169 9867 7275
rect 9903 5321 9915 7275
rect 9927 4169 9939 7275
rect 9951 3929 9963 7275
rect 9735 2033 9747 2619
rect 9759 2033 9771 2835
rect 9783 2033 9795 2163
rect 9831 2033 9843 3387
rect 9855 2033 9867 3795
rect 9879 2033 9891 3171
rect 9975 2849 9987 7275
rect 9999 2417 10011 7275
rect 10071 5465 10083 7275
rect 10023 2633 10035 4251
rect 10095 3977 10107 7275
rect 10143 7121 10155 7275
rect 10119 2633 10131 6819
rect 9951 2033 9963 2403
rect 9999 2033 10011 2211
rect 10047 2033 10059 2115
rect 10095 2033 10107 2619
rect 10143 2033 10155 7083
rect 10167 5489 10179 7275
rect 10191 2033 10203 5691
rect 10215 2033 10227 3651
rect 10239 3593 10251 7275
rect 10263 4313 10275 7275
rect 10287 4961 10299 7275
rect 10311 5489 10323 7275
rect 10323 3593 10335 5187
rect 10239 2033 10251 2307
rect 10287 2033 10299 3579
rect 10359 3089 10371 7275
rect 10383 3281 10395 7275
rect 10407 7145 10419 7275
rect 10455 7169 10467 7275
rect 10479 5705 10491 7275
rect 10503 7193 10515 7275
rect 10551 6257 10563 7275
rect 10311 2033 10323 2619
rect 10407 2033 10419 3579
rect 10503 2033 10515 4539
rect 10527 2033 10539 2091
rect 10551 2033 10563 2067
rect 10575 2057 10587 7275
rect 10599 3689 10611 7275
rect 10647 4289 10659 7275
rect 10671 4889 10683 7275
rect 10695 2681 10707 7275
rect 10719 4889 10731 7275
rect 10767 3089 10779 7275
rect 10599 2033 10611 2187
rect 10647 2033 10659 2571
rect 10791 2465 10803 7275
rect 10815 3689 10827 7275
rect 10863 3089 10875 7275
rect 10887 3329 10899 7275
rect 10911 4145 10923 7275
rect 10959 5057 10971 7275
rect 10983 6833 10995 7275
rect 11007 6617 11019 7275
rect 10839 2033 10851 2043
rect 11007 2033 11019 2835
rect 11031 2033 11043 4251
rect 11055 3881 11067 7275
rect 11079 3665 11091 7275
rect 11103 4505 11115 7275
rect 11127 7217 11139 7275
rect 11079 2033 11091 2043
rect 11127 2033 11139 7179
rect 11175 6617 11187 7275
rect 11151 2057 11163 5331
rect 11175 2033 11187 4131
rect 11199 2201 11211 7275
rect 11247 5057 11259 7275
rect 11295 3617 11307 7275
rect 11343 7193 11355 7275
rect 11415 4481 11427 7275
rect 11439 4649 11451 7275
rect 11463 5897 11475 7275
rect 11247 2033 11259 2811
rect 11295 2033 11307 2811
rect 11367 2033 11379 3315
rect 11391 2033 11403 3651
rect 11415 2033 11427 2451
rect 11463 2033 11475 4587
rect 11487 4241 11499 7275
rect 11487 2033 11499 3963
rect 11511 3593 11523 7275
rect 11559 4649 11571 7275
rect 11583 5225 11595 7275
rect 11607 7241 11619 7275
rect 11559 2033 11571 3147
rect 11583 2033 11595 2475
rect 11607 2033 11619 4659
rect 11655 4097 11667 7275
rect 11679 4961 11691 7275
rect 11727 7265 11739 7275
rect 11631 2033 11643 4011
rect 11703 2033 11715 3603
rect 11727 2033 11739 5379
rect 11751 4697 11763 7251
rect 11751 2873 11763 4635
rect 11775 3545 11787 7275
rect 11799 2033 11811 7203
rect 11823 4121 11835 7275
rect 11847 2825 11859 7227
rect 11823 2033 11835 2259
rect 11871 2033 11883 4635
rect 11895 3401 11907 7275
rect 11919 4985 11931 7275
rect 11943 5225 11955 7275
rect 11991 6473 12003 7275
rect 11955 4121 11967 5115
rect 11919 2033 11931 4107
rect 11943 2033 11955 3579
rect 11991 2033 12003 5475
rect 12015 4505 12027 7275
rect 12015 2033 12027 4107
rect 12063 2033 12075 6315
rect 12111 5273 12123 7275
rect 12087 2033 12099 3507
rect 12111 2033 12123 4947
rect 12183 4097 12195 7275
rect 12207 5705 12219 7275
rect 12231 3809 12243 7275
rect 12255 4505 12267 7275
rect 12279 4985 12291 7275
rect 12327 5825 12339 7275
rect 12351 5057 12363 7275
rect 12399 6305 12411 7275
rect 12447 5129 12459 7275
rect 12471 7217 12483 7275
rect 12183 2033 12195 3531
rect 12207 2033 12219 2811
rect 12279 2033 12291 3795
rect 12303 2033 12315 3387
rect 12375 2033 12387 2283
rect 12399 2033 12411 2523
rect 12471 2033 12483 6627
rect 12495 6185 12507 7275
rect 12543 5009 12555 7275
rect 12567 4217 12579 7275
rect 12591 3833 12603 7275
rect 12639 4625 12651 7275
rect 12687 5273 12699 7275
rect 12831 5489 12843 7275
rect 13191 5633 13203 7275
rect 12519 2033 12531 2667
rect 12591 2033 12603 2715
rect 12663 2033 12675 4803
rect 13239 4577 13251 7275
rect 12735 2033 12747 2331
rect 12807 2033 12819 4083
rect 13335 2033 13347 5115
rect 13383 2657 13395 7275
rect 13407 5129 13419 7275
rect 13431 4409 13443 7275
rect 13455 5633 13467 7275
rect 13599 6761 13611 7275
rect 13383 2033 13395 2523
rect 13527 2033 13539 4227
rect 13551 2033 13563 3507
rect 13575 2033 13587 2355
rect 13599 2033 13611 5355
rect 13647 2033 13659 5763
rect 13671 2033 13683 4611
rect 13695 2033 13707 4395
rect 13743 2033 13755 3819
rect 13767 2033 13779 2667
rect 13839 2033 13851 6699
rect 13887 2033 13899 5427
rect 13959 4265 13971 7275
rect 14007 3521 14019 7275
rect 13959 2033 13971 2355
rect 14031 2033 14043 3627
rect 14079 2033 14091 3795
rect 14127 2033 14139 5931
rect 14151 4289 14163 7275
rect 14175 6185 14187 7275
rect 14199 5993 14211 7275
rect 14223 3137 14235 7275
rect 14295 2249 14307 7275
rect 14319 3809 14331 7275
rect 14343 3401 14355 7275
rect 14367 5993 14379 7275
rect 14415 6761 14427 7275
rect 14379 2297 14391 5571
rect 14439 4529 14451 7275
rect 14463 4433 14475 7275
rect 14511 6713 14523 7275
rect 14535 5465 14547 7275
rect 14583 3953 14595 7275
rect 14631 4193 14643 7275
rect 14679 4793 14691 7275
rect 14751 7241 14763 7275
rect 14343 2033 14355 2283
rect 14703 2033 14715 2691
rect 14751 2033 14763 7203
rect 14775 5825 14787 7275
rect 14799 3401 14811 7275
rect 14823 4145 14835 7275
rect 14871 2081 14883 7275
rect 14895 7217 14907 7275
rect 14895 2033 14907 6435
rect 14919 6209 14931 7275
rect 14943 7265 14955 7275
rect 14991 5561 15003 7275
rect 14943 2033 14955 4947
rect 15015 2033 15027 6243
rect 15039 3041 15051 7275
rect 15111 2921 15123 7275
rect 15135 5513 15147 7275
rect 15063 2033 15075 2427
rect 15135 2033 15147 4755
rect 15159 2033 15171 5979
rect 15183 4769 15195 7275
rect 15231 5897 15243 7275
rect 15255 6953 15267 7275
rect 15279 6137 15291 7275
rect 15183 2033 15195 4731
rect 15207 2033 15219 3123
rect 15291 2873 15303 4755
rect 15327 4673 15339 7275
rect 15279 2033 15291 2547
rect 15327 2033 15339 4515
rect 15351 3329 15363 7275
rect 15399 7241 15411 7275
rect 15447 6809 15459 7275
rect 15399 2033 15411 2763
rect 15423 2033 15435 4419
rect 15447 2033 15459 4131
rect 15471 2513 15483 7275
rect 15495 6449 15507 7275
rect 15615 7265 15627 7275
rect 15519 2033 15531 4851
rect 15543 2033 15555 2499
rect 15615 2033 15627 5355
rect 15639 2033 15651 2643
rect 15735 2033 15747 6315
rect 15759 2033 15771 5187
rect 15807 2033 15819 7107
rect 15831 2033 15843 4947
rect 15855 2033 15867 2379
rect 15903 2033 15915 3939
rect 15927 2033 15939 5043
rect 16023 4769 16035 7275
rect 16023 2033 16035 4731
rect 16047 2033 16059 3195
rect 16071 2105 16083 4755
rect 16143 2033 16155 5427
rect 16167 4553 16179 7275
rect 16191 2729 16203 7275
rect 16215 2609 16227 7275
rect 16239 2033 16251 2979
rect 16263 2321 16275 7275
rect 16287 3521 16299 7275
rect 16311 5129 16323 7275
rect 16359 3905 16371 7275
rect 16383 4745 16395 7275
rect 16263 2033 16275 2283
rect 16311 2033 16323 3627
rect 16359 2033 16371 2643
rect 16383 2033 16395 4467
rect 16407 2297 16419 7275
rect 16455 7049 16467 7275
rect 16479 4865 16491 7275
rect 16431 3761 16443 4731
rect 16503 3833 16515 7275
rect 16407 2033 16419 2235
rect 16455 2033 16467 2907
rect 16527 2033 16539 3531
rect 16551 3401 16563 7275
rect 16575 4265 16587 7275
rect 16599 4673 16611 7275
rect 16623 4745 16635 7275
rect 16671 4289 16683 7275
rect 16695 6401 16707 7275
rect 16599 2033 16611 4227
rect 16623 2033 16635 3915
rect 16695 2033 16707 5931
rect 16719 3641 16731 7275
rect 16743 3137 16755 7275
rect 16815 3185 16827 7275
rect 16839 3857 16851 7275
rect 16863 4313 16875 7275
rect 16887 4505 16899 7275
rect 16911 4937 16923 7275
rect 16719 2033 16731 3027
rect 16815 2033 16827 2979
rect 16863 2033 16875 3915
rect 16923 2993 16935 4275
rect 16959 3545 16971 7275
rect 16983 4529 16995 7275
rect 16983 2033 16995 4035
rect 17007 3929 17019 5595
rect 17031 5201 17043 7275
rect 17031 2033 17043 5163
rect 17055 2033 17067 7155
rect 17079 3017 17091 7275
rect 17103 3617 17115 5187
rect 17127 4337 17139 7275
rect 17199 4769 17211 7275
rect 17223 3329 17235 7275
rect 17247 4937 17259 7275
rect 17271 3185 17283 7179
rect 17295 6425 17307 7275
rect 17319 5129 17331 7275
rect 17343 6041 17355 7275
rect 17391 6521 17403 7275
rect 17415 4241 17427 7275
rect 17439 5705 17451 7275
rect 17463 6833 17475 7275
rect 17487 5177 17499 7275
rect 17535 4937 17547 7275
rect 17223 2033 17235 3171
rect 17559 2225 17571 7275
rect 17583 6761 17595 7275
rect 17631 3065 17643 7275
rect 17655 3017 17667 7275
rect 17679 2993 17691 5571
rect 17703 4937 17715 7275
rect 17751 5297 17763 7275
rect 17775 3521 17787 7275
rect 17799 6545 17811 7275
rect 17631 2033 17643 2979
rect 17775 2033 17787 3171
rect 17799 2033 17811 6291
rect 17847 5201 17859 7275
rect 17871 4241 17883 7275
rect 17895 5369 17907 7275
rect 17823 2033 17835 4059
rect 17895 2033 17907 4203
rect 17919 2033 17931 5691
rect 17943 3881 17955 7275
rect 17967 5393 17979 7275
rect 17991 3209 18003 7275
rect 18039 5849 18051 7275
rect 18063 4793 18075 7275
rect 18087 4385 18099 7275
rect 17967 2033 17979 3171
rect 18015 2033 18027 3339
rect 18039 2033 18051 2307
rect 18063 2033 18075 4131
rect 18111 3185 18123 7011
rect 18135 6833 18147 7275
rect 18135 2033 18147 5691
rect 18159 5393 18171 7275
rect 18255 6929 18267 7275
rect 18327 6857 18339 7275
rect 18351 6569 18363 7275
rect 18399 6737 18411 7275
rect 18231 2033 18243 5691
rect 18327 2033 18339 6291
rect 18351 2033 18363 4659
rect 18423 4529 18435 7155
rect 18399 2033 18411 4515
rect 18447 3449 18459 7275
rect 18471 4001 18483 7275
rect 18495 4145 18507 7275
rect 18519 5585 18531 7275
rect 18447 2033 18459 3171
rect 18471 2033 18483 3915
rect 18519 2033 18531 4515
rect 18543 3185 18555 5859
rect 18567 5393 18579 7275
rect 18591 4505 18603 7275
rect 18615 5609 18627 7275
rect 18663 5897 18675 7275
rect 18687 6593 18699 7275
rect 18711 7001 18723 7275
rect 18567 2033 18579 4227
rect 18591 2033 18603 3651
rect 18615 2033 18627 4755
rect 18663 2033 18675 5403
rect 18735 5225 18747 7275
rect 18711 2033 18723 4083
rect 18759 2657 18771 5883
rect 18807 5129 18819 7275
rect 18783 2033 18795 4587
rect 18831 2897 18843 7275
rect 18855 4697 18867 7275
rect 18879 6185 18891 7275
rect 18879 2033 18891 3075
rect 18903 2033 18915 3387
rect 18927 2273 18939 7275
rect 18951 4697 18963 7275
rect 18975 4769 18987 7275
rect 18975 2033 18987 3387
rect 18999 2033 19011 4227
rect 19023 2585 19035 7275
rect 19047 6617 19059 7275
rect 19023 2033 19035 2427
rect 19047 2033 19059 4083
rect 19071 2969 19083 7275
rect 19071 2033 19083 2907
rect 19095 2441 19107 6315
rect 19119 4961 19131 7275
rect 19143 5705 19155 7275
rect 19167 4649 19179 7275
rect 19191 5393 19203 7275
rect 19215 5201 19227 7275
rect 19239 4601 19251 7227
rect 19263 5465 19275 7275
rect 19311 6809 19323 7275
rect 19335 4649 19347 6891
rect 19383 5897 19395 7275
rect 19119 2033 19131 4587
rect 19143 2033 19155 3843
rect 19167 2033 19179 2211
rect 19311 2033 19323 4635
rect 19359 2033 19371 2499
rect 19383 2033 19395 5379
rect 19407 2129 19419 7275
rect 19431 4721 19443 7275
rect 19443 2081 19455 4683
rect 19467 2273 19479 5883
rect 19551 3737 19563 7275
rect 19407 2033 19419 2067
rect 19503 2033 19515 3411
rect 19575 2033 19587 3267
rect 19599 2033 19611 4227
rect 19623 2033 19635 2835
rect 19791 2033 19803 2883
rect 19839 2033 19851 7059
rect 19887 2033 19899 5427
rect 19911 4697 19923 7275
rect 19911 2033 19923 4083
rect 19935 2033 19947 6483
rect 19959 5777 19971 7275
rect 19983 2033 19995 4635
rect 20019 3929 20031 4683
rect 20007 2033 20019 3123
rect 20103 2273 20115 7275
rect 20151 3977 20163 7275
rect 20223 5897 20235 7275
rect 20175 3929 20187 5235
rect 20151 2033 20163 3915
rect 20199 2033 20211 4539
rect 20223 2033 20235 5763
rect 20247 4697 20259 7275
rect 20295 7121 20307 7275
rect 20247 2033 20259 3555
rect 20271 2225 20283 5883
rect 20295 2033 20307 6459
rect 20343 6257 20355 7275
rect 20367 5201 20379 7275
rect 20391 7217 20403 7275
rect 20439 5009 20451 7275
rect 20463 7025 20475 7275
rect 20319 2033 20331 4059
rect 20415 2033 20427 4851
rect 20487 4793 20499 7275
rect 20439 2033 20451 4587
rect 20487 2033 20499 4539
rect 20511 3041 20523 7275
rect 20535 2033 20547 5403
rect 20559 4481 20571 7275
rect 20583 2801 20595 7275
rect 20631 5297 20643 7275
rect 20607 3497 20619 4683
rect 20631 2033 20643 5187
rect 20655 4601 20667 5859
rect 20679 4697 20691 7275
rect 20703 7241 20715 7275
rect 20679 2033 20691 3291
rect 20703 2033 20715 6267
rect 20727 4913 20739 7275
rect 20727 2033 20739 4587
rect 20751 2033 20763 5475
rect 20775 2873 20787 7275
rect 20799 4721 20811 7275
rect 20823 5153 20835 7275
rect 20871 4961 20883 7275
rect 20799 2033 20811 3507
rect 20835 3089 20847 4683
rect 20895 3521 20907 7275
rect 20919 6425 20931 7275
rect 20895 2033 20907 3435
rect 20943 2225 20955 7275
rect 20967 4169 20979 7275
rect 20919 2033 20931 2187
rect 20967 2033 20979 4131
rect 20991 3449 21003 6603
rect 21015 5921 21027 7275
rect 21039 4985 21051 7275
rect 21063 4913 21075 7275
rect 21063 2033 21075 4827
rect 21087 4145 21099 4611
rect 21111 2177 21123 7275
rect 21135 5537 21147 7275
rect 21135 2033 21147 3315
rect 21159 2033 21171 3195
rect 21183 2945 21195 7275
rect 21207 2849 21219 6675
rect 21231 6665 21243 7275
rect 21255 4025 21267 7275
rect 21279 5105 21291 7275
rect 21183 2033 21195 2835
rect 21255 2033 21267 3987
rect 21303 2033 21315 6963
rect 21327 4001 21339 5355
rect 21351 2249 21363 7275
rect 21375 3521 21387 7275
rect 21399 6881 21411 7275
rect 21411 2177 21423 4899
rect 21447 3617 21459 7275
rect 21471 4865 21483 7275
rect 21495 6353 21507 7275
rect 21351 2033 21363 2163
rect 21399 2033 21411 2091
rect 21471 2033 21483 4803
rect 21543 3857 21555 7275
rect 21567 3881 21579 7275
rect 21615 6233 21627 7275
rect 21591 3833 21603 6099
rect 21543 2033 21555 3819
rect 21663 2897 21675 7275
rect 21687 5273 21699 7275
rect 21711 6785 21723 7275
rect 21759 4769 21771 7275
rect 21783 7097 21795 7275
rect 21807 4913 21819 7275
rect 21855 5777 21867 7275
rect 21879 5945 21891 7275
rect 21903 6377 21915 7275
rect 21615 2033 21627 2115
rect 21735 2033 21747 4083
rect 21807 2033 21819 4851
rect 21831 2153 21843 4899
rect 21855 2033 21867 5667
rect 21879 2033 21891 5907
rect 21915 5033 21927 5763
rect 21951 5657 21963 7275
rect 21975 6017 21987 7275
rect 21903 2033 21915 4491
rect 21975 2033 21987 4179
rect 21999 3953 22011 7275
rect 22023 2033 22035 5115
rect 22047 4073 22059 7275
rect 22071 5897 22083 7275
rect 22071 2033 22083 5859
rect 22095 4193 22107 7275
rect 22119 2033 22131 6459
rect 22143 2921 22155 7275
rect 22167 4457 22179 7275
rect 22191 3473 22203 7275
rect 22215 4361 22227 7275
rect 22263 5393 22275 7275
rect 22311 5657 22323 7275
rect 22191 2033 22203 3435
rect 22215 2033 22227 3531
rect 22239 2033 22251 4083
rect 22275 3449 22287 4779
rect 22263 2033 22275 3099
rect 22311 2033 22323 5547
rect 22335 2033 22347 5379
rect 22359 4505 22371 6939
rect 22383 6713 22395 7275
rect 22407 5777 22419 7275
rect 22455 5849 22467 7275
rect 22407 2033 22419 5571
rect 22431 2033 22443 4491
rect 22479 2033 22491 3219
rect 22503 2537 22515 7275
rect 22527 5681 22539 7275
rect 22551 4649 22563 7275
rect 22575 4625 22587 5883
rect 22599 5801 22611 7275
rect 22623 6161 22635 7275
rect 22551 2033 22563 4083
rect 22623 2033 22635 4635
rect 22647 3713 22659 7275
rect 22671 2225 22683 5643
rect 22695 4481 22707 7275
rect 22719 3089 22731 7275
rect 22743 4673 22755 7275
rect 22767 5321 22779 7275
rect 22815 7265 22827 7275
rect 22791 4649 22803 6315
rect 22719 2033 22731 3051
rect 22743 2033 22755 4611
rect 22767 2033 22779 3243
rect 22815 2033 22827 7227
rect 22839 6953 22851 7275
rect 22863 4697 22875 7275
rect 22911 6089 22923 7275
rect 22839 2033 22851 4251
rect 22863 2033 22875 3363
rect 22887 3065 22899 5955
rect 22935 4529 22947 7275
rect 22959 5729 22971 7275
rect 22983 4409 22995 7275
rect 23007 4721 23019 7275
rect 23031 4625 23043 5595
rect 23055 4073 23067 7275
rect 23079 6065 23091 7275
rect 22911 2033 22923 3795
rect 22935 2033 22947 3147
rect 22959 2033 22971 2739
rect 23055 2033 23067 4035
rect 23103 3497 23115 7275
rect 23127 4769 23139 7275
rect 23127 2033 23139 2859
rect 23151 2033 23163 5379
rect 23175 4121 23187 7275
rect 23199 4049 23211 6315
rect 23223 4433 23235 7275
rect 23295 4769 23307 7275
rect 23319 6161 23331 7275
rect 23223 2033 23235 4395
rect 23247 2633 23259 4755
rect 23271 2033 23283 4683
rect 23319 2033 23331 5739
rect 23343 5369 23355 7275
rect 23391 5849 23403 7275
rect 23343 2033 23355 5331
rect 23367 2033 23379 5163
rect 23415 4697 23427 7275
rect 23439 4409 23451 4923
rect 23463 4505 23475 7275
rect 23415 2033 23427 3771
rect 23463 2033 23475 2955
rect 23487 2033 23499 6459
rect 23511 4577 23523 7275
rect 23535 4601 23547 5355
rect 23559 2033 23571 5811
rect 23583 4817 23595 7275
rect 23583 2033 23595 3315
rect 23607 2033 23619 5931
rect 23655 4769 23667 7275
rect 23631 2561 23643 4683
rect 23655 2033 23667 4707
rect 23679 2033 23691 5835
rect 23703 2033 23715 7251
rect 23727 7145 23739 7275
rect 23775 3353 23787 7275
rect 23847 4241 23859 7275
rect 23871 4673 23883 7275
rect 23919 4217 23931 7275
rect 23967 2897 23979 7275
rect 23991 5513 24003 7275
rect 24015 6713 24027 7275
rect 24063 7121 24075 7275
rect 24087 5465 24099 7275
rect 24111 5777 24123 7275
rect 24159 2465 24171 7275
rect 24207 3161 24219 7275
rect 24279 4553 24291 7275
rect 24303 5081 24315 7275
rect 23823 2033 23835 2403
rect 24183 2033 24195 2787
rect 24231 2033 24243 4227
rect 24327 2825 24339 7275
rect 24375 5705 24387 7275
rect 24399 5969 24411 7275
rect 24375 2033 24387 4659
rect 24399 2033 24411 5691
rect 24423 5609 24435 7275
rect 24447 6665 24459 7275
rect 24447 2033 24459 6627
rect 24471 4673 24483 7131
rect 24495 4865 24507 7275
rect 24519 5057 24531 7275
rect 24495 2033 24507 4731
rect 24519 2033 24531 3675
rect 24543 2681 24555 7275
rect 24567 2033 24579 3003
rect 24591 2489 24603 7275
rect 24615 7241 24627 7275
rect 24639 2369 24651 7275
rect 24663 3593 24675 6651
rect 24687 5705 24699 7275
rect 24711 2801 24723 7275
rect 24735 5633 24747 7275
rect 25071 2033 25083 3315
rect 25119 2033 25131 5691
rect 25143 2057 25155 2187
rect 25167 2081 25179 5379
rect 25191 2105 25203 2331
rect 25215 2129 25227 4755
rect 25239 2153 25251 5787
rect 25263 2177 25275 6099
rect 25359 2033 25559 7275
rect 25612 4876 25683 4888
rect 25613 2164 25683 2176
rect 25613 2140 25683 2152
rect 25613 2116 25683 2128
rect 25613 2092 25683 2104
rect 25613 2068 25683 2080
rect 25613 2044 25683 2056
rect -1500 203 -1430 215
rect -1500 179 -1430 191
rect -1500 155 -1430 167
rect -1500 131 -1430 143
rect -1377 0 -1177 1234
rect -1161 0 -1149 1234
rect -1137 0 -1125 1234
rect -1113 0 -1101 1234
rect -1089 0 -1077 1234
rect 231 192 243 1234
rect 903 192 915 1234
rect 999 192 1011 1234
rect 1215 240 1227 1234
rect 1335 264 1347 1234
rect 2127 288 2139 1234
rect 2151 312 2163 1234
rect 2175 336 2187 1234
rect 916 178 934 192
rect 915 0 927 178
rect 2295 120 2307 1234
rect 2703 360 2715 1234
rect 2751 384 2763 1234
rect 2799 408 2811 1234
rect 2847 432 2859 1234
rect 2871 456 2883 1234
rect 2919 480 2931 1234
rect 3063 528 3075 1234
rect 3135 552 3147 1234
rect 3351 576 3363 1234
rect 3399 600 3411 1234
rect 3615 624 3627 1234
rect 3015 0 3027 490
rect 4167 96 4179 1234
rect 4407 648 4419 1234
rect 4431 672 4443 1234
rect 4575 720 4587 1234
rect 4647 744 4659 1234
rect 4983 768 4995 1234
rect 4491 0 4503 682
rect 5007 624 5019 1234
rect 5079 624 5091 1234
rect 5175 792 5187 1234
rect 5319 816 5331 1234
rect 5439 840 5451 1234
rect 5487 864 5499 1234
rect 5511 744 5523 1234
rect 5607 744 5619 1234
rect 5727 72 5739 1234
rect 6279 912 6291 1234
rect 6423 936 6435 1234
rect 5967 0 5979 874
rect 6543 840 6555 1234
rect 7095 168 7107 1234
rect 7191 768 7203 1234
rect 7479 768 7491 1234
rect 7647 552 7659 1234
rect 7743 840 7755 1234
rect 7815 864 7827 1234
rect 7935 960 7947 1234
rect 8007 552 8019 1234
rect 8103 552 8115 1234
rect 8319 984 8331 1234
rect 8343 1008 8355 1234
rect 8367 240 8379 1234
rect 8439 240 8451 1234
rect 8487 1032 8499 1234
rect 8511 1056 8523 1234
rect 8535 960 8547 1234
rect 8559 1080 8571 1234
rect 8631 1104 8643 1234
rect 8871 1128 8883 1234
rect 8895 1056 8907 1234
rect 7443 0 7455 154
rect 8919 0 8931 1138
rect 8943 1080 8955 1234
rect 8991 1056 9003 1234
rect 9039 1080 9051 1234
rect 9087 48 9099 1234
rect 9207 1104 9219 1234
rect 9351 336 9363 1234
rect 9447 336 9459 1234
rect 9567 1176 9579 1234
rect 9903 1200 9915 1234
rect 9951 24 9963 1234
rect 10023 1128 10035 1234
rect 10095 864 10107 1234
rect 10119 1128 10131 1234
rect 10335 24 10347 1234
rect 10359 1224 10371 1234
rect 10431 336 10443 1234
rect 10455 264 10467 1234
rect 10719 336 10731 1234
rect 10743 264 10755 1234
rect 10791 240 10803 1234
rect 9964 10 9982 24
rect 9963 0 9975 10
rect 10431 0 10443 226
rect 10839 144 10851 1234
rect 10887 384 10899 1234
rect 10935 144 10947 1234
rect 11151 840 11163 1234
rect 11199 840 11211 1234
rect 11271 1056 11283 1234
rect 11319 888 11331 1234
rect 11511 288 11523 1234
rect 11679 864 11691 1234
rect 11751 1008 11763 1234
rect 11967 240 11979 1234
rect 12135 432 12147 1234
rect 12231 888 12243 1234
rect 12327 1008 12339 1234
rect 12423 1056 12435 1234
rect 12831 1128 12843 1234
rect 11907 0 11919 34
rect 12855 24 12867 1234
rect 12975 432 12987 1234
rect 13791 288 13803 1234
rect 13983 768 13995 1234
rect 14007 240 14019 1234
rect 14103 744 14115 1234
rect 14175 360 14187 1234
rect 14199 744 14211 1234
rect 14223 312 14235 1234
rect 15231 504 15243 1234
rect 15471 696 15483 1234
rect 15567 384 15579 1234
rect 15663 696 15675 1234
rect 15711 504 15723 1234
rect 15975 648 15987 1234
rect 14811 0 14823 346
rect 16095 336 16107 1234
rect 16167 1224 16179 1234
rect 16191 648 16203 1234
rect 16263 1152 16275 1234
rect 16479 1128 16491 1234
rect 16575 480 16587 1234
rect 16275 0 16287 370
rect 16671 192 16683 1234
rect 16743 1152 16755 1234
rect 16767 1224 16779 1234
rect 16935 144 16947 1234
rect 16959 1128 16971 1234
rect 17103 768 17115 1234
rect 17847 984 17859 1234
rect 18111 696 18123 1234
rect 18159 696 18171 1234
rect 18207 1008 18219 1234
rect 17739 0 17751 466
rect 18279 264 18291 1234
rect 18495 1104 18507 1234
rect 18807 288 18819 1234
rect 18831 456 18843 1234
rect 18927 240 18939 1234
rect 19191 1152 19203 1234
rect 19239 648 19251 1234
rect 19263 888 19275 1234
rect 19455 1224 19467 1234
rect 19671 648 19683 1234
rect 19695 1200 19707 1234
rect 19743 912 19755 1234
rect 19815 1056 19827 1234
rect 20031 432 20043 1234
rect 20079 1176 20091 1234
rect 20103 600 20115 1234
rect 20367 672 20379 1234
rect 20463 1104 20475 1234
rect 20559 864 20571 1234
rect 20583 552 20595 1234
rect 20631 216 20643 1234
rect 17763 0 17775 106
rect 19227 0 19239 82
rect 20691 0 20703 1066
rect 20823 408 20835 1234
rect 20847 528 20859 1234
rect 20895 624 20907 1234
rect 21015 960 21027 1234
rect 21231 816 21243 1234
rect 21279 936 21291 1234
rect 21351 480 21363 1234
rect 21663 504 21675 1234
rect 21759 864 21771 1234
rect 21927 360 21939 1234
rect 21999 864 22011 1234
rect 22359 648 22371 1234
rect 22431 168 22443 1234
rect 22575 1128 22587 1234
rect 22647 576 22659 1234
rect 23007 864 23019 1234
rect 23175 1032 23187 1234
rect 23223 648 23235 1234
rect 23236 634 23254 648
rect 23235 0 23247 634
rect 23271 384 23283 1234
rect 23391 720 23403 1234
rect 23511 792 23523 1234
rect 23619 0 23631 826
rect 24543 696 24555 1234
rect 24591 648 24603 1234
rect 24711 648 24723 1234
rect 24711 144 24723 610
rect 24711 24 24723 58
rect 24735 48 24747 1114
rect 24759 72 24771 730
rect 24783 96 24795 850
rect 24807 120 24819 1090
rect 25359 0 25559 1234
rect 25613 131 25683 143
rect 25613 107 25683 119
rect 25613 83 25683 95
rect 25613 59 25683 71
rect 25613 35 25683 47
rect 25613 11 25683 23
use leftbuf leftbuf_1
timestamp 1386242881
transform 1 0 -1377 0 1 7275
box 0 0 1464 799
use nand3 g8075
timestamp 1386234893
transform 1 0 87 0 1 7275
box 0 0 120 799
use rowcrosser Rs1Sel_91_1_93_
timestamp 1386086759
transform 1 0 207 0 1 7275
box 0 0 48 799
use nand2 g7994
timestamp 1386234792
transform 1 0 255 0 1 7275
box 0 0 96 799
use nand3 g8032
timestamp 1386234893
transform 1 0 351 0 1 7275
box 0 0 120 799
use nand2 g7941
timestamp 1386234792
transform 1 0 471 0 1 7275
box 0 0 96 799
use nand3 g8197
timestamp 1386234893
transform 1 0 567 0 1 7275
box 0 0 120 799
use nand2 g8043
timestamp 1386234792
transform 1 0 687 0 1 7275
box 0 0 96 799
use nand3 g8112
timestamp 1386234893
transform 1 0 783 0 1 7275
box 0 0 120 799
use nand2 g8060
timestamp 1386234792
transform 1 0 903 0 1 7275
box 0 0 96 799
use nand3 g7942
timestamp 1386234893
transform 1 0 999 0 1 7275
box 0 0 120 799
use nor2 g8066
timestamp 1386235306
transform 1 0 1119 0 1 7275
box 0 0 120 799
use nand2 g8169
timestamp 1386234792
transform 1 0 1239 0 1 7275
box 0 0 96 799
use nand3 g7934
timestamp 1386234893
transform 1 0 1335 0 1 7275
box 0 0 120 799
use nand2 g8107
timestamp 1386234792
transform 1 0 1455 0 1 7275
box 0 0 96 799
use nand2 g8229
timestamp 1386234792
transform 1 0 1551 0 1 7275
box 0 0 96 799
use nand2 g7912
timestamp 1386234792
transform 1 0 1647 0 1 7275
box 0 0 96 799
use nand4 g8039
timestamp 1386234936
transform 1 0 1743 0 1 7275
box 0 0 144 799
use and2 g8046
timestamp 1386234845
transform 1 0 1887 0 1 7275
box 0 0 120 799
use nand3 g8123
timestamp 1386234893
transform 1 0 2007 0 1 7275
box 0 0 120 799
use and2 g8222
timestamp 1386234845
transform 1 0 2127 0 1 7275
box 0 0 120 799
use nand2 g8102
timestamp 1386234792
transform 1 0 2247 0 1 7275
box 0 0 96 799
use nor2 g8098
timestamp 1386235306
transform 1 0 2343 0 1 7275
box 0 0 120 799
use nand3 g8012
timestamp 1386234893
transform 1 0 2463 0 1 7275
box 0 0 120 799
use nor2 g8187
timestamp 1386235306
transform 1 0 2583 0 1 7275
box 0 0 120 799
use inv g7951
timestamp 1386238110
transform 1 0 2703 0 1 7275
box 0 0 120 799
use nand4 g8171
timestamp 1386234936
transform 1 0 2823 0 1 7275
box 0 0 144 799
use nand2 g8135
timestamp 1386234792
transform 1 0 2967 0 1 7275
box 0 0 96 799
use nand2 g8154
timestamp 1386234792
transform 1 0 3063 0 1 7275
box 0 0 96 799
use nor2 g8261
timestamp 1386235306
transform 1 0 3159 0 1 7275
box 0 0 120 799
use nand2 g8276
timestamp 1386234792
transform 1 0 3279 0 1 7275
box 0 0 96 799
use inv g8130
timestamp 1386238110
transform 1 0 3375 0 1 7275
box 0 0 120 799
use nand3 g8027
timestamp 1386234893
transform 1 0 3495 0 1 7275
box 0 0 120 799
use nand3 g8082
timestamp 1386234893
transform 1 0 3615 0 1 7275
box 0 0 120 799
use nand2 g8035
timestamp 1386234792
transform 1 0 3735 0 1 7275
box 0 0 96 799
use inv g8019
timestamp 1386238110
transform 1 0 3831 0 1 7275
box 0 0 120 799
use nand2 g8168
timestamp 1386234792
transform 1 0 3951 0 1 7275
box 0 0 96 799
use nand2 g8238
timestamp 1386234792
transform 1 0 4047 0 1 7275
box 0 0 96 799
use nand2 g7989
timestamp 1386234792
transform 1 0 4143 0 1 7275
box 0 0 96 799
use nand2 g8225
timestamp 1386234792
transform 1 0 4239 0 1 7275
box 0 0 96 799
use mux2 g8143
timestamp 1386235218
transform 1 0 4335 0 1 7275
box 0 0 192 799
use and2 g454
timestamp 1386234845
transform 1 0 4527 0 1 7275
box 0 0 120 799
use trisbuf g2
timestamp 1386237216
transform 1 0 4647 0 1 7275
box 0 0 216 799
use nand3 g8069
timestamp 1386234893
transform 1 0 4863 0 1 7275
box 0 0 120 799
use inv g8042
timestamp 1386238110
transform 1 0 4983 0 1 7275
box 0 0 120 799
use nand2 g8149
timestamp 1386234792
transform 1 0 5103 0 1 7275
box 0 0 96 799
use nand3 g7926
timestamp 1386234893
transform 1 0 5199 0 1 7275
box 0 0 120 799
use nand2 g8280
timestamp 1386234792
transform 1 0 5319 0 1 7275
box 0 0 96 799
use inv g7985
timestamp 1386238110
transform 1 0 5415 0 1 7275
box 0 0 120 799
use nand2 g8249
timestamp 1386234792
transform 1 0 5535 0 1 7275
box 0 0 96 799
use nand2 g8064
timestamp 1386234792
transform 1 0 5631 0 1 7275
box 0 0 96 799
use nor2 g8235
timestamp 1386235306
transform 1 0 5727 0 1 7275
box 0 0 120 799
use nand2 g8058
timestamp 1386234792
transform 1 0 5847 0 1 7275
box 0 0 96 799
use nand4 g7948
timestamp 1386234936
transform 1 0 5943 0 1 7275
box 0 0 144 799
use nand2 g8009
timestamp 1386234792
transform 1 0 6087 0 1 7275
box 0 0 96 799
use nand2 g8055
timestamp 1386234792
transform 1 0 6183 0 1 7275
box 0 0 96 799
use rowcrosser rowcrosser_0
timestamp 1386086759
transform 1 0 6279 0 1 7275
box 0 0 48 799
use nand2 g7939
timestamp 1386234792
transform 1 0 6327 0 1 7275
box 0 0 96 799
use nand3 g8088
timestamp 1386234893
transform 1 0 6423 0 1 7275
box 0 0 120 799
use nand2 g7960
timestamp 1386234792
transform 1 0 6543 0 1 7275
box 0 0 96 799
use nand2 g7947
timestamp 1386234792
transform 1 0 6639 0 1 7275
box 0 0 96 799
use nand2 g8214
timestamp 1386234792
transform 1 0 6735 0 1 7275
box 0 0 96 799
use and2 g8056
timestamp 1386234845
transform 1 0 6831 0 1 7275
box 0 0 120 799
use inv g8269
timestamp 1386238110
transform 1 0 6951 0 1 7275
box 0 0 120 799
use nor2 g8183
timestamp 1386235306
transform 1 0 7071 0 1 7275
box 0 0 120 799
use nand2 g8170
timestamp 1386234792
transform 1 0 7191 0 1 7275
box 0 0 96 799
use nand3 g8124
timestamp 1386234893
transform 1 0 7287 0 1 7275
box 0 0 120 799
use inv g8106
timestamp 1386238110
transform 1 0 7407 0 1 7275
box 0 0 120 799
use nor2 g8119
timestamp 1386235306
transform 1 0 7527 0 1 7275
box 0 0 120 799
use nand2 g8146
timestamp 1386234792
transform 1 0 7647 0 1 7275
box 0 0 96 799
use and2 g8127
timestamp 1386234845
transform 1 0 7743 0 1 7275
box 0 0 120 799
use nand2 g8155
timestamp 1386234792
transform 1 0 7863 0 1 7275
box 0 0 96 799
use nand2 g8033
timestamp 1386234792
transform 1 0 7959 0 1 7275
box 0 0 96 799
use nand3 g7921
timestamp 1386234893
transform 1 0 8055 0 1 7275
box 0 0 120 799
use nand2 g8252
timestamp 1386234792
transform 1 0 8175 0 1 7275
box 0 0 96 799
use nor2 g7978
timestamp 1386235306
transform 1 0 8271 0 1 7275
box 0 0 120 799
use nand3 g8244
timestamp 1386234893
transform 1 0 8391 0 1 7275
box 0 0 120 799
use and2 g7930
timestamp 1386234845
transform 1 0 8511 0 1 7275
box 0 0 120 799
use nand4 g7972
timestamp 1386234936
transform 1 0 8631 0 1 7275
box 0 0 144 799
use inv g8240
timestamp 1386238110
transform 1 0 8775 0 1 7275
box 0 0 120 799
use nor2 g8054
timestamp 1386235306
transform 1 0 8895 0 1 7275
box 0 0 120 799
use and2 g8139
timestamp 1386234845
transform 1 0 9015 0 1 7275
box 0 0 120 799
use nand2 g8023
timestamp 1386234792
transform 1 0 9135 0 1 7275
box 0 0 96 799
use nand2 g8118
timestamp 1386234792
transform 1 0 9231 0 1 7275
box 0 0 96 799
use nand2 g7981
timestamp 1386234792
transform 1 0 9327 0 1 7275
box 0 0 96 799
use nand4 g8111
timestamp 1386234936
transform 1 0 9423 0 1 7275
box 0 0 144 799
use inv g8120
timestamp 1386238110
transform 1 0 9567 0 1 7275
box 0 0 120 799
use nand2 g8091
timestamp 1386234792
transform 1 0 9687 0 1 7275
box 0 0 96 799
use nand2 g7918
timestamp 1386234792
transform 1 0 9783 0 1 7275
box 0 0 96 799
use nand4 g8134
timestamp 1386234936
transform 1 0 9879 0 1 7275
box 0 0 144 799
use mux2 g8050
timestamp 1386235218
transform 1 0 10023 0 1 7275
box 0 0 192 799
use nand3 g8218
timestamp 1386234893
transform 1 0 10215 0 1 7275
box 0 0 120 799
use nand2 g7995
timestamp 1386234792
transform 1 0 10335 0 1 7275
box 0 0 96 799
use nand2 g7945
timestamp 1386234792
transform 1 0 10431 0 1 7275
box 0 0 96 799
use nand2 g7964
timestamp 1386234792
transform 1 0 10527 0 1 7275
box 0 0 96 799
use nand3 g8198
timestamp 1386234893
transform 1 0 10623 0 1 7275
box 0 0 120 799
use nand2 g8199
timestamp 1386234792
transform 1 0 10743 0 1 7275
box 0 0 96 799
use nand2 g8221
timestamp 1386234792
transform 1 0 10839 0 1 7275
box 0 0 96 799
use nand2 g8220
timestamp 1386234792
transform 1 0 10935 0 1 7275
box 0 0 96 799
use nand3 g8230
timestamp 1386234893
transform 1 0 11031 0 1 7275
box 0 0 120 799
use nor2 g8271
timestamp 1386235306
transform 1 0 11151 0 1 7275
box 0 0 120 799
use inv g8004
timestamp 1386238110
transform 1 0 11271 0 1 7275
box 0 0 120 799
use nand4 g8074
timestamp 1386234936
transform 1 0 11391 0 1 7275
box 0 0 144 799
use nand2 g8209
timestamp 1386234792
transform 1 0 11535 0 1 7275
box 0 0 96 799
use and2 g8103
timestamp 1386234845
transform 1 0 11631 0 1 7275
box 0 0 120 799
use inv g8268
timestamp 1386238110
transform 1 0 11751 0 1 7275
box 0 0 120 799
use nand2 g8180
timestamp 1386234792
transform 1 0 11871 0 1 7275
box 0 0 96 799
use xor2 g8005
timestamp 1386237344
transform 1 0 11967 0 1 7275
box 0 0 192 799
use nand4 g8052
timestamp 1386234936
transform 1 0 12159 0 1 7275
box 0 0 144 799
use and2 g8136
timestamp 1386234845
transform 1 0 12303 0 1 7275
box 0 0 120 799
use nand2 g8110
timestamp 1386234792
transform 1 0 12423 0 1 7275
box 0 0 96 799
use nand2 g8153
timestamp 1386234792
transform 1 0 12519 0 1 7275
box 0 0 96 799
use inv StatusReg_reg_91_3_93_
timestamp 1386238110
transform 1 0 12615 0 1 7275
box 0 0 120 799
use scandtype g7922
timestamp 1386241841
transform 1 0 12735 0 1 7275
box 0 0 624 799
use nand4 stateSub_reg_91_2_93_
timestamp 1386234936
transform 1 0 13359 0 1 7275
box 0 0 144 799
use scandtype g7943
timestamp 1386241841
transform 1 0 13503 0 1 7275
box 0 0 624 799
use nand4 g8024
timestamp 1386234936
transform 1 0 14127 0 1 7275
box 0 0 144 799
use nand3 g8099
timestamp 1386234893
transform 1 0 14271 0 1 7275
box 0 0 120 799
use nand2 g8057
timestamp 1386234792
transform 1 0 14391 0 1 7275
box 0 0 96 799
use nor2 g8190
timestamp 1386235306
transform 1 0 14487 0 1 7275
box 0 0 120 799
use inv g8045
timestamp 1386238110
transform 1 0 14607 0 1 7275
box 0 0 120 799
use nand3 g7913
timestamp 1386234893
transform 1 0 14727 0 1 7275
box 0 0 120 799
use nand3 g8018
timestamp 1386234893
transform 1 0 14847 0 1 7275
box 0 0 120 799
use inv g8092
timestamp 1386238110
transform 1 0 14967 0 1 7275
box 0 0 120 799
use nor2 g8081
timestamp 1386235306
transform 1 0 15087 0 1 7275
box 0 0 120 799
use nand2 g8243
timestamp 1386234792
transform 1 0 15207 0 1 7275
box 0 0 96 799
use and2 g8234
timestamp 1386234845
transform 1 0 15303 0 1 7275
box 0 0 120 799
use nand2 StatusReg_reg_91_1_93_
timestamp 1386234792
transform 1 0 15423 0 1 7275
box 0 0 96 799
use scandtype g7933
timestamp 1386241841
transform 1 0 15519 0 1 7275
box 0 0 624 799
use nand2 g8213
timestamp 1386234792
transform 1 0 16143 0 1 7275
box 0 0 96 799
use nand2 g7963
timestamp 1386234792
transform 1 0 16239 0 1 7275
box 0 0 96 799
use nand2 g8096
timestamp 1386234792
transform 1 0 16335 0 1 7275
box 0 0 96 799
use nand2 g8212
timestamp 1386234792
transform 1 0 16431 0 1 7275
box 0 0 96 799
use nand3 g7911
timestamp 1386234893
transform 1 0 16527 0 1 7275
box 0 0 120 799
use nand4 g8015
timestamp 1386234936
transform 1 0 16647 0 1 7275
box 0 0 144 799
use nand4 g8084
timestamp 1386234936
transform 1 0 16791 0 1 7275
box 0 0 144 799
use and2 g8265
timestamp 1386234845
transform 1 0 16935 0 1 7275
box 0 0 120 799
use inv g8200
timestamp 1386238110
transform 1 0 17055 0 1 7275
box 0 0 120 799
use nand2 g8108
timestamp 1386234792
transform 1 0 17175 0 1 7275
box 0 0 96 799
use nand2 g8049
timestamp 1386234792
transform 1 0 17271 0 1 7275
box 0 0 96 799
use nand4 g8144
timestamp 1386234936
transform 1 0 17367 0 1 7275
box 0 0 144 799
use nand2 g8159
timestamp 1386234792
transform 1 0 17511 0 1 7275
box 0 0 96 799
use nor2 g8177
timestamp 1386235306
transform 1 0 17607 0 1 7275
box 0 0 120 799
use nand2 g7996
timestamp 1386234792
transform 1 0 17727 0 1 7275
box 0 0 96 799
use nand2 g8251
timestamp 1386234792
transform 1 0 17823 0 1 7275
box 0 0 96 799
use nand2 g8036
timestamp 1386234792
transform 1 0 17919 0 1 7275
box 0 0 96 799
use nand2 g8226
timestamp 1386234792
transform 1 0 18015 0 1 7275
box 0 0 96 799
use xor2 g7929
timestamp 1386237344
transform 1 0 18111 0 1 7275
box 0 0 192 799
use nor2 g7979
timestamp 1386235306
transform 1 0 18303 0 1 7275
box 0 0 120 799
use nand3 g8264
timestamp 1386234893
transform 1 0 18423 0 1 7275
box 0 0 120 799
use nand2 g7924
timestamp 1386234792
transform 1 0 18543 0 1 7275
box 0 0 96 799
use nand4 g8089
timestamp 1386234936
transform 1 0 18639 0 1 7275
box 0 0 144 799
use nand3 g8206
timestamp 1386234893
transform 1 0 18783 0 1 7275
box 0 0 120 799
use nand2 g8237
timestamp 1386234792
transform 1 0 18903 0 1 7275
box 0 0 96 799
use nand2 g8016
timestamp 1386234792
transform 1 0 18999 0 1 7275
box 0 0 96 799
use nand4 g8278
timestamp 1386234936
transform 1 0 19095 0 1 7275
box 0 0 144 799
use inv g8216
timestamp 1386238110
transform 1 0 19239 0 1 7275
box 0 0 120 799
use nand2 StatusReg_reg_91_0_93_
timestamp 1386234792
transform 1 0 19359 0 1 7275
box 0 0 96 799
use scandtype g8253
timestamp 1386241841
transform 1 0 19455 0 1 7275
box 0 0 624 799
use inv g8186
timestamp 1386238110
transform 1 0 20079 0 1 7275
box 0 0 120 799
use and2 g7946
timestamp 1386234845
transform 1 0 20199 0 1 7275
box 0 0 120 799
use nand2 g8090
timestamp 1386234792
transform 1 0 20319 0 1 7275
box 0 0 96 799
use nand3 g8195
timestamp 1386234893
transform 1 0 20415 0 1 7275
box 0 0 120 799
use and2 g8223
timestamp 1386234845
transform 1 0 20535 0 1 7275
box 0 0 120 799
use nand2 g8077
timestamp 1386234792
transform 1 0 20655 0 1 7275
box 0 0 96 799
use nand2 g8133
timestamp 1386234792
transform 1 0 20751 0 1 7275
box 0 0 96 799
use nand4 g7971
timestamp 1386234936
transform 1 0 20847 0 1 7275
box 0 0 144 799
use nand2 g8041
timestamp 1386234792
transform 1 0 20991 0 1 7275
box 0 0 96 799
use and2 g8002
timestamp 1386234845
transform 1 0 21087 0 1 7275
box 0 0 120 799
use nand3 g8128
timestamp 1386234893
transform 1 0 21207 0 1 7275
box 0 0 120 799
use nand2 g8029
timestamp 1386234792
transform 1 0 21327 0 1 7275
box 0 0 96 799
use nand2 g8100
timestamp 1386234792
transform 1 0 21423 0 1 7275
box 0 0 96 799
use and2 g8117
timestamp 1386234845
transform 1 0 21519 0 1 7275
box 0 0 120 799
use nand2 g8167
timestamp 1386234792
transform 1 0 21639 0 1 7275
box 0 0 96 799
use nand2 g7982
timestamp 1386234792
transform 1 0 21735 0 1 7275
box 0 0 96 799
use nand2 g8227
timestamp 1386234792
transform 1 0 21831 0 1 7275
box 0 0 96 799
use nand2 g8191
timestamp 1386234792
transform 1 0 21927 0 1 7275
box 0 0 96 799
use nand2 g7975
timestamp 1386234792
transform 1 0 22023 0 1 7275
box 0 0 96 799
use nand3 g8270
timestamp 1386234893
transform 1 0 22119 0 1 7275
box 0 0 120 799
use inv g8073
timestamp 1386238110
transform 1 0 22239 0 1 7275
box 0 0 120 799
use nor2 g7967
timestamp 1386235306
transform 1 0 22359 0 1 7275
box 0 0 120 799
use nand2 g7925
timestamp 1386234792
transform 1 0 22479 0 1 7275
box 0 0 96 799
use nand2 g8163
timestamp 1386234792
transform 1 0 22575 0 1 7275
box 0 0 96 799
use nand3 g7969
timestamp 1386234893
transform 1 0 22671 0 1 7275
box 0 0 120 799
use nand2 g8051
timestamp 1386234792
transform 1 0 22791 0 1 7275
box 0 0 96 799
use nand4 g8147
timestamp 1386234936
transform 1 0 22887 0 1 7275
box 0 0 144 799
use nand3 g7955
timestamp 1386234893
transform 1 0 23031 0 1 7275
box 0 0 120 799
use inv g7928
timestamp 1386238110
transform 1 0 23151 0 1 7275
box 0 0 120 799
use nand2 g8030
timestamp 1386234792
transform 1 0 23271 0 1 7275
box 0 0 96 799
use and2 g1
timestamp 1386234845
transform 1 0 23367 0 1 7275
box 0 0 120 799
use trisbuf g8217
timestamp 1386237216
transform 1 0 23487 0 1 7275
box 0 0 216 799
use inv g8248
timestamp 1386238110
transform 1 0 23703 0 1 7275
box 0 0 120 799
use and2 g8114
timestamp 1386234845
transform 1 0 23823 0 1 7275
box 0 0 120 799
use nand2 g8174
timestamp 1386234792
transform 1 0 23943 0 1 7275
box 0 0 96 799
use nand2 g8241
timestamp 1386234792
transform 1 0 24039 0 1 7275
box 0 0 96 799
use inv g8067
timestamp 1386238110
transform 1 0 24135 0 1 7275
box 0 0 120 799
use nand2 g7990
timestamp 1386234792
transform 1 0 24255 0 1 7275
box 0 0 96 799
use nand3 g8158
timestamp 1386234893
transform 1 0 24351 0 1 7275
box 0 0 120 799
use nand2 g8063
timestamp 1386234792
transform 1 0 24471 0 1 7275
box 0 0 96 799
use nand2 g8257
timestamp 1386234792
transform 1 0 24567 0 1 7275
box 0 0 96 799
use nand2 nME
timestamp 1386234792
transform 1 0 24663 0 1 7275
box 0 0 96 799
use rightend rightend_1
timestamp 1386235834
transform 1 0 25239 0 1 7275
box 0 0 320 799
use leftbuf leftbuf_0
timestamp 1386242881
transform 1 0 -1377 0 1 1234
box 0 0 1464 799
use nand3 stateSub_reg_91_0_93_
timestamp 1386234893
transform 1 0 87 0 1 1234
box 0 0 120 799
use rowcrosser PcSel_91_0_93_
timestamp 1386086759
transform 1 0 207 0 1 1234
box 0 0 48 799
use scandtype g8150
timestamp 1386241841
transform 1 0 255 0 1 1234
box 0 0 624 799
use rowcrosser IrWe
timestamp 1386086759
transform 1 0 879 0 1 1234
box 0 0 48 799
use nand2 g8020
timestamp 1386234792
transform 1 0 927 0 1 1234
box 0 0 96 799
use nand2 g8178
timestamp 1386234792
transform 1 0 1023 0 1 1234
box 0 0 96 799
use nand3 state_reg_91_1_93_
timestamp 1386234893
transform 1 0 1119 0 1 1234
box 0 0 120 799
use scandtype g8250
timestamp 1386241841
transform 1 0 1239 0 1 1234
box 0 0 624 799
use inv g8148
timestamp 1386238110
transform 1 0 1863 0 1 1234
box 0 0 120 799
use nand2 g7976
timestamp 1386234792
transform 1 0 1983 0 1 1234
box 0 0 96 799
use nand4 g7993
timestamp 1386234936
transform 1 0 2079 0 1 1234
box 0 0 144 799
use nand2 g8211
timestamp 1386234792
transform 1 0 2223 0 1 1234
box 0 0 96 799
use nand2 g8196
timestamp 1386234792
transform 1 0 2319 0 1 1234
box 0 0 96 799
use nand2 g8175
timestamp 1386234792
transform 1 0 2415 0 1 1234
box 0 0 96 799
use nand3 g8078
timestamp 1386234893
transform 1 0 2511 0 1 1234
box 0 0 120 799
use nand2 g8093
timestamp 1386234792
transform 1 0 2631 0 1 1234
box 0 0 96 799
use nand2 g7974
timestamp 1386234792
transform 1 0 2727 0 1 1234
box 0 0 96 799
use nand3 g8104
timestamp 1386234893
transform 1 0 2823 0 1 1234
box 0 0 120 799
use nand2 g7940
timestamp 1386234792
transform 1 0 2943 0 1 1234
box 0 0 96 799
use nand4 g8160
timestamp 1386234936
transform 1 0 3039 0 1 1234
box 0 0 144 799
use inv g8076
timestamp 1386238110
transform 1 0 3183 0 1 1234
box 0 0 120 799
use and2 g8161
timestamp 1386234845
transform 1 0 3303 0 1 1234
box 0 0 120 799
use nand2 StatusReg_reg_91_2_93_
timestamp 1386234792
transform 1 0 3423 0 1 1234
box 0 0 96 799
use scandtype g8224
timestamp 1386241841
transform 1 0 3519 0 1 1234
box 0 0 624 799
use rowcrosser Flags_91_0_93_
timestamp 1386086759
transform 1 0 4143 0 1 1234
box 0 0 48 799
use xor2 g8094
timestamp 1386237344
transform 1 0 4191 0 1 1234
box 0 0 192 799
use nor2 g8121
timestamp 1386235306
transform 1 0 4383 0 1 1234
box 0 0 120 799
use nand2 g8037
timestamp 1386234792
transform 1 0 4503 0 1 1234
box 0 0 96 799
use nand2 g8266
timestamp 1386234792
transform 1 0 4599 0 1 1234
box 0 0 96 799
use nand2 g8125
timestamp 1386234792
transform 1 0 4695 0 1 1234
box 0 0 96 799
use nand3 g7915
timestamp 1386234893
transform 1 0 4791 0 1 1234
box 0 0 120 799
use nand3 g8232
timestamp 1386234893
transform 1 0 4911 0 1 1234
box 0 0 120 799
use nor2 g8152
timestamp 1386235306
transform 1 0 5031 0 1 1234
box 0 0 120 799
use nand2 g8080
timestamp 1386234792
transform 1 0 5151 0 1 1234
box 0 0 96 799
use nand2 g7997
timestamp 1386234792
transform 1 0 5247 0 1 1234
box 0 0 96 799
use nand3 g8267
timestamp 1386234893
transform 1 0 5343 0 1 1234
box 0 0 120 799
use and2 g8282
timestamp 1386234845
transform 1 0 5463 0 1 1234
box 0 0 120 799
use inv g8274
timestamp 1386238110
transform 1 0 5583 0 1 1234
box 0 0 120 799
use inv g8236
timestamp 1386238110
transform 1 0 5703 0 1 1234
box 0 0 120 799
use inv g8101
timestamp 1386238110
transform 1 0 5823 0 1 1234
box 0 0 120 799
use inv g8011
timestamp 1386238110
transform 1 0 5943 0 1 1234
box 0 0 120 799
use nand4 g7919
timestamp 1386234936
transform 1 0 6063 0 1 1234
box 0 0 144 799
use nand4 g8185
timestamp 1386234936
transform 1 0 6207 0 1 1234
box 0 0 144 799
use nand2 IntReq_reg
timestamp 1386234792
transform 1 0 6351 0 1 1234
box 0 0 96 799
use scandtype g7927
timestamp 1386241841
transform 1 0 6447 0 1 1234
box 0 0 624 799
use rowcrosser LrEn
timestamp 1386086759
transform 1 0 7071 0 1 1234
box 0 0 48 799
use nand2 g8255
timestamp 1386234792
transform 1 0 7119 0 1 1234
box 0 0 96 799
use inv g8086
timestamp 1386238110
transform 1 0 7215 0 1 1234
box 0 0 120 799
use nor2 g7962
timestamp 1386235306
transform 1 0 7335 0 1 1234
box 0 0 120 799
use nor2 g8192
timestamp 1386235306
transform 1 0 7455 0 1 1234
box 0 0 120 799
use nand2 g7988
timestamp 1386234792
transform 1 0 7575 0 1 1234
box 0 0 96 799
use nand2 g8254
timestamp 1386234792
transform 1 0 7671 0 1 1234
box 0 0 96 799
use nand2 g8116
timestamp 1386234792
transform 1 0 7767 0 1 1234
box 0 0 96 799
use nand2 g8145
timestamp 1386234792
transform 1 0 7863 0 1 1234
box 0 0 96 799
use nor2 g8166
timestamp 1386235306
transform 1 0 7959 0 1 1234
box 0 0 120 799
use nand2 g8014
timestamp 1386234792
transform 1 0 8079 0 1 1234
box 0 0 96 799
use nand2 g7959
timestamp 1386234792
transform 1 0 8175 0 1 1234
box 0 0 96 799
use nand4 g8001
timestamp 1386234936
transform 1 0 8271 0 1 1234
box 0 0 144 799
use rowcrosser Flags_91_1_93_
timestamp 1386086759
transform 1 0 8415 0 1 1234
box 0 0 48 799
use nand3 g7998
timestamp 1386234893
transform 1 0 8463 0 1 1234
box 0 0 120 799
use and2 g7987
timestamp 1386234845
transform 1 0 8583 0 1 1234
box 0 0 120 799
use nand3 g8072
timestamp 1386234893
transform 1 0 8703 0 1 1234
box 0 0 120 799
use nand2 g7966
timestamp 1386234792
transform 1 0 8823 0 1 1234
box 0 0 96 799
use nand2 g8105
timestamp 1386234792
transform 1 0 8919 0 1 1234
box 0 0 96 799
use rowcrosser Flags_91_2_93_
timestamp 1386086759
transform 1 0 9015 0 1 1234
box 0 0 48 799
use inv g8259
timestamp 1386238110
transform 1 0 9063 0 1 1234
box 0 0 120 799
use nand2 g8122
timestamp 1386234792
transform 1 0 9183 0 1 1234
box 0 0 96 799
use nand2 g8129
timestamp 1386234792
transform 1 0 9279 0 1 1234
box 0 0 96 799
use nand2 g8059
timestamp 1386234792
transform 1 0 9375 0 1 1234
box 0 0 96 799
use nor2 g8097
timestamp 1386235306
transform 1 0 9471 0 1 1234
box 0 0 120 799
use inv g8062
timestamp 1386238110
transform 1 0 9591 0 1 1234
box 0 0 120 799
use nand2 g8025
timestamp 1386234792
transform 1 0 9711 0 1 1234
box 0 0 96 799
use nand3 g8247
timestamp 1386234893
transform 1 0 9807 0 1 1234
box 0 0 120 799
use rowcrosser ImmSel
timestamp 1386086759
transform 1 0 9927 0 1 1234
box 0 0 48 799
use nand2 g8263
timestamp 1386234792
transform 1 0 9975 0 1 1234
box 0 0 96 799
use nand2 g8256
timestamp 1386234792
transform 1 0 10071 0 1 1234
box 0 0 96 799
use nand2 g8087
timestamp 1386234792
transform 1 0 10167 0 1 1234
box 0 0 96 799
use nand3 g7970
timestamp 1386234893
transform 1 0 10263 0 1 1234
box 0 0 120 799
use nand2 g7932
timestamp 1386234792
transform 1 0 10383 0 1 1234
box 0 0 96 799
use nand2 g8286
timestamp 1386234792
transform 1 0 10479 0 1 1234
box 0 0 96 799
use inv g7991
timestamp 1386238110
transform 1 0 10575 0 1 1234
box 0 0 120 799
use nor2 g8137
timestamp 1386235306
transform 1 0 10695 0 1 1234
box 0 0 120 799
use rowcrosser AluEn
timestamp 1386086759
transform 1 0 10815 0 1 1234
box 0 0 48 799
use inv g8201
timestamp 1386238110
transform 1 0 10863 0 1 1234
box 0 0 120 799
use and2 g7952
timestamp 1386234845
transform 1 0 10983 0 1 1234
box 0 0 120 799
use nand3 g7936
timestamp 1386234893
transform 1 0 11103 0 1 1234
box 0 0 120 799
use nand3 g8242
timestamp 1386234893
transform 1 0 11223 0 1 1234
box 0 0 120 799
use nand2 g8207
timestamp 1386234792
transform 1 0 11343 0 1 1234
box 0 0 96 799
use nand2 g8044
timestamp 1386234792
transform 1 0 11439 0 1 1234
box 0 0 96 799
use nand3 g8006
timestamp 1386234893
transform 1 0 11535 0 1 1234
box 0 0 120 799
use nand3 g8173
timestamp 1386234893
transform 1 0 11655 0 1 1234
box 0 0 120 799
use and2 g7956
timestamp 1386234845
transform 1 0 11775 0 1 1234
box 0 0 120 799
use nand4 g8157
timestamp 1386234936
transform 1 0 11895 0 1 1234
box 0 0 144 799
use nand3 g8040
timestamp 1386234893
transform 1 0 12039 0 1 1234
box 0 0 120 799
use nand2 g8068
timestamp 1386234792
transform 1 0 12159 0 1 1234
box 0 0 96 799
use nand2 g8140
timestamp 1386234792
transform 1 0 12255 0 1 1234
box 0 0 96 799
use nand2 g8141
timestamp 1386234792
transform 1 0 12351 0 1 1234
box 0 0 96 799
use inv g452
timestamp 1386238110
transform 1 0 12447 0 1 1234
box 0 0 120 799
use trisbuf g8210
timestamp 1386237216
transform 1 0 12567 0 1 1234
box 0 0 216 799
use nand2 InISR_reg
timestamp 1386234792
transform 1 0 12783 0 1 1234
box 0 0 96 799
use scandtype g8003
timestamp 1386241841
transform 1 0 12879 0 1 1234
box 0 0 624 799
use nand3 g8203
timestamp 1386234893
transform 1 0 13503 0 1 1234
box 0 0 120 799
use nand2 g8065
timestamp 1386234792
transform 1 0 13623 0 1 1234
box 0 0 96 799
use nand2 g8113
timestamp 1386234792
transform 1 0 13719 0 1 1234
box 0 0 96 799
use inv g7977
timestamp 1386238110
transform 1 0 13815 0 1 1234
box 0 0 120 799
use nand3 g8070
timestamp 1386234893
transform 1 0 13935 0 1 1234
box 0 0 120 799
use nand2 g8038
timestamp 1386234792
transform 1 0 14055 0 1 1234
box 0 0 96 799
use nand2 IRQ2_reg
timestamp 1386234792
transform 1 0 14151 0 1 1234
box 0 0 96 799
use scandtype g8233
timestamp 1386241841
transform 1 0 14247 0 1 1234
box 0 0 624 799
use inv g7980
timestamp 1386238110
transform 1 0 14871 0 1 1234
box 0 0 120 799
use inv g7954
timestamp 1386238110
transform 1 0 14991 0 1 1234
box 0 0 120 799
use nand4 g8151
timestamp 1386234936
transform 1 0 15111 0 1 1234
box 0 0 144 799
use inv g7920
timestamp 1386238110
transform 1 0 15255 0 1 1234
box 0 0 120 799
use nand3 g8138
timestamp 1386234893
transform 1 0 15375 0 1 1234
box 0 0 120 799
use nand2 g7968
timestamp 1386234792
transform 1 0 15495 0 1 1234
box 0 0 96 799
use nand2 g8188
timestamp 1386234792
transform 1 0 15591 0 1 1234
box 0 0 96 799
use nand2 g8176
timestamp 1386234792
transform 1 0 15687 0 1 1234
box 0 0 96 799
use nand2 g8172
timestamp 1386234792
transform 1 0 15783 0 1 1234
box 0 0 96 799
use and2 g8026
timestamp 1386234845
transform 1 0 15879 0 1 1234
box 0 0 120 799
use nor2 g8031
timestamp 1386235306
transform 1 0 15999 0 1 1234
box 0 0 120 799
use nand2 g7935
timestamp 1386234792
transform 1 0 16119 0 1 1234
box 0 0 96 799
use nor2 g8162
timestamp 1386235306
transform 1 0 16215 0 1 1234
box 0 0 120 799
use nand2 g8095
timestamp 1386234792
transform 1 0 16335 0 1 1234
box 0 0 96 799
use nor2 g7950
timestamp 1386235306
transform 1 0 16431 0 1 1234
box 0 0 120 799
use nand2 g8008
timestamp 1386234792
transform 1 0 16551 0 1 1234
box 0 0 96 799
use nand4 g8013
timestamp 1386234936
transform 1 0 16647 0 1 1234
box 0 0 144 799
use inv g8126
timestamp 1386238110
transform 1 0 16791 0 1 1234
box 0 0 120 799
use nand2 g7984
timestamp 1386234792
transform 1 0 16911 0 1 1234
box 0 0 96 799
use nor2 IRQ1_reg
timestamp 1386235306
transform 1 0 17007 0 1 1234
box 0 0 120 799
use scandtype g7986
timestamp 1386241841
transform 1 0 17127 0 1 1234
box 0 0 624 799
use nand3 g8205
timestamp 1386234893
transform 1 0 17751 0 1 1234
box 0 0 120 799
use and2 g8164
timestamp 1386234845
transform 1 0 17871 0 1 1234
box 0 0 120 799
use nand2 g7949
timestamp 1386234792
transform 1 0 17991 0 1 1234
box 0 0 96 799
use nand2 g8017
timestamp 1386234792
transform 1 0 18087 0 1 1234
box 0 0 96 799
use nor2 g8010
timestamp 1386235306
transform 1 0 18183 0 1 1234
box 0 0 120 799
use and2 g8165
timestamp 1386234845
transform 1 0 18303 0 1 1234
box 0 0 120 799
use nand3 g8245
timestamp 1386234893
transform 1 0 18423 0 1 1234
box 0 0 120 799
use nand2 g8260
timestamp 1386234792
transform 1 0 18543 0 1 1234
box 0 0 96 799
use inv g8034
timestamp 1386238110
transform 1 0 18639 0 1 1234
box 0 0 120 799
use nand2 g8215
timestamp 1386234792
transform 1 0 18759 0 1 1234
box 0 0 96 799
use nand2 g8343
timestamp 1386234792
transform 1 0 18855 0 1 1234
box 0 0 96 799
use nand4 g8079
timestamp 1386234936
transform 1 0 18951 0 1 1234
box 0 0 144 799
use nand3 g7999
timestamp 1386234893
transform 1 0 19095 0 1 1234
box 0 0 120 799
use and2 g8239
timestamp 1386234845
transform 1 0 19215 0 1 1234
box 0 0 120 799
use nand2 g8007
timestamp 1386234792
transform 1 0 19335 0 1 1234
box 0 0 96 799
use inv g8262
timestamp 1386238110
transform 1 0 19431 0 1 1234
box 0 0 120 799
use nand2 g7965
timestamp 1386234792
transform 1 0 19551 0 1 1234
box 0 0 96 799
use and2 g8109
timestamp 1386234845
transform 1 0 19647 0 1 1234
box 0 0 120 799
use nand2 g8085
timestamp 1386234792
transform 1 0 19767 0 1 1234
box 0 0 96 799
use nand2 g7944
timestamp 1386234792
transform 1 0 19863 0 1 1234
box 0 0 96 799
use nand2 g8021
timestamp 1386234792
transform 1 0 19959 0 1 1234
box 0 0 96 799
use nor2 g7931
timestamp 1386235306
transform 1 0 20055 0 1 1234
box 0 0 120 799
use nand2 g8184
timestamp 1386234792
transform 1 0 20175 0 1 1234
box 0 0 96 799
use and2 g8132
timestamp 1386234845
transform 1 0 20271 0 1 1234
box 0 0 120 799
use nand3 g8219
timestamp 1386234893
transform 1 0 20391 0 1 1234
box 0 0 120 799
use nand2 g7916
timestamp 1386234792
transform 1 0 20511 0 1 1234
box 0 0 96 799
use rowcrosser PcEn
timestamp 1386086759
transform 1 0 20607 0 1 1234
box 0 0 48 799
use nand3 g8061
timestamp 1386234893
transform 1 0 20655 0 1 1234
box 0 0 120 799
use nand2 g8258
timestamp 1386234792
transform 1 0 20775 0 1 1234
box 0 0 96 799
use and2 g8115
timestamp 1386234845
transform 1 0 20871 0 1 1234
box 0 0 120 799
use inv g8202
timestamp 1386238110
transform 1 0 20991 0 1 1234
box 0 0 120 799
use nand2 g7973
timestamp 1386234792
transform 1 0 21111 0 1 1234
box 0 0 96 799
use nand3 g453
timestamp 1386234893
transform 1 0 21207 0 1 1234
box 0 0 120 799
use rowcrosser Flags_91_3_93_
timestamp 1386086759
transform 1 0 21327 0 1 1234
box 0 0 48 799
use trisbuf g8246
timestamp 1386237216
transform 1 0 21375 0 1 1234
box 0 0 216 799
use inv g8208
timestamp 1386238110
transform 1 0 21591 0 1 1234
box 0 0 120 799
use and2 g7958
timestamp 1386234845
transform 1 0 21711 0 1 1234
box 0 0 120 799
use nand3 g8156
timestamp 1386234893
transform 1 0 21831 0 1 1234
box 0 0 120 799
use nand2 g8231
timestamp 1386234792
transform 1 0 21951 0 1 1234
box 0 0 96 799
use inv g8047
timestamp 1386238110
transform 1 0 22047 0 1 1234
box 0 0 120 799
use nand3 g7992
timestamp 1386234893
transform 1 0 22167 0 1 1234
box 0 0 120 799
use nand2 g7957
timestamp 1386234792
transform 1 0 22287 0 1 1234
box 0 0 96 799
use nor2 g8179
timestamp 1386235306
transform 1 0 22383 0 1 1234
box 0 0 120 799
use mux2 g8022
timestamp 1386235218
transform 1 0 22503 0 1 1234
box 0 0 192 799
use nand2 g8193
timestamp 1386234792
transform 1 0 22695 0 1 1234
box 0 0 96 799
use nand2 g8071
timestamp 1386234792
transform 1 0 22791 0 1 1234
box 0 0 96 799
use nand2 g8285
timestamp 1386234792
transform 1 0 22887 0 1 1234
box 0 0 96 799
use inv g8083
timestamp 1386238110
transform 1 0 22983 0 1 1234
box 0 0 120 799
use nand2 g7953
timestamp 1386234792
transform 1 0 23103 0 1 1234
box 0 0 96 799
use rowcrosser PcWe
timestamp 1386086759
transform 1 0 23199 0 1 1234
box 0 0 48 799
use rowcrosser g7914
timestamp 1386086759
transform 1 0 23247 0 1 1234
box 0 0 48 799
use nand4 g8204
timestamp 1386234936
transform 1 0 23295 0 1 1234
box 0 0 144 799
use nand2 g8053
timestamp 1386234792
transform 1 0 23439 0 1 1234
box 0 0 96 799
use nand2 g8000
timestamp 1386234792
transform 1 0 23535 0 1 1234
box 0 0 96 799
use nand2 state_reg_91_0_93_
timestamp 1386234792
transform 1 0 23631 0 1 1234
box 0 0 96 799
use scandtype g8142
timestamp 1386241841
transform 1 0 23727 0 1 1234
box 0 0 624 799
use nor2 g7917
timestamp 1386235306
transform 1 0 24351 0 1 1234
box 0 0 120 799
use nand4 stateSub_reg_91_1_93_
timestamp 1386234936
transform 1 0 24471 0 1 1234
box 0 0 144 799
use scandtype LrSel
timestamp 1386241841
transform 1 0 24615 0 1 1234
box 0 0 624 799
use rightend rightend_0
timestamp 1386235834
transform 1 0 25239 0 1 1234
box 0 0 320 799
<< labels >>
rlabel m2contact 25269 6106 25269 6106 6 SysBus[1]
rlabel m2contact 25269 2170 25269 2170 6 SysBus[1]
rlabel m2contact 25245 5794 25245 5794 6 SysBus[0]
rlabel m2contact 25245 2146 25245 2146 6 SysBus[0]
rlabel m2contact 25221 4762 25221 4762 6 SysBus[3]
rlabel m2contact 25221 2122 25221 2122 6 SysBus[3]
rlabel m2contact 25197 2338 25197 2338 6 SysBus[2]
rlabel m2contact 25197 2098 25197 2098 6 SysBus[2]
rlabel m2contact 25173 5386 25173 5386 6 OpcodeCondIn[3]
rlabel m2contact 25173 2074 25173 2074 6 OpcodeCondIn[3]
rlabel m2contact 25149 2194 25149 2194 6 OpcodeCondIn[1]
rlabel m2contact 25149 2050 25149 2050 6 OpcodeCondIn[1]
rlabel m2contact 25125 5698 25125 5698 6 stateSub[1]
rlabel m2contact 25077 3322 25077 3322 6 n_163
rlabel m2contact 24741 5626 24741 5626 6 n_13
rlabel m2contact 24717 2794 24717 2794 6 n_39
rlabel m2contact 24693 5698 24693 5698 6 stateSub[1]
rlabel m2contact 24669 6658 24669 6658 6 n_302
rlabel m2contact 24669 3586 24669 3586 6 n_302
rlabel m2contact 24645 2362 24645 2362 6 n_218
rlabel m2contact 24621 7234 24621 7234 6 n_184
rlabel m2contact 24597 2482 24597 2482 6 n_217
rlabel m2contact 24573 3010 24573 3010 6 n_323
rlabel m2contact 24549 2674 24549 2674 6 n_88
rlabel m2contact 24525 3682 24525 3682 6 n_33
rlabel m2contact 24525 5050 24525 5050 6 n_132
rlabel m2contact 24501 4738 24501 4738 6 n_31
rlabel m2contact 24501 4858 24501 4858 6 n_268
rlabel m2contact 24477 7138 24477 7138 6 n_75
rlabel m2contact 24477 4666 24477 4666 6 n_75
rlabel m2contact 24453 6658 24453 6658 6 n_302
rlabel m2contact 24453 6634 24453 6634 6 n_113
rlabel m2contact 24429 5602 24429 5602 6 n_273
rlabel m2contact 24405 5962 24405 5962 6 n_274
rlabel m2contact 24405 5698 24405 5698 6 stateSub[1]
rlabel m2contact 24381 4666 24381 4666 6 n_75
rlabel m2contact 24381 5698 24381 5698 6 stateSub[1]
rlabel m2contact 24333 2818 24333 2818 6 n_159
rlabel m2contact 24309 5074 24309 5074 6 n_139
rlabel m2contact 24285 4546 24285 4546 6 n_101
rlabel m2contact 24237 4234 24237 4234 6 state[0]
rlabel m2contact 24213 3154 24213 3154 6 n_214
rlabel m2contact 24189 2794 24189 2794 6 n_39
rlabel m2contact 24165 2458 24165 2458 6 n_40
rlabel m2contact 24117 5770 24117 5770 6 n_64
rlabel m2contact 24093 5458 24093 5458 6 OpcodeCondIn[4]
rlabel m2contact 24069 7114 24069 7114 6 n_63
rlabel m2contact 24021 6706 24021 6706 6 n_222
rlabel m2contact 23997 5506 23997 5506 6 OpcodeCondIn[5]
rlabel m2contact 23973 2890 23973 2890 6 n_191
rlabel m2contact 23925 4210 23925 4210 6 n_148
rlabel m2contact 23877 4666 23877 4666 6 n_193
rlabel m2contact 23853 4234 23853 4234 6 state[0]
rlabel m2contact 23829 2410 23829 2410 6 n_344
rlabel m2contact 23781 3346 23781 3346 6 n_110
rlabel m2contact 23733 7138 23733 7138 6 n_75
rlabel m2contact 23709 7258 23709 7258 6 n_260
rlabel m2contact 23685 5842 23685 5842 6 n_253
rlabel m2contact 23661 4762 23661 4762 6 SysBus[3]
rlabel m2contact 23661 4714 23661 4714 6 n_209
rlabel m2contact 23637 4690 23637 4690 6 n_128
rlabel m2contact 23637 2554 23637 2554 6 n_128
rlabel m2contact 23613 5938 23613 5938 6 n_164
rlabel m2contact 23589 4810 23589 4810 6 n_237
rlabel m2contact 23589 3322 23589 3322 6 n_163
rlabel m2contact 23565 5818 23565 5818 6 n_165
rlabel m2contact 23541 5362 23541 5362 6 n_311
rlabel m2contact 23541 4594 23541 4594 6 n_311
rlabel m2contact 23517 4570 23517 4570 6 StatusReg[3]
rlabel m2contact 23493 6466 23493 6466 6 n_79
rlabel m2contact 23469 4498 23469 4498 6 Op1Sel
rlabel m2contact 23469 2962 23469 2962 6 n_80
rlabel m2contact 23445 4930 23445 4930 6 IrWe
rlabel m2contact 23445 4402 23445 4402 6 IrWe
rlabel m2contact 23421 4690 23421 4690 6 n_128
rlabel m2contact 23421 3778 23421 3778 6 nME
rlabel m2contact 23397 5842 23397 5842 6 n_253
rlabel m2contact 23373 5170 23373 5170 6 n_144
rlabel m2contact 23349 5362 23349 5362 6 n_311
rlabel m2contact 23349 5338 23349 5338 6 n_72
rlabel m2contact 23325 6154 23325 6154 6 n_312
rlabel m2contact 23325 5746 23325 5746 6 n_24
rlabel m2contact 23301 4762 23301 4762 6 SysBus[3]
rlabel m2contact 23277 4690 23277 4690 6 PcSel[0]
rlabel m2contact 23253 4762 23253 4762 6 n_95
rlabel m2contact 23253 2626 23253 2626 6 n_95
rlabel m2contact 23229 4402 23229 4402 6 IrWe
rlabel m2contact 23229 4426 23229 4426 6 n_355
rlabel m2contact 23205 6322 23205 6322 6 n_89
rlabel m2contact 23205 4042 23205 4042 6 n_89
rlabel m2contact 23181 4114 23181 4114 6 n_354
rlabel m2contact 23157 5386 23157 5386 6 OpcodeCondIn[3]
rlabel m2contact 23133 4762 23133 4762 6 n_95
rlabel m2contact 23133 2866 23133 2866 6 n_206
rlabel m2contact 23109 3490 23109 3490 6 n_182
rlabel m2contact 23085 6058 23085 6058 6 n_93
rlabel m2contact 23061 4042 23061 4042 6 n_89
rlabel m2contact 23061 4066 23061 4066 6 n_220
rlabel m2contact 23037 5602 23037 5602 6 n_273
rlabel m2contact 23037 4618 23037 4618 6 n_273
rlabel m2contact 23013 4714 23013 4714 6 n_209
rlabel m2contact 22989 4402 22989 4402 6 n_23
rlabel m2contact 22965 5722 22965 5722 6 n_141
rlabel m2contact 22965 2746 22965 2746 6 n_215
rlabel m2contact 22941 4522 22941 4522 6 n_48
rlabel m2contact 22941 3154 22941 3154 6 n_214
rlabel m2contact 22917 3802 22917 3802 6 n_231
rlabel m2contact 22917 6082 22917 6082 6 n_94
rlabel m2contact 22893 5962 22893 5962 6 n_274
rlabel m2contact 22893 3058 22893 3058 6 n_274
rlabel m2contact 22869 4690 22869 4690 6 PcSel[0]
rlabel m2contact 22869 3370 22869 3370 6 n_42
rlabel m2contact 22845 6946 22845 6946 6 n_293
rlabel m2contact 22845 4258 22845 4258 6 n_177
rlabel m2contact 22821 7258 22821 7258 6 n_260
rlabel m2contact 22821 7234 22821 7234 6 n_184
rlabel m2contact 22797 6322 22797 6322 6 n_89
rlabel m2contact 22797 4642 22797 4642 6 n_89
rlabel m2contact 22773 5314 22773 5314 6 n_68
rlabel m2contact 22773 3250 22773 3250 6 n_275
rlabel m2contact 22749 4618 22749 4618 6 n_273
rlabel m2contact 22749 4666 22749 4666 6 n_193
rlabel m2contact 22725 3058 22725 3058 6 n_274
rlabel m2contact 22725 3082 22725 3082 6 n_76
rlabel m2contact 22701 4474 22701 4474 6 n_197
rlabel m2contact 22677 5650 22677 5650 6 n_175
rlabel m2contact 22677 2218 22677 2218 6 n_175
rlabel m2contact 22653 3706 22653 3706 6 n_310
rlabel m2contact 22629 4642 22629 4642 6 n_89
rlabel m2contact 22629 6154 22629 6154 6 n_312
rlabel m2contact 22605 5794 22605 5794 6 SysBus[0]
rlabel m2contact 22581 5890 22581 5890 6 n_22
rlabel m2contact 22581 4618 22581 4618 6 n_22
rlabel m2contact 22557 4642 22557 4642 6 n_285
rlabel m2contact 22557 4090 22557 4090 6 n_234
rlabel m2contact 22533 5674 22533 5674 6 n_284
rlabel m2contact 22509 2530 22509 2530 6 InISR
rlabel m2contact 22485 3226 22485 3226 6 n_343
rlabel m2contact 22461 5842 22461 5842 6 n_253
rlabel m2contact 22437 4498 22437 4498 6 Op1Sel
rlabel m2contact 22413 5770 22413 5770 6 n_64
rlabel m2contact 22413 5578 22413 5578 6 n_329
rlabel m2contact 22389 6706 22389 6706 6 n_222
rlabel m2contact 22365 6946 22365 6946 6 n_293
rlabel m2contact 22365 4498 22365 4498 6 n_293
rlabel m2contact 22341 5386 22341 5386 6 OpcodeCondIn[3]
rlabel m2contact 22317 5650 22317 5650 6 n_175
rlabel m2contact 22317 5554 22317 5554 6 n_286
rlabel m2contact 22281 4786 22281 4786 6 n_248
rlabel m2contact 22281 3442 22281 3442 6 n_248
rlabel m2contact 22269 5386 22269 5386 6 OpcodeCondIn[3]
rlabel m2contact 22269 3106 22269 3106 6 n_223
rlabel m2contact 22245 4090 22245 4090 6 n_234
rlabel m2contact 22221 3538 22221 3538 6 n_202
rlabel m2contact 22221 4354 22221 4354 6 n_224
rlabel m2contact 22197 3442 22197 3442 6 n_248
rlabel m2contact 22197 3466 22197 3466 6 n_183
rlabel m2contact 22173 4450 22173 4450 6 n_178
rlabel m2contact 22149 2914 22149 2914 6 n_479
rlabel m2contact 22125 6466 22125 6466 6 n_79
rlabel m2contact 22101 4186 22101 4186 6 n_70
rlabel m2contact 22077 5890 22077 5890 6 n_22
rlabel m2contact 22077 5866 22077 5866 6 n_100
rlabel m2contact 22053 4066 22053 4066 6 n_220
rlabel m2contact 22029 5122 22029 5122 6 n_124
rlabel m2contact 22005 3946 22005 3946 6 n_47
rlabel m2contact 21981 4186 21981 4186 6 n_70
rlabel m2contact 21981 6010 21981 6010 6 n_45
rlabel m2contact 21957 5650 21957 5650 6 n_46
rlabel m2contact 21921 5770 21921 5770 6 n_195
rlabel m2contact 21921 5026 21921 5026 6 n_195
rlabel m2contact 21909 4498 21909 4498 6 n_293
rlabel m2contact 21909 6370 21909 6370 6 n_244
rlabel m2contact 21885 5938 21885 5938 6 n_164
rlabel m2contact 21885 5914 21885 5914 6 n_478
rlabel m2contact 21861 5770 21861 5770 6 n_195
rlabel m2contact 21861 5674 21861 5674 6 n_284
rlabel m2contact 21837 4906 21837 4906 6 n_87
rlabel m2contact 21837 2146 21837 2146 6 n_87
rlabel m2contact 21813 4906 21813 4906 6 n_87
rlabel m2contact 21813 4858 21813 4858 6 n_268
rlabel m2contact 21789 7090 21789 7090 6 n_6
rlabel m2contact 21765 4762 21765 4762 6 n_38
rlabel m2contact 21741 4090 21741 4090 6 n_234
rlabel m2contact 21717 6778 21717 6778 6 n_171
rlabel m2contact 21693 5266 21693 5266 6 n_109
rlabel m2contact 21669 2890 21669 2890 6 n_191
rlabel m2contact 21621 2122 21621 2122 6 n_26
rlabel m2contact 21621 6226 21621 6226 6 n_154
rlabel m2contact 21597 6106 21597 6106 6 SysBus[1]
rlabel m2contact 21597 3826 21597 3826 6 SysBus[1]
rlabel m2contact 21573 3874 21573 3874 6 n_264
rlabel m2contact 21549 3826 21549 3826 6 SysBus[1]
rlabel m2contact 21549 3850 21549 3850 6 n_168
rlabel m2contact 21501 6346 21501 6346 6 n_227
rlabel m2contact 21477 4858 21477 4858 6 n_268
rlabel m2contact 21477 4810 21477 4810 6 n_237
rlabel m2contact 21453 3610 21453 3610 6 n_226
rlabel m2contact 21417 4906 21417 4906 6 LrEn
rlabel m2contact 21417 2170 21417 2170 6 LrEn
rlabel m2contact 21405 2098 21405 2098 6 CFlag
rlabel m2contact 21405 6874 21405 6874 6 n_117
rlabel m2contact 21381 3514 21381 3514 6 stateSub[2]
rlabel m2contact 21357 2170 21357 2170 6 LrEn
rlabel m2contact 21357 2242 21357 2242 6 n_69
rlabel m2contact 21333 5362 21333 5362 6 n_174
rlabel m2contact 21333 3994 21333 3994 6 n_174
rlabel m2contact 21309 6970 21309 6970 6 n_228
rlabel m2contact 21285 5098 21285 5098 6 n_62
rlabel m2contact 21261 3994 21261 3994 6 n_174
rlabel m2contact 21261 4018 21261 4018 6 n_300
rlabel m2contact 21237 6658 21237 6658 6 n_134
rlabel m2contact 21213 6682 21213 6682 6 n_55
rlabel m2contact 21213 2842 21213 2842 6 n_55
rlabel m2contact 21189 2842 21189 2842 6 n_55
rlabel m2contact 21189 2938 21189 2938 6 n_212
rlabel m2contact 21165 3202 21165 3202 6 n_54
rlabel m2contact 21141 5530 21141 5530 6 n_130
rlabel m2contact 21141 3322 21141 3322 6 n_163
rlabel m2contact 21117 2170 21117 2170 6 n_179
rlabel m2contact 21093 4618 21093 4618 6 n_22
rlabel m2contact 21093 4138 21093 4138 6 n_22
rlabel m2contact 21069 4906 21069 4906 6 LrEn
rlabel m2contact 21069 4834 21069 4834 6 n_267
rlabel m2contact 21045 4978 21045 4978 6 n_235
rlabel m2contact 21021 5914 21021 5914 6 n_478
rlabel m2contact 20997 6610 20997 6610 6 OpcodeCondIn[0]
rlabel m2contact 20997 3442 20997 3442 6 OpcodeCondIn[0]
rlabel m2contact 20973 4138 20973 4138 6 n_22
rlabel m2contact 20973 4162 20973 4162 6 n_99
rlabel m2contact 20949 2218 20949 2218 6 n_175
rlabel m2contact 20925 2194 20925 2194 6 OpcodeCondIn[1]
rlabel m2contact 20925 6418 20925 6418 6 n_120
rlabel m2contact 20901 3442 20901 3442 6 OpcodeCondIn[0]
rlabel m2contact 20901 3514 20901 3514 6 stateSub[2]
rlabel m2contact 20877 4954 20877 4954 6 n_172
rlabel m2contact 20841 4690 20841 4690 6 n_76
rlabel m2contact 20841 3082 20841 3082 6 n_76
rlabel m2contact 20829 5146 20829 5146 6 n_205
rlabel m2contact 20805 4714 20805 4714 6 n_92
rlabel m2contact 20805 3514 20805 3514 6 stateSub[2]
rlabel m2contact 20781 2866 20781 2866 6 n_206
rlabel m2contact 20757 5482 20757 5482 6 n_368
rlabel m2contact 20733 4594 20733 4594 6 n_311
rlabel m2contact 20733 4906 20733 4906 6 n_49
rlabel m2contact 20709 7234 20709 7234 6 n_184
rlabel m2contact 20709 6274 20709 6274 6 n_345
rlabel m2contact 20685 4690 20685 4690 6 n_76
rlabel m2contact 20685 3298 20685 3298 6 n_305
rlabel m2contact 20661 5866 20661 5866 6 n_100
rlabel m2contact 20661 4594 20661 4594 6 n_100
rlabel m2contact 20637 5194 20637 5194 6 Flags[1]
rlabel m2contact 20637 5290 20637 5290 6 n_105
rlabel m2contact 20613 4690 20613 4690 6 n_182
rlabel m2contact 20613 3490 20613 3490 6 n_182
rlabel m2contact 20589 2794 20589 2794 6 n_39
rlabel m2contact 20565 4474 20565 4474 6 n_197
rlabel m2contact 20541 5410 20541 5410 6 n_11
rlabel m2contact 20517 3034 20517 3034 6 n_156
rlabel m2contact 20493 4546 20493 4546 6 n_101
rlabel m2contact 20493 4786 20493 4786 6 n_248
rlabel m2contact 20469 7018 20469 7018 6 n_161
rlabel m2contact 20445 4594 20445 4594 6 n_100
rlabel m2contact 20445 5002 20445 5002 6 n_152
rlabel m2contact 20421 4858 20421 4858 6 n_268
rlabel m2contact 20397 7210 20397 7210 6 n_352
rlabel m2contact 20373 5194 20373 5194 6 Flags[1]
rlabel m2contact 20349 6250 20349 6250 6 n_351
rlabel m2contact 20325 4066 20325 4066 6 n_220
rlabel m2contact 20301 7114 20301 7114 6 n_63
rlabel m2contact 20301 6466 20301 6466 6 n_79
rlabel m2contact 20277 5890 20277 5890 6 n_175
rlabel m2contact 20277 2218 20277 2218 6 n_175
rlabel m2contact 20253 4690 20253 4690 6 n_182
rlabel m2contact 20253 3562 20253 3562 6 n_309
rlabel m2contact 20229 5890 20229 5890 6 n_175
rlabel m2contact 20229 5770 20229 5770 6 StatusReg[0]
rlabel m2contact 20205 4546 20205 4546 6 n_307
rlabel m2contact 20181 5242 20181 5242 6 n_257
rlabel m2contact 20181 3922 20181 3922 6 n_257
rlabel m2contact 20157 3922 20157 3922 6 n_257
rlabel m2contact 20157 3970 20157 3970 6 n_249
rlabel m2contact 20109 2266 20109 2266 6 n_44
rlabel m2contact 20025 4690 20025 4690 6 n_477
rlabel m2contact 20025 3922 20025 3922 6 n_477
rlabel m2contact 20013 3130 20013 3130 6 n_334
rlabel m2contact 19989 4642 19989 4642 6 n_285
rlabel m2contact 19965 5770 19965 5770 6 StatusReg[0]
rlabel m2contact 19941 6490 19941 6490 6 n_236
rlabel m2contact 19917 4690 19917 4690 6 n_477
rlabel m2contact 19917 4090 19917 4090 6 n_234
rlabel m2contact 19893 5434 19893 5434 6 n_240
rlabel m2contact 19845 7066 19845 7066 6 n_173
rlabel m2contact 19797 2890 19797 2890 6 n_191
rlabel m2contact 19629 2842 19629 2842 6 n_32
rlabel m2contact 19605 4234 19605 4234 6 state[0]
rlabel m2contact 19581 3274 19581 3274 6 state[1]
rlabel m2contact 19557 3730 19557 3730 6 n_360
rlabel m2contact 19509 3418 19509 3418 6 n_288
rlabel m2contact 19473 5890 19473 5890 6 n_44
rlabel m2contact 19473 2266 19473 2266 6 n_44
rlabel m2contact 19449 4690 19449 4690 6 n_9
rlabel m2contact 19449 2074 19449 2074 6 n_9
rlabel m2contact 19437 4714 19437 4714 6 n_92
rlabel m2contact 19413 2074 19413 2074 6 n_9
rlabel m2contact 19413 2122 19413 2122 6 n_26
rlabel m2contact 19389 5890 19389 5890 6 n_44
rlabel m2contact 19389 5386 19389 5386 6 OpcodeCondIn[3]
rlabel m2contact 19365 2506 19365 2506 6 n_19
rlabel m2contact 19341 6898 19341 6898 6 n_277
rlabel m2contact 19341 4642 19341 4642 6 n_277
rlabel m2contact 19317 4642 19317 4642 6 n_277
rlabel m2contact 19317 6802 19317 6802 6 n_20
rlabel m2contact 19269 5458 19269 5458 6 OpcodeCondIn[4]
rlabel m2contact 19245 7234 19245 7234 6 n_184
rlabel m2contact 19245 4594 19245 4594 6 n_184
rlabel m2contact 19221 5194 19221 5194 6 n_131
rlabel m2contact 19197 5386 19197 5386 6 OpcodeCondIn[3]
rlabel m2contact 19173 4642 19173 4642 6 n_65
rlabel m2contact 19173 2218 19173 2218 6 n_175
rlabel m2contact 19149 5698 19149 5698 6 stateSub[1]
rlabel m2contact 19149 3850 19149 3850 6 n_168
rlabel m2contact 19125 4594 19125 4594 6 n_184
rlabel m2contact 19125 4954 19125 4954 6 n_172
rlabel m2contact 19101 6322 19101 6322 6 n_89
rlabel m2contact 19101 2434 19101 2434 6 n_89
rlabel m2contact 19077 2914 19077 2914 6 n_479
rlabel m2contact 19077 2962 19077 2962 6 n_80
rlabel m2contact 19053 6610 19053 6610 6 OpcodeCondIn[0]
rlabel m2contact 19053 4090 19053 4090 6 n_234
rlabel m2contact 19029 2434 19029 2434 6 n_89
rlabel m2contact 19029 2578 19029 2578 6 n_10
rlabel m2contact 19005 4234 19005 4234 6 state[0]
rlabel m2contact 18981 4762 18981 4762 6 n_38
rlabel m2contact 18981 3394 18981 3394 6 stateSub[0]
rlabel m2contact 18957 4690 18957 4690 6 n_9
rlabel m2contact 18933 2266 18933 2266 6 n_44
rlabel m2contact 18909 3394 18909 3394 6 stateSub[0]
rlabel m2contact 18885 6178 18885 6178 6 n_199
rlabel m2contact 18885 3082 18885 3082 6 n_76
rlabel m2contact 18861 4690 18861 4690 6 n_190
rlabel m2contact 18837 2890 18837 2890 6 n_191
rlabel m2contact 18813 5122 18813 5122 6 n_124
rlabel m2contact 18789 4594 18789 4594 6 n_136
rlabel m2contact 18765 5890 18765 5890 6 n_317
rlabel m2contact 18765 2650 18765 2650 6 n_317
rlabel m2contact 18741 5218 18741 5218 6 n_7
rlabel m2contact 18717 6994 18717 6994 6 n_254
rlabel m2contact 18717 4090 18717 4090 6 n_234
rlabel m2contact 18693 6586 18693 6586 6 n_122
rlabel m2contact 18669 5890 18669 5890 6 n_317
rlabel m2contact 18669 5410 18669 5410 6 n_11
rlabel m2contact 18621 5602 18621 5602 6 n_273
rlabel m2contact 18621 4762 18621 4762 6 n_16
rlabel m2contact 18597 4498 18597 4498 6 OpcodeCondIn[2]
rlabel m2contact 18597 3658 18597 3658 6 n_29
rlabel m2contact 18573 5386 18573 5386 6 OpcodeCondIn[3]
rlabel m2contact 18573 4234 18573 4234 6 state[0]
rlabel m2contact 18549 5866 18549 5866 6 n_100
rlabel m2contact 18549 3178 18549 3178 6 n_100
rlabel m2contact 18525 5578 18525 5578 6 n_329
rlabel m2contact 18525 4522 18525 4522 6 n_48
rlabel m2contact 18501 4138 18501 4138 6 n_328
rlabel m2contact 18477 3922 18477 3922 6 n_477
rlabel m2contact 18477 3994 18477 3994 6 n_251
rlabel m2contact 18453 3178 18453 3178 6 n_100
rlabel m2contact 18453 3442 18453 3442 6 n_233
rlabel m2contact 18429 7162 18429 7162 6 n_238
rlabel m2contact 18429 4522 18429 4522 6 n_238
rlabel m2contact 18405 4522 18405 4522 6 n_238
rlabel m2contact 18405 6730 18405 6730 6 n_340
rlabel m2contact 18357 6562 18357 6562 6 PcSel[2]
rlabel m2contact 18357 4666 18357 4666 6 n_193
rlabel m2contact 18333 6850 18333 6850 6 n_314
rlabel m2contact 18333 6298 18333 6298 6 n_194
rlabel m2contact 18261 6922 18261 6922 6 n_18
rlabel m2contact 18237 5698 18237 5698 6 stateSub[1]
rlabel m2contact 18165 5386 18165 5386 6 OpcodeCondIn[3]
rlabel m2contact 18141 6826 18141 6826 6 OpcodeCondIn[7]
rlabel m2contact 18141 5698 18141 5698 6 stateSub[1]
rlabel m2contact 18117 7018 18117 7018 6 n_161
rlabel m2contact 18117 3178 18117 3178 6 n_161
rlabel m2contact 18093 4378 18093 4378 6 n_270
rlabel m2contact 18069 4138 18069 4138 6 n_328
rlabel m2contact 18069 4786 18069 4786 6 n_248
rlabel m2contact 18045 2314 18045 2314 6 n_51
rlabel m2contact 18045 5842 18045 5842 6 n_253
rlabel m2contact 18021 3346 18021 3346 6 n_110
rlabel m2contact 17997 3202 17997 3202 6 n_54
rlabel m2contact 17973 3178 17973 3178 6 n_161
rlabel m2contact 17973 5386 17973 5386 6 OpcodeCondIn[3]
rlabel m2contact 17949 3874 17949 3874 6 n_264
rlabel m2contact 17925 5698 17925 5698 6 stateSub[1]
rlabel m2contact 17901 5362 17901 5362 6 n_174
rlabel m2contact 17901 4210 17901 4210 6 n_148
rlabel m2contact 17877 4234 17877 4234 6 state[0]
rlabel m2contact 17853 5194 17853 5194 6 n_131
rlabel m2contact 17829 4066 17829 4066 6 n_220
rlabel m2contact 17805 6538 17805 6538 6 n_145
rlabel m2contact 17805 6298 17805 6298 6 n_194
rlabel m2contact 17781 3178 17781 3178 6 n_161
rlabel m2contact 17781 3514 17781 3514 6 stateSub[2]
rlabel m2contact 17757 5290 17757 5290 6 n_105
rlabel m2contact 17709 4930 17709 4930 6 IrWe
rlabel m2contact 17685 5578 17685 5578 6 IRQ1
rlabel m2contact 17685 2986 17685 2986 6 IRQ1
rlabel m2contact 17661 3010 17661 3010 6 n_323
rlabel m2contact 17637 2986 17637 2986 6 IRQ1
rlabel m2contact 17637 3058 17637 3058 6 n_34
rlabel m2contact 17589 6754 17589 6754 6 n_104
rlabel m2contact 17565 2218 17565 2218 6 n_175
rlabel m2contact 17541 4930 17541 4930 6 n_56
rlabel m2contact 17493 5170 17493 5170 6 n_144
rlabel m2contact 17469 6826 17469 6826 6 OpcodeCondIn[7]
rlabel m2contact 17445 5698 17445 5698 6 stateSub[1]
rlabel m2contact 17421 4234 17421 4234 6 state[0]
rlabel m2contact 17397 6514 17397 6514 6 n_66
rlabel m2contact 17349 6034 17349 6034 6 n_125
rlabel m2contact 17325 5122 17325 5122 6 n_124
rlabel m2contact 17301 6418 17301 6418 6 n_120
rlabel m2contact 17277 7186 17277 7186 6 n_5
rlabel m2contact 17277 3178 17277 3178 6 n_5
rlabel m2contact 17253 4930 17253 4930 6 n_56
rlabel m2contact 17229 3178 17229 3178 6 n_5
rlabel m2contact 17229 3322 17229 3322 6 n_163
rlabel m2contact 17205 4762 17205 4762 6 n_16
rlabel m2contact 17133 4330 17133 4330 6 n_12
rlabel m2contact 17109 5194 17109 5194 6 n_226
rlabel m2contact 17109 3610 17109 3610 6 n_226
rlabel m2contact 17085 3010 17085 3010 6 n_323
rlabel m2contact 17061 7162 17061 7162 6 n_238
rlabel m2contact 17037 5194 17037 5194 6 n_226
rlabel m2contact 17037 5170 17037 5170 6 n_278
rlabel m2contact 17013 5602 17013 5602 6 n_261
rlabel m2contact 17013 3922 17013 3922 6 n_261
rlabel m2contact 16989 4522 16989 4522 6 n_129
rlabel m2contact 16989 4042 16989 4042 6 n_147
rlabel m2contact 16965 3538 16965 3538 6 n_202
rlabel m2contact 16929 4282 16929 4282 6 n_321
rlabel m2contact 16929 2986 16929 2986 6 n_321
rlabel m2contact 16917 4930 16917 4930 6 n_167
rlabel m2contact 16893 4498 16893 4498 6 OpcodeCondIn[2]
rlabel m2contact 16869 3922 16869 3922 6 n_261
rlabel m2contact 16869 4306 16869 4306 6 n_192
rlabel m2contact 16845 3850 16845 3850 6 n_168
rlabel m2contact 16821 2986 16821 2986 6 n_321
rlabel m2contact 16821 3178 16821 3178 6 n_245
rlabel m2contact 16749 3130 16749 3130 6 n_334
rlabel m2contact 16725 3034 16725 3034 6 n_156
rlabel m2contact 16725 3634 16725 3634 6 n_338
rlabel m2contact 16701 6394 16701 6394 6 n_243
rlabel m2contact 16701 5938 16701 5938 6 n_242
rlabel m2contact 16677 4282 16677 4282 6 n_321
rlabel m2contact 16629 4738 16629 4738 6 n_31
rlabel m2contact 16629 3922 16629 3922 6 n_290
rlabel m2contact 16605 4666 16605 4666 6 n_193
rlabel m2contact 16605 4234 16605 4234 6 state[0]
rlabel m2contact 16581 4258 16581 4258 6 n_177
rlabel m2contact 16557 3394 16557 3394 6 stateSub[0]
rlabel m2contact 16533 3538 16533 3538 6 n_202
rlabel m2contact 16509 3826 16509 3826 6 n_126
rlabel m2contact 16485 4858 16485 4858 6 n_268
rlabel m2contact 16461 7042 16461 7042 6 n_71
rlabel m2contact 16461 2914 16461 2914 6 n_155
rlabel m2contact 16437 4738 16437 4738 6 n_169
rlabel m2contact 16437 3754 16437 3754 6 n_169
rlabel m2contact 16413 2242 16413 2242 6 n_69
rlabel m2contact 16413 2290 16413 2290 6 WdSel
rlabel m2contact 16389 4738 16389 4738 6 n_169
rlabel m2contact 16389 4474 16389 4474 6 n_197
rlabel m2contact 16365 3898 16365 3898 6 n_266
rlabel m2contact 16365 2650 16365 2650 6 n_317
rlabel m2contact 16317 3634 16317 3634 6 n_338
rlabel m2contact 16317 5122 16317 5122 6 n_52
rlabel m2contact 16293 3514 16293 3514 6 stateSub[2]
rlabel m2contact 16269 2290 16269 2290 6 WdSel
rlabel m2contact 16269 2314 16269 2314 6 n_51
rlabel m2contact 16245 2986 16245 2986 6 n_316
rlabel m2contact 16221 2602 16221 2602 6 n_306
rlabel m2contact 16197 2722 16197 2722 6 StatusReg[2]
rlabel m2contact 16173 4546 16173 4546 6 n_307
rlabel m2contact 16149 5434 16149 5434 6 n_240
rlabel m2contact 16077 4762 16077 4762 6 CFlag
rlabel m2contact 16077 2098 16077 2098 6 CFlag
rlabel m2contact 16053 3202 16053 3202 6 n_54
rlabel m2contact 16029 4762 16029 4762 6 CFlag
rlabel m2contact 16029 4738 16029 4738 6 n_298
rlabel m2contact 15933 5050 15933 5050 6 n_132
rlabel m2contact 15909 3946 15909 3946 6 n_47
rlabel m2contact 15861 2386 15861 2386 6 n_61
rlabel m2contact 15837 4954 15837 4954 6 n_172
rlabel m2contact 15813 7114 15813 7114 6 n_63
rlabel m2contact 15765 5194 15765 5194 6 n_82
rlabel m2contact 15741 6322 15741 6322 6 n_89
rlabel m2contact 15645 2650 15645 2650 6 n_317
rlabel m2contact 15621 7258 15621 7258 6 n_361
rlabel m2contact 15621 5362 15621 5362 6 n_282
rlabel m2contact 15549 2506 15549 2506 6 n_19
rlabel m2contact 15525 4858 15525 4858 6 n_268
rlabel m2contact 15501 6442 15501 6442 6 n_21
rlabel m2contact 15477 2506 15477 2506 6 n_19
rlabel m2contact 15453 4138 15453 4138 6 n_328
rlabel m2contact 15453 6802 15453 6802 6 n_20
rlabel m2contact 15429 4426 15429 4426 6 n_355
rlabel m2contact 15405 7234 15405 7234 6 n_184
rlabel m2contact 15405 2770 15405 2770 6 n_362
rlabel m2contact 15357 3322 15357 3322 6 n_163
rlabel m2contact 15333 4522 15333 4522 6 n_129
rlabel m2contact 15333 4666 15333 4666 6 n_193
rlabel m2contact 15297 4762 15297 4762 6 n_206
rlabel m2contact 15297 2866 15297 2866 6 n_206
rlabel m2contact 15285 6130 15285 6130 6 n_213
rlabel m2contact 15285 2554 15285 2554 6 n_128
rlabel m2contact 15261 6946 15261 6946 6 n_293
rlabel m2contact 15237 5890 15237 5890 6 IntReq
rlabel m2contact 15213 3130 15213 3130 6 n_334
rlabel m2contact 15189 4762 15189 4762 6 n_206
rlabel m2contact 15189 4738 15189 4738 6 n_298
rlabel m2contact 15165 5986 15165 5986 6 n_232
rlabel m2contact 15141 5506 15141 5506 6 OpcodeCondIn[5]
rlabel m2contact 15141 4762 15141 4762 6 n_363
rlabel m2contact 15117 2914 15117 2914 6 n_155
rlabel m2contact 15069 2434 15069 2434 6 n_336
rlabel m2contact 15045 3034 15045 3034 6 n_287
rlabel m2contact 15021 6250 15021 6250 6 n_351
rlabel m2contact 14997 5554 14997 5554 6 n_286
rlabel m2contact 14949 7258 14949 7258 6 n_361
rlabel m2contact 14949 4954 14949 4954 6 n_172
rlabel m2contact 14925 6202 14925 6202 6 n_315
rlabel m2contact 14901 7210 14901 7210 6 n_352
rlabel m2contact 14901 6442 14901 6442 6 n_21
rlabel m2contact 14877 2074 14877 2074 6 n_308
rlabel m2contact 14829 4138 14829 4138 6 n_185
rlabel m2contact 14805 3394 14805 3394 6 stateSub[0]
rlabel m2contact 14781 5818 14781 5818 6 n_165
rlabel m2contact 14757 7234 14757 7234 6 n_184
rlabel m2contact 14757 7210 14757 7210 6 IRQ2
rlabel m2contact 14709 2698 14709 2698 6 n_473
rlabel m2contact 14685 4786 14685 4786 6 n_248
rlabel m2contact 14637 4186 14637 4186 6 n_70
rlabel m2contact 14589 3946 14589 3946 6 n_250
rlabel m2contact 14541 5458 14541 5458 6 OpcodeCondIn[4]
rlabel m2contact 14517 6706 14517 6706 6 n_222
rlabel m2contact 14469 4426 14469 4426 6 n_138
rlabel m2contact 14445 4522 14445 4522 6 n_86
rlabel m2contact 14421 6754 14421 6754 6 n_104
rlabel m2contact 14385 5578 14385 5578 6 IRQ1
rlabel m2contact 14385 2290 14385 2290 6 IRQ1
rlabel m2contact 14373 5986 14373 5986 6 n_232
rlabel m2contact 14349 2290 14349 2290 6 IRQ1
rlabel m2contact 14349 3394 14349 3394 6 stateSub[0]
rlabel m2contact 14325 3802 14325 3802 6 n_231
rlabel m2contact 14301 2242 14301 2242 6 n_91
rlabel m2contact 14229 3130 14229 3130 6 n_334
rlabel m2contact 14205 5986 14205 5986 6 n_291
rlabel m2contact 14181 6178 14181 6178 6 n_199
rlabel m2contact 14157 4282 14157 4282 6 n_321
rlabel m2contact 14133 5938 14133 5938 6 n_242
rlabel m2contact 14085 3802 14085 3802 6 n_231
rlabel m2contact 14037 3634 14037 3634 6 nWE
rlabel m2contact 14013 3514 14013 3514 6 stateSub[2]
rlabel m2contact 13965 2362 13965 2362 6 n_218
rlabel m2contact 13965 4258 13965 4258 6 n_177
rlabel m2contact 13893 5434 13893 5434 6 n_240
rlabel m2contact 13845 6706 13845 6706 6 n_222
rlabel m2contact 13773 2674 13773 2674 6 n_88
rlabel m2contact 13749 3826 13749 3826 6 n_126
rlabel m2contact 13701 4402 13701 4402 6 n_23
rlabel m2contact 13677 4618 13677 4618 6 n_22
rlabel m2contact 13653 5770 13653 5770 6 StatusReg[0]
rlabel m2contact 13605 6754 13605 6754 6 n_304
rlabel m2contact 13605 5362 13605 5362 6 n_282
rlabel m2contact 13581 2362 13581 2362 6 n_200
rlabel m2contact 13557 3514 13557 3514 6 stateSub[2]
rlabel m2contact 13533 4234 13533 4234 6 state[0]
rlabel m2contact 13461 5626 13461 5626 6 n_13
rlabel m2contact 13437 4402 13437 4402 6 n_303
rlabel m2contact 13413 5122 13413 5122 6 n_52
rlabel m2contact 13389 2530 13389 2530 6 InISR
rlabel m2contact 13389 2650 13389 2650 6 n_317
rlabel m2contact 13341 5122 13341 5122 6 n_476
rlabel m2contact 13245 4570 13245 4570 6 StatusReg[3]
rlabel m2contact 13197 5626 13197 5626 6 n_475
rlabel m2contact 12837 5482 12837 5482 6 n_368
rlabel m2contact 12813 4090 12813 4090 6 n_234
rlabel m2contact 12741 2338 12741 2338 6 SysBus[2]
rlabel m2contact 12693 5266 12693 5266 6 n_109
rlabel m2contact 12669 4810 12669 4810 6 n_237
rlabel m2contact 12645 4618 12645 4618 6 n_108
rlabel m2contact 12597 2722 12597 2722 6 StatusReg[2]
rlabel m2contact 12597 3826 12597 3826 6 n_149
rlabel m2contact 12573 4210 12573 4210 6 n_148
rlabel m2contact 12549 5002 12549 5002 6 n_152
rlabel m2contact 12525 2674 12525 2674 6 n_320
rlabel m2contact 12501 6178 12501 6178 6 n_97
rlabel m2contact 12477 7210 12477 7210 6 IRQ2
rlabel m2contact 12477 6634 12477 6634 6 n_113
rlabel m2contact 12453 5122 12453 5122 6 n_476
rlabel m2contact 12405 6298 12405 6298 6 n_194
rlabel m2contact 12405 2530 12405 2530 6 n_15
rlabel m2contact 12381 2290 12381 2290 6 n_37
rlabel m2contact 12357 5050 12357 5050 4 n_132
rlabel m2contact 12333 5818 12333 5818 4 n_165
rlabel m2contact 12309 3394 12309 3394 4 stateSub[0]
rlabel m2contact 12285 4978 12285 4978 4 n_235
rlabel m2contact 12285 3802 12285 3802 4 n_231
rlabel m2contact 12261 4498 12261 4498 4 OpcodeCondIn[2]
rlabel m2contact 12237 3802 12237 3802 4 n_231
rlabel m2contact 12213 2818 12213 2818 4 n_159
rlabel m2contact 12213 5698 12213 5698 4 stateSub[1]
rlabel m2contact 12189 3538 12189 3538 4 n_202
rlabel m2contact 12189 4090 12189 4090 4 n_234
rlabel m2contact 12117 5266 12117 5266 4 n_84
rlabel m2contact 12117 4954 12117 4954 4 n_172
rlabel m2contact 12093 3514 12093 3514 4 stateSub[2]
rlabel m2contact 12069 6322 12069 6322 4 n_89
rlabel m2contact 12021 4114 12021 4114 4 n_354
rlabel m2contact 12021 4498 12021 4498 4 OpcodeCondIn[2]
rlabel m2contact 11997 5482 11997 5482 4 n_181
rlabel m2contact 11997 6466 11997 6466 4 n_79
rlabel m2contact 11961 5122 11961 5122 4 n_269
rlabel m2contact 11961 4114 11961 4114 4 n_269
rlabel m2contact 11949 5218 11949 5218 4 n_7
rlabel m2contact 11949 3586 11949 3586 4 n_302
rlabel m2contact 11925 4114 11925 4114 4 n_269
rlabel m2contact 11925 4978 11925 4978 4 OpcodeCondIn[6]
rlabel m2contact 11901 3394 11901 3394 4 stateSub[0]
rlabel m2contact 11877 4642 11877 4642 4 n_65
rlabel m2contact 11853 7234 11853 7234 4 n_207
rlabel m2contact 11853 2818 11853 2818 4 n_207
rlabel m2contact 11829 4114 11829 4114 4 n_151
rlabel m2contact 11829 2266 11829 2266 4 n_44
rlabel m2contact 11805 7210 11805 7210 4 n_30
rlabel m2contact 11781 3538 11781 3538 4 n_150
rlabel m2contact 11757 7258 11757 7258 4 n_190
rlabel m2contact 11757 4690 11757 4690 4 n_190
rlabel m2contact 11757 4642 11757 4642 4 n_206
rlabel m2contact 11757 2866 11757 2866 4 n_206
rlabel m2contact 11733 7258 11733 7258 4 n_190
rlabel m2contact 11733 5386 11733 5386 4 OpcodeCondIn[3]
rlabel m2contact 11709 3610 11709 3610 4 n_226
rlabel m2contact 11685 4954 11685 4954 4 n_172
rlabel m2contact 11661 4090 11661 4090 4 n_234
rlabel m2contact 11637 4018 11637 4018 4 n_300
rlabel m2contact 11613 7234 11613 7234 4 n_207
rlabel m2contact 11613 4666 11613 4666 4 n_193
rlabel m2contact 11589 2482 11589 2482 4 n_217
rlabel m2contact 11589 5218 11589 5218 4 n_83
rlabel m2contact 11565 4642 11565 4642 4 n_206
rlabel m2contact 11565 3154 11565 3154 4 n_214
rlabel m2contact 11517 3586 11517 3586 4 n_198
rlabel m2contact 11493 4234 11493 4234 4 state[0]
rlabel m2contact 11493 3970 11493 3970 4 n_249
rlabel m2contact 11469 5890 11469 5890 4 IntReq
rlabel m2contact 11469 4594 11469 4594 4 n_136
rlabel m2contact 11445 4642 11445 4642 4 n_137
rlabel m2contact 11421 2458 11421 2458 4 n_40
rlabel m2contact 11421 4474 11421 4474 4 n_197
rlabel m2contact 11397 3658 11397 3658 4 n_29
rlabel m2contact 11373 3322 11373 3322 4 n_163
rlabel m2contact 11349 7186 11349 7186 4 n_5
rlabel m2contact 11301 2818 11301 2818 4 n_207
rlabel m2contact 11301 3610 11301 3610 4 nIRQ
rlabel m2contact 11253 2818 11253 2818 4 n_255
rlabel m2contact 11253 5050 11253 5050 4 n_132
rlabel m2contact 11205 2194 11205 2194 4 OpcodeCondIn[1]
rlabel m2contact 11181 6610 11181 6610 4 OpcodeCondIn[0]
rlabel m2contact 11181 4138 11181 4138 4 n_185
rlabel m2contact 11157 5338 11157 5338 4 n_72
rlabel m2contact 11157 2050 11157 2050 4 n_72
rlabel m2contact 11133 7210 11133 7210 4 n_30
rlabel m2contact 11133 7186 11133 7186 4 n_239
rlabel m2contact 11109 4498 11109 4498 4 OpcodeCondIn[2]
rlabel m2contact 11085 2050 11085 2050 4 n_72
rlabel m2contact 11085 3658 11085 3658 4 n_29
rlabel m2contact 11061 3874 11061 3874 4 n_264
rlabel m2contact 11037 4258 11037 4258 4 n_177
rlabel m2contact 11013 2842 11013 2842 4 n_32
rlabel m2contact 11013 6610 11013 6610 4 n_25
rlabel m2contact 10989 6826 10989 6826 4 OpcodeCondIn[7]
rlabel m2contact 10965 5050 10965 5050 4 n_132
rlabel m2contact 10917 4138 10917 4138 4 n_57
rlabel m2contact 10893 3322 10893 3322 4 n_163
rlabel m2contact 10869 3082 10869 3082 4 n_76
rlabel m2contact 10845 2050 10845 2050 4 Flags[0]
rlabel m2contact 10821 3682 10821 3682 4 n_33
rlabel m2contact 10797 2458 10797 2458 4 n_40
rlabel m2contact 10773 3082 10773 3082 4 n_76
rlabel m2contact 10725 4882 10725 4882 4 AluOR[1]
rlabel m2contact 10701 2674 10701 2674 4 n_320
rlabel m2contact 10677 4882 10677 4882 4 n_280
rlabel m2contact 10653 4282 10653 4282 4 n_321
rlabel m2contact 10653 2578 10653 2578 4 n_10
rlabel m2contact 10605 2194 10605 2194 4 OpcodeCondIn[1]
rlabel m2contact 10605 3682 10605 3682 4 n_353
rlabel m2contact 10581 2050 10581 2050 4 Flags[0]
rlabel m2contact 10557 2074 10557 2074 4 n_308
rlabel m2contact 10557 6250 10557 6250 4 n_351
rlabel m2contact 10533 2098 10533 2098 4 CFlag
rlabel m2contact 10509 7186 10509 7186 4 n_239
rlabel m2contact 10509 4546 10509 4546 4 n_307
rlabel m2contact 10485 5698 10485 5698 4 stateSub[1]
rlabel m2contact 10461 7162 10461 7162 4 n_238
rlabel m2contact 10413 7138 10413 7138 4 n_75
rlabel m2contact 10413 3586 10413 3586 4 n_198
rlabel m2contact 10389 3274 10389 3274 4 state[1]
rlabel m2contact 10365 3082 10365 3082 4 n_76
rlabel m2contact 10329 5194 10329 5194 4 n_82
rlabel m2contact 10329 3586 10329 3586 4 n_82
rlabel m2contact 10317 5482 10317 5482 4 n_181
rlabel m2contact 10317 2626 10317 2626 4 n_95
rlabel m2contact 10293 3586 10293 3586 4 n_82
rlabel m2contact 10293 4954 10293 4954 4 n_172
rlabel m2contact 10269 4306 10269 4306 4 n_192
rlabel m2contact 10245 3586 10245 3586 4 n_140
rlabel m2contact 10245 2314 10245 2314 4 n_51
rlabel m2contact 10221 3658 10221 3658 4 n_29
rlabel m2contact 10197 5698 10197 5698 4 stateSub[1]
rlabel m2contact 10173 5482 10173 5482 4 n_98
rlabel m2contact 10149 7114 10149 7114 4 n_63
rlabel m2contact 10149 7090 10149 7090 4 n_6
rlabel m2contact 10125 6826 10125 6826 4 OpcodeCondIn[7]
rlabel m2contact 10125 2626 10125 2626 4 OpcodeCondIn[7]
rlabel m2contact 10101 2626 10101 2626 4 OpcodeCondIn[7]
rlabel m2contact 10101 3970 10101 3970 4 n_249
rlabel m2contact 10077 5458 10077 5458 4 OpcodeCondIn[4]
rlabel m2contact 10053 2122 10053 2122 4 n_26
rlabel m2contact 10029 4258 10029 4258 4 n_177
rlabel m2contact 10029 2626 10029 2626 4 n_177
rlabel m2contact 10005 2410 10005 2410 4 n_344
rlabel m2contact 10005 2218 10005 2218 4 n_175
rlabel m2contact 9981 2842 9981 2842 4 n_32
rlabel m2contact 9957 3922 9957 3922 4 n_290
rlabel m2contact 9957 2410 9957 2410 4 PcEn
rlabel m2contact 9933 4162 9933 4162 4 n_99
rlabel m2contact 9909 5314 9909 5314 4 n_68
rlabel m2contact 9885 3178 9885 3178 4 n_245
rlabel m2contact 9861 3802 9861 3802 4 n_231
rlabel m2contact 9861 4162 9861 4162 4 n_127
rlabel m2contact 9837 3394 9837 3394 4 stateSub[0]
rlabel m2contact 9813 5314 9813 5314 4 n_73
rlabel m2contact 9789 2170 9789 2170 4 n_179
rlabel m2contact 9765 2842 9765 2842 4 n_133
rlabel m2contact 9765 3922 9765 3922 4 n_170
rlabel m2contact 9741 2626 9741 2626 4 n_177
rlabel m2contact 9741 3970 9741 3970 4 n_249
rlabel m2contact 9717 2890 9717 2890 4 n_191
rlabel m2contact 9693 6706 9693 6706 4 n_222
rlabel m2contact 9693 2170 9693 2170 4 n_222
rlabel m2contact 9669 3586 9669 3586 4 n_140
rlabel m2contact 9645 3802 9645 3802 4 n_231
rlabel m2contact 9621 5074 9621 5074 4 n_139
rlabel m2contact 9597 3802 9597 3802 4 n_201
rlabel m2contact 9573 6538 9573 6538 4 n_145
rlabel m2contact 9573 3586 9573 3586 4 n_145
rlabel m2contact 9549 6250 9549 6250 4 n_351
rlabel m2contact 9525 7066 9525 7066 4 n_173
rlabel m2contact 9525 6922 9525 6922 4 n_18
rlabel m2contact 9501 2170 9501 2170 4 n_222
rlabel m2contact 9501 2626 9501 2626 4 n_246
rlabel m2contact 9477 6490 9477 6490 4 n_236
rlabel m2contact 9453 5146 9453 5146 4 n_205
rlabel m2contact 9429 3274 9429 3274 4 state[1]
rlabel m2contact 9405 3586 9405 3586 4 n_145
rlabel m2contact 9405 5146 9405 5146 4 n_123
rlabel m2contact 9381 5698 9381 5698 4 stateSub[1]
rlabel m2contact 9357 3586 9357 3586 4 n_121
rlabel m2contact 9333 2146 9333 2146 4 n_87
rlabel m2contact 9333 6490 9333 6490 4 n_8
rlabel m2contact 9333 2170 9333 2170 4 n_8
rlabel m2contact 9309 6922 9309 6922 4 n_256
rlabel m2contact 9309 3514 9309 3514 4 stateSub[2]
rlabel m2contact 9285 3490 9285 3490 4 n_182
rlabel m2contact 9261 2170 9261 2170 4 n_8
rlabel m2contact 9261 3946 9261 3946 4 n_250
rlabel m2contact 9237 2194 9237 2194 4 OpcodeCondIn[1]
rlabel m2contact 9213 7042 9213 7042 4 n_71
rlabel m2contact 9189 6802 9189 6802 4 n_20
rlabel m2contact 9165 4186 9165 4186 4 n_70
rlabel m2contact 9141 6946 9141 6946 4 n_293
rlabel m2contact 9117 4186 9117 4186 4 n_162
rlabel m2contact 9093 6562 9093 6562 4 PcSel[2]
rlabel m2contact 9069 5818 9069 5818 4 n_165
rlabel m2contact 9045 7018 9045 7018 4 n_161
rlabel m2contact 9045 6946 9045 6946 4 ImmSel
rlabel m2contact 8997 4594 8997 4594 4 n_136
rlabel m2contact 8973 3970 8973 3970 4 n_249
rlabel m2contact 8949 5506 8949 5506 4 OpcodeCondIn[5]
rlabel m2contact 8925 4258 8925 4258 4 n_177
rlabel m2contact 8877 5458 8877 5458 4 OpcodeCondIn[4]
rlabel m2contact 8853 6994 8853 6994 4 n_254
rlabel m2contact 8853 5434 8853 5434 4 n_240
rlabel m2contact 8805 6970 8805 6970 4 n_228
rlabel m2contact 8805 3898 8805 3898 4 n_266
rlabel m2contact 8781 2218 8781 2218 4 n_175
rlabel m2contact 8757 6946 8757 6946 4 ImmSel
rlabel m2contact 8757 3898 8757 3898 4 n_263
rlabel m2contact 8733 5986 8733 5986 4 n_291
rlabel m2contact 8733 3874 8733 3874 4 n_264
rlabel m2contact 8709 3034 8709 3034 4 n_287
rlabel m2contact 8685 6922 8685 6922 4 n_256
rlabel m2contact 8685 6154 8685 6154 4 n_312
rlabel m2contact 8661 6898 8661 6898 4 n_277
rlabel m2contact 8661 5602 8661 5602 4 n_261
rlabel m2contact 8661 3034 8661 3034 4 n_261
rlabel m2contact 8637 4498 8637 4498 4 OpcodeCondIn[2]
rlabel m2contact 8613 3034 8613 3034 4 n_261
rlabel m2contact 8613 3082 8613 3082 4 n_76
rlabel m2contact 8565 2794 8565 2794 4 n_39
rlabel m2contact 8541 4258 8541 4258 4 n_177
rlabel m2contact 8493 6754 8493 6754 4 n_304
rlabel m2contact 8469 5362 8469 5362 4 n_282
rlabel m2contact 8445 6874 8445 6874 4 n_117
rlabel m2contact 8445 6754 8445 6754 4 PcWe
rlabel m2contact 8421 3034 8421 3034 4 n_77
rlabel m2contact 8397 6850 8397 6850 4 n_314
rlabel m2contact 8373 5362 8373 5362 4 n_14
rlabel m2contact 8325 6826 8325 6826 4 OpcodeCondIn[7]
rlabel m2contact 8301 6802 8301 6802 4 n_20
rlabel m2contact 8301 6778 8301 6778 4 n_171
rlabel m2contact 8253 6754 8253 6754 4 PcWe
rlabel m2contact 8253 4282 8253 4282 4 n_321
rlabel m2contact 8229 6706 8229 6706 4 n_222
rlabel m2contact 8229 4306 8229 4306 4 n_192
rlabel m2contact 8205 6730 8205 6730 4 n_340
rlabel m2contact 8205 6298 8205 6298 4 n_194
rlabel m2contact 8181 6706 8181 6706 4 n_190
rlabel m2contact 8181 4690 8181 4690 4 n_190
rlabel m2contact 8157 4762 8157 4762 4 n_363
rlabel m2contact 8157 4282 8157 4282 4 n_118
rlabel m2contact 8133 6706 8133 6706 4 n_190
rlabel m2contact 8133 4954 8133 4954 4 n_172
rlabel m2contact 8109 2890 8109 2890 4 n_191
rlabel m2contact 8085 4114 8085 4114 4 n_151
rlabel m2contact 8061 3850 8061 3850 4 n_168
rlabel m2contact 8037 2242 8037 2242 4 n_91
rlabel m2contact 8013 4114 8013 4114 4 n_43
rlabel m2contact 7989 6682 7989 6682 4 n_55
rlabel m2contact 7989 3514 7989 3514 4 stateSub[2]
rlabel m2contact 7941 6658 7941 6658 4 n_134
rlabel m2contact 7941 4954 7941 4954 4 n_172
rlabel m2contact 7941 2242 7941 2242 4 n_172
rlabel m2contact 7917 2242 7917 2242 4 n_172
rlabel m2contact 7917 3394 7917 3394 4 stateSub[0]
rlabel m2contact 7893 6634 7893 6634 4 n_113
rlabel m2contact 7893 2890 7893 2890 4 n_191
rlabel m2contact 7845 2266 7845 2266 4 n_44
rlabel m2contact 7845 3586 7845 3586 4 n_121
rlabel m2contact 7797 6610 7797 6610 4 n_25
rlabel m2contact 7797 3874 7797 3874 4 n_264
rlabel m2contact 7773 4258 7773 4258 4 n_177
rlabel m2contact 7725 6586 7725 6586 4 n_122
rlabel m2contact 7725 2458 7725 2458 4 n_40
rlabel m2contact 7701 6418 7701 6418 4 n_120
rlabel m2contact 7701 5170 7701 5170 4 n_278
rlabel m2contact 7677 3586 7677 3586 4 n_121
rlabel m2contact 7629 6562 7629 6562 4 PcSel[2]
rlabel m2contact 7629 4954 7629 4954 4 n_172
rlabel m2contact 7605 6322 7605 6322 4 n_89
rlabel m2contact 7581 4666 7581 4666 4 n_193
rlabel m2contact 7557 6538 7557 6538 4 n_145
rlabel m2contact 7557 3586 7557 3586 4 ENB
rlabel m2contact 7509 3010 7509 3010 4 n_323
rlabel m2contact 7485 5818 7485 5818 4 n_165
rlabel m2contact 7437 5818 7437 5818 4 n_102
rlabel m2contact 7437 3898 7437 3898 4 n_263
rlabel m2contact 7389 6514 7389 6514 4 n_66
rlabel m2contact 7389 3010 7389 3010 4 n_323
rlabel m2contact 7365 6490 7365 6490 4 n_8
rlabel m2contact 7365 3802 7365 3802 4 n_201
rlabel m2contact 7341 2962 7341 2962 4 n_80
rlabel m2contact 7317 6466 7317 6466 4 n_79
rlabel m2contact 7293 4474 7293 4474 4 n_197
rlabel m2contact 7269 2290 7269 2290 4 n_37
rlabel m2contact 7245 2314 7245 2314 4 n_51
rlabel m2contact 7245 6322 7245 6322 4 n_89
rlabel m2contact 7221 6442 7221 6442 4 n_21
rlabel m2contact 7173 6418 7173 6418 4 n_120
rlabel m2contact 7173 6154 7173 6154 4 n_312
rlabel m2contact 7149 2338 7149 2338 4 SysBus[2]
rlabel m2contact 7125 3874 7125 3874 4 n_264
rlabel m2contact 7101 2338 7101 2338 4 Flags[2]
rlabel m2contact 7101 2794 7101 2794 4 n_39
rlabel m2contact 7029 6394 7029 6394 4 n_243
rlabel m2contact 6981 3946 6981 3946 4 n_250
rlabel m2contact 6957 5890 6957 5890 4 IntReq
rlabel m2contact 6933 4306 6933 4306 4 n_192
rlabel m2contact 6885 4474 6885 4474 4 n_197
rlabel m2contact 6861 4210 6861 4210 4 n_148
rlabel m2contact 6813 5890 6813 5890 4 n_347
rlabel m2contact 6789 2338 6789 2338 4 Flags[2]
rlabel m2contact 6765 6250 6765 6250 4 n_351
rlabel m2contact 6717 2770 6717 2770 4 n_362
rlabel m2contact 6693 4210 6693 4210 4 n_148
rlabel m2contact 6669 6370 6669 6370 4 n_244
rlabel m2contact 6621 2362 6621 2362 4 n_200
rlabel m2contact 6597 2386 6597 2386 4 n_61
rlabel m2contact 6573 4042 6573 4042 4 n_147
rlabel m2contact 6525 2410 6525 2410 4 PcEn
rlabel m2contact 6501 4042 6501 4042 4 n_348
rlabel m2contact 6477 2434 6477 2434 4 n_336
rlabel m2contact 6453 6346 6453 6346 4 n_227
rlabel m2contact 6429 4762 6429 4762 4 n_363
rlabel m2contact 6429 2434 6429 2434 4 n_363
rlabel m2contact 6405 2794 6405 2794 4 n_39
rlabel m2contact 6405 4738 6405 4738 4 n_298
rlabel m2contact 6381 6322 6381 6322 4 n_89
rlabel m2contact 6381 2458 6381 2458 4 n_40
rlabel m2contact 6357 4834 6357 4834 4 n_267
rlabel m2contact 6333 6322 6333 6322 4 Rs1Sel[1]
rlabel m2contact 6309 6322 6309 6322 4 Rs1Sel[1]
rlabel m2contact 6309 2674 6309 2674 4 n_320
rlabel m2contact 6285 4306 6285 4306 4 n_192
rlabel m2contact 6285 2458 6285 2458 4 n_192
rlabel m2contact 6261 5026 6261 5026 4 n_195
rlabel m2contact 6261 2770 6261 2770 4 n_362
rlabel m2contact 6237 2434 6237 2434 4 n_363
rlabel m2contact 6237 3658 6237 3658 4 n_29
rlabel m2contact 6213 6298 6213 6298 4 n_194
rlabel m2contact 6213 5026 6213 5026 4 n_153
rlabel m2contact 6213 2770 6213 2770 4 n_153
rlabel m2contact 6189 3754 6189 3754 4 n_169
rlabel m2contact 6165 6274 6165 6274 4 n_345
rlabel m2contact 6165 4066 6165 4066 4 n_220
rlabel m2contact 6141 2458 6141 2458 4 n_192
rlabel m2contact 6141 3754 6141 3754 4 Flags[3]
rlabel m2contact 6117 6250 6117 6250 4 n_351
rlabel m2contact 6117 3850 6117 3850 4 n_168
rlabel m2contact 6093 3178 6093 3178 4 n_245
rlabel m2contact 6069 5122 6069 5122 4 n_269
rlabel m2contact 6045 4498 6045 4498 4 OpcodeCondIn[2]
rlabel m2contact 6021 2482 6021 2482 4 n_217
rlabel m2contact 6021 4834 6021 4834 4 n_267
rlabel m2contact 5997 5866 5997 5866 4 n_100
rlabel m2contact 5973 2770 5973 2770 4 n_153
rlabel m2contact 5973 4858 5973 4858 4 n_268
rlabel m2contact 5949 6058 5949 6058 4 n_93
rlabel m2contact 5949 2482 5949 2482 4 n_93
rlabel m2contact 5925 6010 5925 6010 4 n_45
rlabel m2contact 5901 2482 5901 2482 4 n_93
rlabel m2contact 5901 2770 5901 2770 4 n_474
rlabel m2contact 5877 4570 5877 4570 4 StatusReg[3]
rlabel m2contact 5853 2962 5853 2962 4 n_80
rlabel m2contact 5829 5122 5829 5122 4 n_208
rlabel m2contact 5781 2506 5781 2506 4 n_19
rlabel m2contact 5781 3082 5781 3082 4 n_76
rlabel m2contact 5757 6226 5757 6226 4 n_154
rlabel m2contact 5733 5506 5733 5506 4 OpcodeCondIn[5]
rlabel m2contact 5709 2530 5709 2530 4 n_15
rlabel m2contact 5685 5458 5685 5458 4 OpcodeCondIn[4]
rlabel m2contact 5661 3874 5661 3874 4 n_264
rlabel m2contact 5589 2674 5589 2674 4 n_320
rlabel m2contact 5565 4882 5565 4882 4 n_280
rlabel m2contact 5565 3490 5565 3490 4 n_182
rlabel m2contact 5493 4066 5493 4066 4 n_220
rlabel m2contact 5445 4498 5445 4498 4 OpcodeCondIn[2]
rlabel m2contact 5421 2674 5421 2674 4 n_107
rlabel m2contact 5397 6202 5397 6202 4 n_315
rlabel m2contact 5397 6178 5397 6178 4 n_97
rlabel m2contact 5373 6154 5373 6154 4 n_312
rlabel m2contact 5373 6130 5373 6130 4 n_213
rlabel m2contact 5349 6106 5349 6106 4 SysBus[1]
rlabel m2contact 5301 6082 5301 6082 4 n_94
rlabel m2contact 5301 3514 5301 3514 4 stateSub[2]
rlabel m2contact 5277 6058 5277 6058 4 n_93
rlabel m2contact 5277 6034 5277 6034 4 n_125
rlabel m2contact 5253 5650 5253 5650 4 n_46
rlabel m2contact 5229 6010 5229 6010 4 n_45
rlabel m2contact 5229 2554 5229 2554 4 n_128
rlabel m2contact 5205 4066 5205 4066 4 n_220
rlabel m2contact 5181 5986 5181 5986 4 n_291
rlabel m2contact 5181 5866 5181 5866 4 n_100
rlabel m2contact 5181 2554 5181 2554 4 n_100
rlabel m2contact 5157 3178 5157 3178 4 n_245
rlabel m2contact 5133 2554 5133 2554 4 n_100
rlabel m2contact 5133 3898 5133 3898 4 n_263
rlabel m2contact 5061 5962 5061 5962 4 n_274
rlabel m2contact 5061 2578 5061 2578 4 n_10
rlabel m2contact 5013 5938 5013 5938 4 n_242
rlabel m2contact 4965 5914 4965 5914 4 n_478
rlabel m2contact 4965 5890 4965 5890 4 n_347
rlabel m2contact 4941 2602 4941 2602 4 n_306
rlabel m2contact 4941 4066 4941 4066 4 n_220
rlabel m2contact 4917 5866 4917 5866 4 n_100
rlabel m2contact 4893 5842 4893 5842 4 n_253
rlabel m2contact 4893 5818 4893 5818 4 n_102
rlabel m2contact 4869 4954 4869 4954 4 n_172
rlabel m2contact 4845 4258 4845 4258 4 n_177
rlabel m2contact 4821 5794 4821 5794 4 SysBus[0]
rlabel m2contact 4821 4858 4821 4858 4 n_268
rlabel m2contact 4773 3010 4773 3010 4 n_323
rlabel m2contact 4749 4810 4749 4810 4 n_237
rlabel m2contact 4749 3394 4749 3394 4 stateSub[0]
rlabel m2contact 4725 5698 4725 5698 4 stateSub[1]
rlabel m2contact 4677 5770 4677 5770 4 StatusReg[0]
rlabel m2contact 4677 2626 4677 2626 4 n_246
rlabel m2contact 4653 4978 4653 4978 4 OpcodeCondIn[6]
rlabel m2contact 4629 5002 4629 5002 4 n_152
rlabel m2contact 4629 3946 4629 3946 4 n_250
rlabel m2contact 4593 4282 4593 4282 4 n_118
rlabel m2contact 4593 2626 4593 2626 4 n_118
rlabel m2contact 4581 4690 4581 4690 4 n_190
rlabel m2contact 4557 2626 4557 2626 4 n_118
rlabel m2contact 4557 4258 4557 4258 4 n_177
rlabel m2contact 4533 4234 4533 4234 4 state[0]
rlabel m2contact 4485 5746 4485 5746 4 n_24
rlabel m2contact 4485 5722 4485 5722 4 n_141
rlabel m2contact 4461 3394 4461 3394 4 stateSub[0]
rlabel m2contact 4413 5698 4413 5698 4 stateSub[1]
rlabel m2contact 4389 4666 4389 4666 4 n_193
rlabel m2contact 4341 2650 4341 2650 4 n_317
rlabel m2contact 4317 5674 4317 5674 4 n_284
rlabel m2contact 4293 4066 4293 4066 4 n_220
rlabel m2contact 4269 5602 4269 5602 4 n_261
rlabel m2contact 4245 2794 4245 2794 4 n_39
rlabel m2contact 4221 5650 4221 5650 4 n_46
rlabel m2contact 4221 4666 4221 4666 4 n_193
rlabel m2contact 4197 5626 4197 5626 4 n_475
rlabel m2contact 4197 5602 4197 5602 4 StatusReg[2]
rlabel m2contact 4197 2722 4197 2722 4 StatusReg[2]
rlabel m2contact 4173 5602 4173 5602 4 StatusReg[2]
rlabel m2contact 4173 2794 4173 2794 4 LrSel
rlabel m2contact 4125 2674 4125 2674 4 n_107
rlabel m2contact 4101 2698 4101 2698 4 n_473
rlabel m2contact 4077 5578 4077 5578 4 IRQ1
rlabel m2contact 4029 5554 4029 5554 4 n_286
rlabel m2contact 4029 2722 4029 2722 4 StatusReg[2]
rlabel m2contact 4005 2746 4005 2746 4 n_215
rlabel m2contact 3981 2770 3981 2770 4 n_474
rlabel m2contact 3981 4738 3981 4738 4 n_298
rlabel m2contact 3909 2794 3909 2794 4 LrSel
rlabel m2contact 3861 4378 3861 4378 4 n_270
rlabel m2contact 3813 5530 3813 5530 4 n_130
rlabel m2contact 3789 5506 3789 5506 4 OpcodeCondIn[5]
rlabel m2contact 3765 5482 3765 5482 4 n_98
rlabel m2contact 3717 2818 3717 2818 4 n_255
rlabel m2contact 3693 5458 3693 5458 4 OpcodeCondIn[4]
rlabel m2contact 3669 5434 3669 5434 4 n_240
rlabel m2contact 3645 3178 3645 3178 4 n_245
rlabel m2contact 3597 2842 3597 2842 4 n_133
rlabel m2contact 3573 4498 3573 4498 4 OpcodeCondIn[2]
rlabel m2contact 3549 4690 3549 4690 4 n_190
rlabel m2contact 3525 5050 3525 5050 4 n_132
rlabel m2contact 3501 2914 3501 2914 4 n_155
rlabel m2contact 3477 3514 3477 3514 4 stateSub[2]
rlabel m2contact 3453 4306 3453 4306 4 n_192
rlabel m2contact 3453 4690 3453 4690 4 n_3
rlabel m2contact 3357 5410 3357 5410 4 n_11
rlabel m2contact 3333 5386 3333 5386 4 OpcodeCondIn[3]
rlabel m2contact 3333 2866 3333 2866 4 n_206
rlabel m2contact 3309 4978 3309 4978 4 OpcodeCondIn[6]
rlabel m2contact 3261 2890 3261 2890 4 n_191
rlabel m2contact 3261 4618 3261 4618 4 n_108
rlabel m2contact 3213 5362 3213 5362 4 n_14
rlabel m2contact 3213 2914 3213 2914 4 n_155
rlabel m2contact 3189 4714 3189 4714 4 n_92
rlabel m2contact 3165 4546 3165 4546 4 n_307
rlabel m2contact 3141 5314 3141 5314 4 n_73
rlabel m2contact 3117 2938 3117 2938 4 n_212
rlabel m2contact 3117 4714 3117 4714 4 n_17
rlabel m2contact 3093 5338 3093 5338 4 n_72
rlabel m2contact 3093 4306 3093 4306 4 n_192
rlabel m2contact 3069 5314 3069 5314 4 state[1]
rlabel m2contact 3069 3274 3069 3274 4 state[1]
rlabel m2contact 3045 4306 3045 4306 4 n_106
rlabel m2contact 3021 5314 3021 5314 4 state[1]
rlabel m2contact 3021 3538 3021 3538 4 n_150
rlabel m2contact 2997 5290 2997 5290 4 n_105
rlabel m2contact 2997 2962 2997 2962 4 n_80
rlabel m2contact 2973 5266 2973 5266 4 n_84
rlabel m2contact 2949 2986 2949 2986 4 n_316
rlabel m2contact 2925 3922 2925 3922 4 n_170
rlabel m2contact 2901 5242 2901 5242 4 n_257
rlabel m2contact 2901 4474 2901 4474 4 n_197
rlabel m2contact 2877 3106 2877 3106 4 n_223
rlabel m2contact 2853 3922 2853 3922 4 n_265
rlabel m2contact 2781 5218 2781 5218 4 n_83
rlabel m2contact 2781 3106 2781 3106 4 n_67
rlabel m2contact 2733 5194 2733 5194 4 n_82
rlabel m2contact 2685 5170 2685 5170 4 n_278
rlabel m2contact 2685 3010 2685 3010 4 n_323
rlabel m2contact 2661 5146 2661 5146 4 n_123
rlabel m2contact 2637 3274 2637 3274 4 state[1]
rlabel m2contact 2613 5122 2613 5122 4 n_208
rlabel m2contact 2613 5098 2613 5098 4 n_62
rlabel m2contact 2589 4666 2589 4666 4 n_193
rlabel m2contact 2565 5074 2565 5074 4 n_139
rlabel m2contact 2565 3082 2565 3082 4 n_76
rlabel m2contact 2541 5050 2541 5050 4 n_132
rlabel m2contact 2541 3154 2541 3154 4 n_214
rlabel m2contact 2517 4858 2517 4858 4 n_268
rlabel m2contact 2493 3058 2493 3058 4 n_34
rlabel m2contact 2493 4066 2493 4066 4 n_220
rlabel m2contact 2469 4666 2469 4666 4 n_193
rlabel m2contact 2445 5026 2445 5026 4 n_153
rlabel m2contact 2445 3082 2445 3082 4 n_76
rlabel m2contact 2397 5002 2397 5002 4 n_152
rlabel m2contact 2397 3034 2397 3034 4 n_77
rlabel m2contact 2397 4474 2397 4474 4 n_197
rlabel m2contact 2397 3058 2397 3058 4 n_197
rlabel m2contact 2373 3058 2373 3058 4 n_197
rlabel m2contact 2373 3850 2373 3850 4 n_168
rlabel m2contact 2349 3082 2349 3082 4 n_76
rlabel m2contact 2325 3106 2325 3106 4 n_67
rlabel m2contact 2301 4978 2301 4978 4 OpcodeCondIn[6]
rlabel m2contact 2277 4954 2277 4954 4 n_172
rlabel m2contact 2277 4930 2277 4930 4 n_167
rlabel m2contact 2253 4378 2253 4378 4 n_270
rlabel m2contact 2229 4042 2229 4042 4 n_348
rlabel m2contact 2205 4378 2205 4378 4 n_247
rlabel m2contact 2181 4906 2181 4906 4 n_49
rlabel m2contact 2157 4306 2157 4306 4 n_106
rlabel m2contact 2109 4882 2109 4882 4 n_280
rlabel m2contact 2109 4306 2109 4306 4 n_143
rlabel m2contact 2085 4858 2085 4858 4 n_268
rlabel m2contact 2061 4834 2061 4834 4 n_267
rlabel m2contact 2061 3130 2061 3130 4 n_334
rlabel m2contact 2037 3154 2037 3154 4 n_214
rlabel m2contact 2037 4786 2037 4786 4 n_248
rlabel m2contact 2013 3346 2013 3346 4 n_110
rlabel m2contact 1989 4810 1989 4810 4 n_237
rlabel m2contact 1941 4786 1941 4786 4 n_248
rlabel m2contact 1941 3178 1941 3178 4 n_245
rlabel m2contact 1917 4186 1917 4186 4 n_162
rlabel m2contact 1893 3202 1893 3202 4 n_54
rlabel m2contact 1869 4186 1869 4186 4 AluEn
rlabel m2contact 1845 4762 1845 4762 4 n_363
rlabel m2contact 1821 3226 1821 3226 4 n_343
rlabel m2contact 1797 4738 1797 4738 4 n_298
rlabel m2contact 1773 3250 1773 3250 4 n_275
rlabel m2contact 1749 3274 1749 3274 4 state[1]
rlabel m2contact 1725 4714 1725 4714 4 n_17
rlabel m2contact 1701 4690 1701 4690 4 n_3
rlabel m2contact 1701 4666 1701 4666 4 n_193
rlabel m2contact 1677 4666 1677 4666 4 n_193
rlabel m2contact 1629 4642 1629 4642 4 n_137
rlabel m2contact 1605 4618 1605 4618 4 n_108
rlabel m2contact 1581 4594 1581 4594 4 n_136
rlabel m2contact 1533 3298 1533 3298 4 n_305
rlabel m2contact 1509 4570 1509 4570 4 StatusReg[3]
rlabel m2contact 1485 4546 1485 4546 4 n_307
rlabel m2contact 1437 4522 1437 4522 4 n_86
rlabel m2contact 1413 4498 1413 4498 4 OpcodeCondIn[2]
rlabel m2contact 1389 4474 1389 4474 4 n_197
rlabel m2contact 1365 3874 1365 3874 4 n_264
rlabel m2contact 1317 4450 1317 4450 4 n_178
rlabel m2contact 1293 4258 1293 4258 4 n_177
rlabel m2contact 1269 4426 1269 4426 4 n_138
rlabel m2contact 1221 4402 1221 4402 4 n_303
rlabel m2contact 1197 4258 1197 4258 4 n_177
rlabel m2contact 1173 4378 1173 4378 4 n_247
rlabel m2contact 1173 4210 1173 4210 4 n_148
rlabel m2contact 1149 4354 1149 4354 4 n_224
rlabel m2contact 1149 4330 1149 4330 4 n_12
rlabel m2contact 1101 4306 1101 4306 4 n_143
rlabel m2contact 1101 3442 1101 3442 4 n_233
rlabel m2contact 1077 4282 1077 4282 4 n_118
rlabel m2contact 1077 3322 1077 3322 4 n_163
rlabel m2contact 1053 4258 1053 4258 4 n_177
rlabel m2contact 1053 3442 1053 3442 4 n_210
rlabel m2contact 1029 4234 1029 4234 4 state[0]
rlabel m2contact 981 3394 981 3394 4 stateSub[0]
rlabel m2contact 981 3802 981 3802 4 n_201
rlabel m2contact 957 4210 957 4210 4 n_148
rlabel m2contact 957 3346 957 3346 4 n_110
rlabel m2contact 933 3850 933 3850 4 n_168
rlabel m2contact 909 4186 909 4186 4 AluEn
rlabel m2contact 885 3850 885 3850 4 n_186
rlabel m2contact 861 3370 861 3370 4 n_42
rlabel m2contact 837 4162 837 4162 4 n_127
rlabel m2contact 813 4138 813 4138 4 n_57
rlabel m2contact 765 3394 765 3394 4 stateSub[0]
rlabel m2contact 765 4114 765 4114 4 n_43
rlabel m2contact 741 4090 741 4090 4 n_234
rlabel m2contact 717 4066 717 4066 4 n_220
rlabel m2contact 717 3658 717 3658 4 n_29
rlabel m2contact 669 3658 669 3658 4 nOE
rlabel m2contact 645 4042 645 4042 4 n_348
rlabel m2contact 621 3418 621 3418 4 n_288
rlabel m2contact 597 4018 597 4018 4 n_300
rlabel m2contact 549 3994 549 3994 4 n_251
rlabel m2contact 525 3970 525 3970 4 n_249
rlabel m2contact 501 3946 501 3946 4 n_250
rlabel m2contact 453 3922 453 3922 4 n_265
rlabel m2contact 405 3898 405 3898 4 n_263
rlabel m2contact 381 3874 381 3874 4 n_264
rlabel m2contact 357 3850 357 3850 4 n_186
rlabel m2contact 333 3442 333 3442 4 n_210
rlabel m2contact 309 3826 309 3826 4 n_149
rlabel m2contact 285 3802 285 3802 4 n_201
rlabel m2contact 237 3778 237 3778 4 nME
rlabel m2contact 237 3754 237 3754 4 Flags[3]
rlabel m2contact 189 3466 189 3466 4 n_183
rlabel m2contact 189 3730 189 3730 4 n_360
rlabel m2contact 165 3490 165 3490 4 n_182
rlabel m2contact 165 3706 165 3706 4 n_310
rlabel m2contact 141 3514 141 3514 4 stateSub[2]
rlabel m2contact 141 3682 141 3682 4 n_353
rlabel m2contact 117 3538 117 3538 4 n_150
rlabel m2contact 117 3562 117 3562 4 n_309
rlabel m2contact 24813 1097 24813 1097 6 OpcodeCondIn[2]
rlabel m2contact 24813 113 24813 113 8 OpcodeCondIn[2]
rlabel m2contact 24789 857 24789 857 6 OpcodeCondIn[7]
rlabel m2contact 24789 89 24789 89 8 OpcodeCondIn[7]
rlabel m2contact 24765 737 24765 737 8 OpcodeCondIn[6]
rlabel m2contact 24765 65 24765 65 8 OpcodeCondIn[6]
rlabel m2contact 24741 1121 24741 1121 6 OpcodeCondIn[4]
rlabel m2contact 24741 41 24741 41 8 OpcodeCondIn[4]
rlabel m2contact 24717 617 24717 617 8 OpcodeCondIn[0]
rlabel m2contact 24717 137 24717 137 8 OpcodeCondIn[0]
rlabel m2contact 24717 65 24717 65 8 OpcodeCondIn[5]
rlabel m2contact 24717 17 24717 17 8 OpcodeCondIn[5]
rlabel m2contact 24717 641 24717 641 8 n_359
rlabel m2contact 24597 641 24597 641 8 n_359
rlabel m2contact 24549 689 24549 689 8 n_331
rlabel m2contact 23625 833 23625 833 6 MemEn
rlabel m2contact 23517 785 23517 785 8 n_81
rlabel m2contact 23397 713 23397 713 8 n_119
rlabel m2contact 23277 377 23277 377 8 PcSel[0]
rlabel metal2 23247 641 23247 641 8 IrWe
rlabel m2contact 23229 641 23229 641 8 IrWe
rlabel m2contact 23181 1025 23181 1025 6 n_203
rlabel m2contact 23013 857 23013 857 6 OpcodeCondIn[7]
rlabel m2contact 22653 569 22653 569 8 n_60
rlabel m2contact 22581 1121 22581 1121 6 OpcodeCondIn[4]
rlabel m2contact 22437 161 22437 161 8 Op1Sel
rlabel m2contact 22365 641 22365 641 8 n_326
rlabel m2contact 22005 857 22005 857 6 OpcodeCondIn[7]
rlabel m2contact 21933 353 21933 353 8 PcSel[1]
rlabel m2contact 21765 857 21765 857 6 OpcodeCondIn[7]
rlabel m2contact 21669 497 21669 497 8 n_27
rlabel m2contact 21357 473 21357 473 8 LrEn
rlabel m2contact 21285 929 21285 929 6 n_41
rlabel m2contact 21237 809 21237 809 6 n_158
rlabel m2contact 21021 953 21021 953 6 n_196
rlabel m2contact 20901 617 20901 617 8 OpcodeCondIn[0]
rlabel m2contact 20853 521 20853 521 8 n_180
rlabel m2contact 20829 401 20829 401 8 n_142
rlabel m2contact 20697 1073 20697 1073 6 ImmSel
rlabel m2contact 20637 209 20637 209 8 Flags[1]
rlabel m2contact 20589 545 20589 545 8 n_28
rlabel m2contact 20565 857 20565 857 6 OpcodeCondIn[7]
rlabel m2contact 20469 1097 20469 1097 6 OpcodeCondIn[2]
rlabel m2contact 20373 665 20373 665 8 n_58
rlabel m2contact 20109 593 20109 593 8 n_211
rlabel m2contact 20085 1169 20085 1169 6 n_219
rlabel m2contact 20037 425 20037 425 8 n_335
rlabel m2contact 19821 1049 19821 1049 6 n_96
rlabel m2contact 19749 905 19749 905 6 n_341
rlabel m2contact 19701 1193 19701 1193 6 n_230
rlabel m2contact 19677 641 19677 641 8 n_326
rlabel m2contact 19461 1217 19461 1217 6 n_276
rlabel m2contact 19269 881 19269 881 6 n_187
rlabel m2contact 19245 641 19245 641 8 n_225
rlabel m2contact 19233 89 19233 89 8 LrSel
rlabel m2contact 19197 1145 19197 1145 6 n_176
rlabel m2contact 18933 233 18933 233 8 n_50
rlabel m2contact 18837 449 18837 449 8 n_189
rlabel m2contact 18813 281 18813 281 8 n_160
rlabel m2contact 18501 1097 18501 1097 6 OpcodeCondIn[2]
rlabel m2contact 18285 257 18285 257 8 n_258
rlabel m2contact 18213 1001 18213 1001 6 n_216
rlabel m2contact 18165 689 18165 689 8 n_331
rlabel m2contact 18117 689 18117 689 8 n_283
rlabel m2contact 17853 977 17853 977 6 n_221
rlabel m2contact 17769 113 17769 113 8 LrWe
rlabel m2contact 17745 473 17745 473 8 LrEn
rlabel m2contact 17109 761 17109 761 8 n_324
rlabel m2contact 16965 1121 16965 1121 6 OpcodeCondIn[4]
rlabel m2contact 16941 137 16941 137 8 n_115
rlabel m2contact 16773 1217 16773 1217 6 n_276
rlabel m2contact 16749 1145 16749 1145 6 n_176
rlabel m2contact 16677 185 16677 185 8 n_111
rlabel m2contact 16581 473 16581 473 8 n_252
rlabel m2contact 16485 1121 16485 1121 6 OpcodeCondIn[4]
rlabel m2contact 16281 377 16281 377 8 PcSel[0]
rlabel m2contact 16269 1145 16269 1145 6 WdSel
rlabel m2contact 16197 641 16197 641 8 n_225
rlabel m2contact 16173 1217 16173 1217 6 n_157
rlabel m2contact 16101 329 16101 329 8 n_272
rlabel m2contact 15981 641 15981 641 8 n_85
rlabel m2contact 15717 497 15717 497 8 n_27
rlabel m2contact 15669 689 15669 689 8 n_283
rlabel m2contact 15573 377 15573 377 8 n_114
rlabel m2contact 15477 689 15477 689 8 Op2Sel[1]
rlabel m2contact 15237 497 15237 497 8 AluWe
rlabel m2contact 14817 353 14817 353 8 PcSel[1]
rlabel m2contact 14229 305 14229 305 8 n_188
rlabel m2contact 14205 737 14205 737 8 OpcodeCondIn[6]
rlabel m2contact 14181 353 14181 353 8 n_166
rlabel m2contact 14109 737 14109 737 8 OpcodeCondIn[6]
rlabel m2contact 14013 233 14013 233 8 n_50
rlabel m2contact 13989 761 13989 761 8 n_324
rlabel m2contact 13797 281 13797 281 8 n_160
rlabel m2contact 12981 425 12981 425 8 n_335
rlabel m2contact 12861 17 12861 17 8 n_53
rlabel m2contact 12837 1121 12837 1121 6 OpcodeCondIn[4]
rlabel m2contact 12429 1049 12429 1049 6 n_96
rlabel m2contact 12333 1001 12333 1001 4 n_216
rlabel m2contact 12237 881 12237 881 4 n_187
rlabel m2contact 12141 425 12141 425 2 n_90
rlabel m2contact 11973 233 11973 233 2 n_327
rlabel m2contact 11913 41 11913 41 2 PcSel[2]
rlabel m2contact 11757 1001 11757 1001 4 n_259
rlabel m2contact 11685 857 11685 857 4 OpcodeCondIn[7]
rlabel m2contact 11517 281 11517 281 2 n_78
rlabel m2contact 11325 881 11325 881 4 Op2Sel[0]
rlabel m2contact 11277 1049 11277 1049 4 n_330
rlabel m2contact 11205 833 11205 833 4 MemEn
rlabel m2contact 11157 833 11157 833 4 n_279
rlabel m2contact 10941 137 10941 137 2 n_115
rlabel m2contact 10893 377 10893 377 2 n_114
rlabel m2contact 10845 137 10845 137 2 Flags[0]
rlabel m2contact 10797 233 10797 233 2 n_327
rlabel m2contact 10749 257 10749 257 2 n_258
rlabel m2contact 10725 329 10725 329 2 n_272
rlabel m2contact 10461 257 10461 257 2 n_229
rlabel m2contact 10437 329 10437 329 2 n_146
rlabel m2contact 10437 233 10437 233 2 PcWe
rlabel m2contact 10365 1217 10365 1217 4 n_157
rlabel m2contact 10341 17 10341 17 2 n_53
rlabel m2contact 10125 1121 10125 1121 4 OpcodeCondIn[4]
rlabel m2contact 10101 857 10101 857 4 OpcodeCondIn[7]
rlabel m2contact 10029 1121 10029 1121 4 OpcodeCondIn[4]
rlabel metal2 9975 17 9975 17 2 PcEn
rlabel m2contact 9957 17 9957 17 2 PcEn
rlabel m2contact 9909 1193 9909 1193 4 n_230
rlabel m2contact 9573 1169 9573 1169 4 n_219
rlabel m2contact 9453 329 9453 329 2 n_146
rlabel m2contact 9357 329 9357 329 2 n_135
rlabel m2contact 9213 1097 9213 1097 4 OpcodeCondIn[2]
rlabel m2contact 9093 41 9093 41 2 PcSel[2]
rlabel m2contact 9045 1073 9045 1073 4 ImmSel
rlabel m2contact 8997 1049 8997 1049 4 n_330
rlabel m2contact 8949 1073 8949 1073 4 n_289
rlabel m2contact 8925 1145 8925 1145 4 WdSel
rlabel m2contact 8901 1049 8901 1049 4 n_241
rlabel m2contact 8877 1121 8877 1121 4 OpcodeCondIn[4]
rlabel m2contact 8637 1097 8637 1097 4 OpcodeCondIn[2]
rlabel m2contact 8565 1073 8565 1073 4 n_289
rlabel m2contact 8541 953 8541 953 4 n_196
rlabel m2contact 8517 1049 8517 1049 4 n_241
rlabel m2contact 8493 1025 8493 1025 4 n_203
rlabel m2contact 8445 233 8445 233 2 PcWe
rlabel m2contact 8373 233 8373 233 2 n_74
rlabel m2contact 8349 1001 8349 1001 4 n_259
rlabel m2contact 8325 977 8325 977 4 n_221
rlabel m2contact 8109 545 8109 545 2 n_28
rlabel m2contact 8013 545 8013 545 2 n_112
rlabel m2contact 7941 953 7941 953 4 n_196
rlabel m2contact 7821 857 7821 857 4 OpcodeCondIn[7]
rlabel m2contact 7749 833 7749 833 4 n_279
rlabel m2contact 7653 545 7653 545 2 n_112
rlabel m2contact 7485 761 7485 761 2 n_324
rlabel m2contact 7449 161 7449 161 2 Op1Sel
rlabel m2contact 7197 761 7197 761 2 n_313
rlabel m2contact 7101 161 7101 161 2 Flags[2]
rlabel m2contact 6549 833 6549 833 4 n_262
rlabel m2contact 6429 929 6429 929 4 n_41
rlabel m2contact 6285 905 6285 905 4 n_341
rlabel m2contact 5973 881 5973 881 4 Op2Sel[0]
rlabel m2contact 5733 65 5733 65 2 OpcodeCondIn[5]
rlabel m2contact 5613 737 5613 737 2 OpcodeCondIn[6]
rlabel m2contact 5517 737 5517 737 2 OpcodeCondIn[6]
rlabel m2contact 5493 857 5493 857 4 OpcodeCondIn[7]
rlabel m2contact 5445 833 5445 833 4 n_262
rlabel m2contact 5325 809 5325 809 4 n_158
rlabel m2contact 5181 785 5181 785 2 n_81
rlabel m2contact 5085 617 5085 617 2 OpcodeCondIn[0]
rlabel m2contact 5013 617 5013 617 2 n_367
rlabel m2contact 4989 761 4989 761 2 n_313
rlabel m2contact 4653 737 4653 737 2 OpcodeCondIn[6]
rlabel m2contact 4581 713 4581 713 2 n_119
rlabel m2contact 4497 689 4497 689 2 Op2Sel[1]
rlabel m2contact 4437 665 4437 665 2 n_58
rlabel m2contact 4413 641 4413 641 2 n_85
rlabel m2contact 4173 89 4173 89 2 LrSel
rlabel m2contact 3621 617 3621 617 2 n_367
rlabel m2contact 3405 593 3405 593 2 n_211
rlabel m2contact 3357 569 3357 569 2 n_60
rlabel m2contact 3141 545 3141 545 2 n_112
rlabel m2contact 3069 521 3069 521 2 n_180
rlabel m2contact 3021 497 3021 497 2 AluWe
rlabel m2contact 2925 473 2925 473 2 n_252
rlabel m2contact 2877 449 2877 449 2 n_189
rlabel m2contact 2853 425 2853 425 2 n_90
rlabel m2contact 2805 401 2805 401 2 n_142
rlabel m2contact 2757 377 2757 377 2 n_114
rlabel m2contact 2709 353 2709 353 2 n_166
rlabel m2contact 2301 113 2301 113 2 LrWe
rlabel m2contact 2181 329 2181 329 2 n_135
rlabel m2contact 2157 305 2157 305 2 n_188
rlabel m2contact 2133 281 2133 281 2 n_78
rlabel m2contact 1341 257 1341 257 2 n_229
rlabel m2contact 1221 233 1221 233 2 n_74
rlabel m2contact 1005 185 1005 185 2 n_111
rlabel metal2 927 185 927 185 2 AluEn
rlabel m2contact 909 185 909 185 2 AluEn
rlabel m2contact 237 185 237 185 2 Flags[3]
rlabel m2contact 21477 8235 21477 8235 6 AluOR[0]
rlabel m2contact 21477 8091 21477 8091 6 AluOR[0]
rlabel m2contact 21453 8187 21453 8187 6 RwSel[0]
rlabel m2contact 21453 8091 21453 8091 6 RwSel[0]
rlabel m2contact 21429 8187 21429 8187 6 Rs1Sel[0]
rlabel m2contact 21429 8115 21429 8115 6 Rs1Sel[0]
rlabel m2contact 21405 8211 21405 8211 6 RegWe
rlabel m2contact 21405 8115 21405 8115 6 RegWe
rlabel m2contact 21381 8211 21381 8211 6 Rs1Sel[1]
rlabel m2contact 21381 8163 21381 8163 6 Rs1Sel[1]
rlabel m2contact 21357 8163 21357 8163 6 RwSel[1]
rlabel m2contact 21357 8139 21357 8139 6 RwSel[1]
rlabel m2contact 21333 8259 21333 8259 6 CFlag
rlabel m2contact 21333 8139 21333 8139 6 CFlag
rlabel m2contact 21309 8259 21309 8259 6 ALE
rlabel m2contact 18765 8091 18765 8091 6 RwSel[0]
rlabel m2contact 16773 8115 16773 8115 6 RegWe
rlabel m2contact 16029 8139 16029 8139 6 CFlag
rlabel m2contact 14253 8163 14253 8163 6 RwSel[1]
rlabel m2contact 13485 8187 13485 8187 6 Rs1Sel[0]
rlabel m2contact 6309 8211 6309 8211 4 Rs1Sel[1]
rlabel m2contact 5613 8235 5613 8235 4 AluOR[0]
rlabel m2contact 3405 8211 3405 8211 4 nWait
rlabel m2contact 429 8211 429 8211 4 nWait
rlabel m2contact 237 8235 237 8235 4 nME
rlabel metal2 23619 0 23631 0 8 MemEn
rlabel metal2 23235 0 23247 0 8 IrWe
rlabel metal2 20691 0 20703 0 8 ImmSel
rlabel metal2 19227 0 19239 0 8 LrSel
rlabel metal2 17763 0 17775 0 8 LrWe
rlabel metal2 17739 0 17751 0 8 LrEn
rlabel metal2 16275 0 16287 0 8 PcSel[0]
rlabel metal2 14811 0 14823 0 8 PcSel[1]
rlabel metal2 11907 0 11919 0 2 PcSel[2]
rlabel metal2 10431 0 10443 0 2 PcWe
rlabel metal2 9963 0 9975 0 2 PcEn
rlabel metal2 8919 0 8931 0 2 WdSel
rlabel metal2 7443 0 7455 0 2 Op1Sel
rlabel metal2 5967 0 5979 0 2 Op2Sel[0]
rlabel metal2 4491 0 4503 0 2 Op2Sel[1]
rlabel metal2 3015 0 3027 0 2 AluWe
rlabel metal2 915 0 927 0 2 AluEn
rlabel metal2 25683 2164 25683 2176 6 SysBus[1]
rlabel metal2 25683 2140 25683 2152 6 SysBus[0]
rlabel metal2 25683 2116 25683 2128 6 SysBus[3]
rlabel metal2 25683 2092 25683 2104 6 SysBus[2]
rlabel metal2 25683 2068 25683 2080 6 OpcodeCondIn[3]
rlabel metal2 25683 2044 25683 2056 6 OpcodeCondIn[1]
rlabel metal2 25683 131 25683 143 8 OpcodeCondIn[0]
rlabel metal2 25683 107 25683 119 8 OpcodeCondIn[2]
rlabel metal2 25683 83 25683 95 8 OpcodeCondIn[7]
rlabel metal2 25683 59 25683 71 8 OpcodeCondIn[6]
rlabel metal2 25683 35 25683 47 8 OpcodeCondIn[4]
rlabel metal2 25683 11 25683 23 8 OpcodeCondIn[5]
rlabel metal2 25683 8253 25683 8265 6 CFlag
rlabel metal2 25683 8205 25683 8217 6 RegWe
rlabel metal2 25683 8181 25683 8193 6 RwSel[0]
rlabel metal2 25683 8157 25683 8169 6 Rs1Sel[1]
rlabel metal2 25683 8133 25683 8145 6 RwSel[1]
rlabel metal2 25683 8109 25683 8121 6 Rs1Sel[0]
rlabel metal2 25683 8085 25683 8097 6 AluOR[0]
rlabel metal2 25359 0 25559 0 1 GND!
rlabel space 25359 8276 25560 8276 5 GND!
rlabel metal2 -1500 203 -1500 215 2 Flags[1]
rlabel metal2 -1500 179 -1500 191 2 Flags[3]
rlabel metal2 -1500 155 -1500 167 2 Flags[2]
rlabel metal2 -1500 131 -1500 143 2 Flags[0]
rlabel metal2 -1500 8253 -1500 8265 4 ALE
rlabel metal2 -1500 8229 -1500 8241 4 nME
rlabel metal2 -1500 8205 -1500 8217 4 nWait
rlabel metal2 -1500 3652 -1500 3664 4 nOE
rlabel metal2 -1500 3628 -1500 3640 4 nWE
rlabel metal2 -1500 3604 -1500 3616 4 nIRQ
rlabel metal2 -1500 3580 -1500 3592 4 ENB
rlabel metal2 -1377 0 -1177 0 1 Vdd!
rlabel metal2 -1377 8276 -1177 8276 5 Vdd!
rlabel metal2 25683 4876 25683 4888 6 AluOR[1]
rlabel metal2 -1161 8276 -1149 8276 5 SDO
rlabel metal2 -1113 8276 -1101 8276 5 Clock
rlabel metal2 -1137 8276 -1125 8276 5 Test
rlabel metal2 -1089 8276 -1077 8276 5 nReset
rlabel metal2 -1161 0 -1149 0 1 SDI
rlabel metal2 -1137 0 -1125 0 1 Test
rlabel metal2 -1113 0 -1101 0 1 Clock
rlabel metal2 -1089 0 -1077 0 1 nReset
<< end >>
